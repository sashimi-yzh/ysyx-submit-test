//Generate the verilog at 2025-12-27T22:02:25 by iSTA.
module ysyx_25080222 (
clock,
io_interrupt,
io_master_arready,
io_master_arvalid,
io_master_awready,
io_master_awvalid,
io_master_bready,
io_master_bvalid,
io_master_rlast,
io_master_rready,
io_master_rvalid,
io_master_wlast,
io_master_wready,
io_master_wvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_awready,
io_slave_awvalid,
io_slave_bready,
io_slave_bvalid,
io_slave_rlast,
io_slave_rready,
io_slave_rvalid,
io_slave_wlast,
io_slave_wready,
io_slave_wvalid,
reset,
io_master_araddr,
io_master_arburst,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_awaddr,
io_master_awburst,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_bid,
io_master_bresp,
io_master_rdata,
io_master_rid,
io_master_rresp,
io_master_wdata,
io_master_wstrb,
io_slave_araddr,
io_slave_arburst,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_awaddr,
io_slave_awburst,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_bid,
io_slave_bresp,
io_slave_rdata,
io_slave_rid,
io_slave_rresp,
io_slave_wdata,
io_slave_wstrb
);

input clock ;
input io_interrupt ;
input io_master_arready ;
output io_master_arvalid ;
input io_master_awready ;
output io_master_awvalid ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_rlast ;
output io_master_rready ;
input io_master_rvalid ;
output io_master_wlast ;
input io_master_wready ;
output io_master_wvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
output io_slave_awready ;
input io_slave_awvalid ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_rlast ;
input io_slave_rready ;
output io_slave_rvalid ;
input io_slave_wlast ;
output io_slave_wready ;
input io_slave_wvalid ;
input reset ;
output [31:0] io_master_araddr ;
output [1:0] io_master_arburst ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [31:0] io_master_awaddr ;
output [1:0] io_master_awburst ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
input [3:0] io_master_bid ;
input [1:0] io_master_bresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [1:0] io_master_rresp ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [31:0] io_slave_araddr ;
input [1:0] io_slave_arburst ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [31:0] io_slave_awaddr ;
input [1:0] io_slave_awburst ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
output [3:0] io_slave_bid ;
output [1:0] io_slave_bresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;
output [1:0] io_slave_rresp ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;

wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire _08922_ ;
wire _08923_ ;
wire _08924_ ;
wire _08925_ ;
wire _08926_ ;
wire _08927_ ;
wire _08928_ ;
wire _08929_ ;
wire _08930_ ;
wire _08931_ ;
wire _08932_ ;
wire _08933_ ;
wire _08934_ ;
wire _08935_ ;
wire _08936_ ;
wire _08937_ ;
wire _08938_ ;
wire _08939_ ;
wire _08940_ ;
wire _08941_ ;
wire _08942_ ;
wire _08943_ ;
wire _08944_ ;
wire _08945_ ;
wire _08946_ ;
wire _08947_ ;
wire _08948_ ;
wire _08949_ ;
wire _08950_ ;
wire _08951_ ;
wire _08952_ ;
wire _08953_ ;
wire _08954_ ;
wire _08955_ ;
wire _08956_ ;
wire _08957_ ;
wire _08958_ ;
wire _08959_ ;
wire _08960_ ;
wire _08961_ ;
wire _08962_ ;
wire _08963_ ;
wire _08964_ ;
wire _08965_ ;
wire _08966_ ;
wire _08967_ ;
wire _08968_ ;
wire _08969_ ;
wire _08970_ ;
wire _08971_ ;
wire _08972_ ;
wire _08973_ ;
wire _08974_ ;
wire _08975_ ;
wire _08976_ ;
wire _08977_ ;
wire _08978_ ;
wire _08979_ ;
wire _08980_ ;
wire _08981_ ;
wire _08982_ ;
wire _08983_ ;
wire _08984_ ;
wire _08985_ ;
wire _08986_ ;
wire _08987_ ;
wire _08988_ ;
wire _08989_ ;
wire _08990_ ;
wire _08991_ ;
wire _08992_ ;
wire _08993_ ;
wire _08994_ ;
wire _08995_ ;
wire _08996_ ;
wire _08997_ ;
wire _08998_ ;
wire _08999_ ;
wire _09000_ ;
wire _09001_ ;
wire _09002_ ;
wire _09003_ ;
wire _09004_ ;
wire _09005_ ;
wire _09006_ ;
wire _09007_ ;
wire _09008_ ;
wire _09009_ ;
wire _09010_ ;
wire _09011_ ;
wire _09012_ ;
wire _09013_ ;
wire _09014_ ;
wire _09015_ ;
wire _09016_ ;
wire _09017_ ;
wire _09018_ ;
wire _09019_ ;
wire _09020_ ;
wire _09021_ ;
wire _09022_ ;
wire _09023_ ;
wire _09024_ ;
wire _09025_ ;
wire _09026_ ;
wire _09027_ ;
wire _09028_ ;
wire _09029_ ;
wire _09030_ ;
wire _09031_ ;
wire _09032_ ;
wire _09033_ ;
wire _09034_ ;
wire _09035_ ;
wire _09036_ ;
wire _09037_ ;
wire _09038_ ;
wire _09039_ ;
wire _09040_ ;
wire _09041_ ;
wire _09042_ ;
wire _09043_ ;
wire _09044_ ;
wire _09045_ ;
wire _09046_ ;
wire _09047_ ;
wire _09048_ ;
wire _09049_ ;
wire _09050_ ;
wire _09051_ ;
wire _09052_ ;
wire _09053_ ;
wire _09054_ ;
wire _09055_ ;
wire _09056_ ;
wire _09057_ ;
wire _09058_ ;
wire _09059_ ;
wire _09060_ ;
wire _09061_ ;
wire _09062_ ;
wire _09063_ ;
wire _09064_ ;
wire _09065_ ;
wire _09066_ ;
wire _09067_ ;
wire _09068_ ;
wire _09069_ ;
wire _09070_ ;
wire _09071_ ;
wire _09072_ ;
wire _09073_ ;
wire _09074_ ;
wire _09075_ ;
wire _09076_ ;
wire _09077_ ;
wire _09078_ ;
wire _09079_ ;
wire _09080_ ;
wire _09081_ ;
wire _09082_ ;
wire _09083_ ;
wire _09084_ ;
wire _09085_ ;
wire _09086_ ;
wire _09087_ ;
wire _09088_ ;
wire _09089_ ;
wire _09090_ ;
wire _09091_ ;
wire _09092_ ;
wire _09093_ ;
wire _09094_ ;
wire _09095_ ;
wire _09096_ ;
wire _09097_ ;
wire _09098_ ;
wire _09099_ ;
wire _09100_ ;
wire _09101_ ;
wire _09102_ ;
wire _09103_ ;
wire _09104_ ;
wire _09105_ ;
wire _09106_ ;
wire _09107_ ;
wire _09108_ ;
wire _09109_ ;
wire _09110_ ;
wire _09111_ ;
wire _09112_ ;
wire _09113_ ;
wire _09114_ ;
wire _09115_ ;
wire _09116_ ;
wire _09117_ ;
wire _09118_ ;
wire _09119_ ;
wire _09120_ ;
wire _09121_ ;
wire _09122_ ;
wire _09123_ ;
wire _09124_ ;
wire _09125_ ;
wire _09126_ ;
wire _09127_ ;
wire _09128_ ;
wire _09129_ ;
wire _09130_ ;
wire _09131_ ;
wire _09132_ ;
wire _09133_ ;
wire _09134_ ;
wire _09135_ ;
wire _09136_ ;
wire _09137_ ;
wire _09138_ ;
wire _09139_ ;
wire _09140_ ;
wire _09141_ ;
wire _09142_ ;
wire _09143_ ;
wire _09144_ ;
wire _09145_ ;
wire _09146_ ;
wire _09147_ ;
wire _09148_ ;
wire _09149_ ;
wire _09150_ ;
wire _09151_ ;
wire _09152_ ;
wire _09153_ ;
wire _09154_ ;
wire _09155_ ;
wire _09156_ ;
wire _09157_ ;
wire _09158_ ;
wire _09159_ ;
wire _09160_ ;
wire _09161_ ;
wire _09162_ ;
wire _09163_ ;
wire _09164_ ;
wire _09165_ ;
wire _09166_ ;
wire _09167_ ;
wire _09168_ ;
wire _09169_ ;
wire _09170_ ;
wire _09171_ ;
wire _09172_ ;
wire _09173_ ;
wire _09174_ ;
wire _09175_ ;
wire _09176_ ;
wire _09177_ ;
wire _09178_ ;
wire _09179_ ;
wire _09180_ ;
wire _09181_ ;
wire _09182_ ;
wire _09183_ ;
wire _09184_ ;
wire _09185_ ;
wire _09186_ ;
wire _09187_ ;
wire _09188_ ;
wire _09189_ ;
wire _09190_ ;
wire _09191_ ;
wire _09192_ ;
wire _09193_ ;
wire _09194_ ;
wire _09195_ ;
wire _09196_ ;
wire _09197_ ;
wire _09198_ ;
wire _09199_ ;
wire _09200_ ;
wire _09201_ ;
wire _09202_ ;
wire _09203_ ;
wire _09204_ ;
wire _09205_ ;
wire _09206_ ;
wire _09207_ ;
wire _09208_ ;
wire _09209_ ;
wire _09210_ ;
wire _09211_ ;
wire _09212_ ;
wire _09213_ ;
wire _09214_ ;
wire _09215_ ;
wire _09216_ ;
wire _09217_ ;
wire _09218_ ;
wire _09219_ ;
wire _09220_ ;
wire _09221_ ;
wire _09222_ ;
wire _09223_ ;
wire _09224_ ;
wire _09225_ ;
wire _09226_ ;
wire _09227_ ;
wire _09228_ ;
wire _09229_ ;
wire _09230_ ;
wire _09231_ ;
wire _09232_ ;
wire _09233_ ;
wire _09234_ ;
wire _09235_ ;
wire _09236_ ;
wire _09237_ ;
wire _09238_ ;
wire _09239_ ;
wire _09240_ ;
wire _09241_ ;
wire _09242_ ;
wire _09243_ ;
wire _09244_ ;
wire _09245_ ;
wire _09246_ ;
wire _09247_ ;
wire _09248_ ;
wire _09249_ ;
wire _09250_ ;
wire _09251_ ;
wire _09252_ ;
wire _09253_ ;
wire _09254_ ;
wire _09255_ ;
wire _09256_ ;
wire _09257_ ;
wire _09258_ ;
wire _09259_ ;
wire _09260_ ;
wire _09261_ ;
wire _09262_ ;
wire _09263_ ;
wire _09264_ ;
wire _09265_ ;
wire _09266_ ;
wire _09267_ ;
wire _09268_ ;
wire _09269_ ;
wire _09270_ ;
wire _09271_ ;
wire _09272_ ;
wire _09273_ ;
wire _09274_ ;
wire _09275_ ;
wire _09276_ ;
wire _09277_ ;
wire _09278_ ;
wire _09279_ ;
wire _09280_ ;
wire _09281_ ;
wire _09282_ ;
wire _09283_ ;
wire _09284_ ;
wire _09285_ ;
wire _09286_ ;
wire _09287_ ;
wire _09288_ ;
wire _09289_ ;
wire _09290_ ;
wire _09291_ ;
wire _09292_ ;
wire _09293_ ;
wire _09294_ ;
wire _09295_ ;
wire _09296_ ;
wire _09297_ ;
wire _09298_ ;
wire _09299_ ;
wire _09300_ ;
wire _09301_ ;
wire _09302_ ;
wire _09303_ ;
wire _09304_ ;
wire _09305_ ;
wire _09306_ ;
wire _09307_ ;
wire _09308_ ;
wire _09309_ ;
wire _09310_ ;
wire _09311_ ;
wire _09312_ ;
wire _09313_ ;
wire _09314_ ;
wire _09315_ ;
wire _09316_ ;
wire _09317_ ;
wire _09318_ ;
wire _09319_ ;
wire _09320_ ;
wire _09321_ ;
wire _09322_ ;
wire _09323_ ;
wire _09324_ ;
wire _09325_ ;
wire _09326_ ;
wire _09327_ ;
wire _09328_ ;
wire _09329_ ;
wire _09330_ ;
wire _09331_ ;
wire _09332_ ;
wire _09333_ ;
wire _09334_ ;
wire _09335_ ;
wire _09336_ ;
wire _09337_ ;
wire _09338_ ;
wire _09339_ ;
wire _09340_ ;
wire _09341_ ;
wire _09342_ ;
wire _09343_ ;
wire _09344_ ;
wire _09345_ ;
wire _09346_ ;
wire _09347_ ;
wire _09348_ ;
wire _09349_ ;
wire _09350_ ;
wire _09351_ ;
wire _09352_ ;
wire _09353_ ;
wire _09354_ ;
wire _09355_ ;
wire _09356_ ;
wire _09357_ ;
wire _09358_ ;
wire _09359_ ;
wire _09360_ ;
wire _09361_ ;
wire _09362_ ;
wire _09363_ ;
wire _09364_ ;
wire _09365_ ;
wire _09366_ ;
wire _09367_ ;
wire _09368_ ;
wire _09369_ ;
wire _09370_ ;
wire _09371_ ;
wire _09372_ ;
wire _09373_ ;
wire _09374_ ;
wire _09375_ ;
wire _09376_ ;
wire _09377_ ;
wire _09378_ ;
wire _09379_ ;
wire _09380_ ;
wire _09381_ ;
wire _09382_ ;
wire _09383_ ;
wire _09384_ ;
wire _09385_ ;
wire _09386_ ;
wire _09387_ ;
wire _09388_ ;
wire _09389_ ;
wire _09390_ ;
wire _09391_ ;
wire _09392_ ;
wire _09393_ ;
wire _09394_ ;
wire _09395_ ;
wire _09396_ ;
wire _09397_ ;
wire _09398_ ;
wire _09399_ ;
wire _09400_ ;
wire _09401_ ;
wire _09402_ ;
wire _09403_ ;
wire _09404_ ;
wire _09405_ ;
wire _09406_ ;
wire _09407_ ;
wire _09408_ ;
wire _09409_ ;
wire _09410_ ;
wire _09411_ ;
wire _09412_ ;
wire _09413_ ;
wire _09414_ ;
wire _09415_ ;
wire _09416_ ;
wire _09417_ ;
wire _09418_ ;
wire _09419_ ;
wire _09420_ ;
wire _09421_ ;
wire _09422_ ;
wire _09423_ ;
wire _09424_ ;
wire _09425_ ;
wire _09426_ ;
wire _09427_ ;
wire _09428_ ;
wire _09429_ ;
wire _09430_ ;
wire _09431_ ;
wire _09432_ ;
wire _09433_ ;
wire _09434_ ;
wire _09435_ ;
wire _09436_ ;
wire _09437_ ;
wire _09438_ ;
wire _09439_ ;
wire _09440_ ;
wire _09441_ ;
wire _09442_ ;
wire _09443_ ;
wire _09444_ ;
wire _09445_ ;
wire _09446_ ;
wire _09447_ ;
wire _09448_ ;
wire _09449_ ;
wire _09450_ ;
wire _09451_ ;
wire _09452_ ;
wire _09453_ ;
wire _09454_ ;
wire _09455_ ;
wire _09456_ ;
wire _09457_ ;
wire _09458_ ;
wire _09459_ ;
wire _09460_ ;
wire _09461_ ;
wire _09462_ ;
wire _09463_ ;
wire _09464_ ;
wire _09465_ ;
wire _09466_ ;
wire _09467_ ;
wire _09468_ ;
wire _09469_ ;
wire _09470_ ;
wire _09471_ ;
wire _09472_ ;
wire _09473_ ;
wire _09474_ ;
wire _09475_ ;
wire _09476_ ;
wire _09477_ ;
wire _09478_ ;
wire _09479_ ;
wire _09480_ ;
wire _09481_ ;
wire _09482_ ;
wire _09483_ ;
wire _09484_ ;
wire _09485_ ;
wire _09486_ ;
wire _09487_ ;
wire _09488_ ;
wire _09489_ ;
wire _09490_ ;
wire _09491_ ;
wire _09492_ ;
wire _09493_ ;
wire _09494_ ;
wire _09495_ ;
wire _09496_ ;
wire _09497_ ;
wire _09498_ ;
wire _09499_ ;
wire _09500_ ;
wire _09501_ ;
wire _09502_ ;
wire _09503_ ;
wire _09504_ ;
wire _09505_ ;
wire _09506_ ;
wire _09507_ ;
wire _09508_ ;
wire _09509_ ;
wire _09510_ ;
wire _09511_ ;
wire _09512_ ;
wire _09513_ ;
wire _09514_ ;
wire _09515_ ;
wire _09516_ ;
wire _09517_ ;
wire _09518_ ;
wire _09519_ ;
wire _09520_ ;
wire _09521_ ;
wire _09522_ ;
wire _09523_ ;
wire _09524_ ;
wire _09525_ ;
wire _09526_ ;
wire _09527_ ;
wire _09528_ ;
wire _09529_ ;
wire _09530_ ;
wire _09531_ ;
wire _09532_ ;
wire _09533_ ;
wire _09534_ ;
wire _09535_ ;
wire _09536_ ;
wire _09537_ ;
wire _09538_ ;
wire _09539_ ;
wire _09540_ ;
wire _09541_ ;
wire _09542_ ;
wire _09543_ ;
wire _09544_ ;
wire _09545_ ;
wire _09546_ ;
wire _09547_ ;
wire _09548_ ;
wire _09549_ ;
wire _09550_ ;
wire _09551_ ;
wire _09552_ ;
wire _09553_ ;
wire _09554_ ;
wire _09555_ ;
wire _09556_ ;
wire _09557_ ;
wire _09558_ ;
wire _09559_ ;
wire _09560_ ;
wire _09561_ ;
wire _09562_ ;
wire _09563_ ;
wire _09564_ ;
wire _09565_ ;
wire _09566_ ;
wire _09567_ ;
wire _09568_ ;
wire _09569_ ;
wire _09570_ ;
wire _09571_ ;
wire _09572_ ;
wire _09573_ ;
wire _09574_ ;
wire _09575_ ;
wire _09576_ ;
wire _09577_ ;
wire _09578_ ;
wire _09579_ ;
wire _09580_ ;
wire _09581_ ;
wire _09582_ ;
wire _09583_ ;
wire _09584_ ;
wire _09585_ ;
wire _09586_ ;
wire _09587_ ;
wire _09588_ ;
wire _09589_ ;
wire _09590_ ;
wire _09591_ ;
wire _09592_ ;
wire _09593_ ;
wire _09594_ ;
wire _09595_ ;
wire _09596_ ;
wire _09597_ ;
wire _09598_ ;
wire _09599_ ;
wire _09600_ ;
wire _09601_ ;
wire _09602_ ;
wire _09603_ ;
wire _09604_ ;
wire _09605_ ;
wire _09606_ ;
wire _09607_ ;
wire _09608_ ;
wire _09609_ ;
wire _09610_ ;
wire _09611_ ;
wire _09612_ ;
wire _09613_ ;
wire _09614_ ;
wire _09615_ ;
wire _09616_ ;
wire _09617_ ;
wire _09618_ ;
wire _09619_ ;
wire _09620_ ;
wire _09621_ ;
wire _09622_ ;
wire _09623_ ;
wire _09624_ ;
wire _09625_ ;
wire _09626_ ;
wire _09627_ ;
wire _09628_ ;
wire _09629_ ;
wire _09630_ ;
wire _09631_ ;
wire _09632_ ;
wire _09633_ ;
wire _09634_ ;
wire _09635_ ;
wire _09636_ ;
wire _09637_ ;
wire _09638_ ;
wire _09639_ ;
wire _09640_ ;
wire _09641_ ;
wire _09642_ ;
wire _09643_ ;
wire _09644_ ;
wire _09645_ ;
wire _09646_ ;
wire _09647_ ;
wire _09648_ ;
wire _09649_ ;
wire _09650_ ;
wire _09651_ ;
wire _09652_ ;
wire _09653_ ;
wire _09654_ ;
wire _09655_ ;
wire _09656_ ;
wire _09657_ ;
wire _09658_ ;
wire _09659_ ;
wire _09660_ ;
wire _09661_ ;
wire _09662_ ;
wire _09663_ ;
wire _09664_ ;
wire _09665_ ;
wire _09666_ ;
wire _09667_ ;
wire _09668_ ;
wire _09669_ ;
wire _09670_ ;
wire _09671_ ;
wire _09672_ ;
wire _09673_ ;
wire _09674_ ;
wire _09675_ ;
wire _09676_ ;
wire _09677_ ;
wire _09678_ ;
wire _09679_ ;
wire _09680_ ;
wire _09681_ ;
wire _09682_ ;
wire _09683_ ;
wire _09684_ ;
wire _09685_ ;
wire _09686_ ;
wire _09687_ ;
wire _09688_ ;
wire _09689_ ;
wire _09690_ ;
wire _09691_ ;
wire _09692_ ;
wire _09693_ ;
wire _09694_ ;
wire _09695_ ;
wire _09696_ ;
wire _09697_ ;
wire _09698_ ;
wire _09699_ ;
wire _09700_ ;
wire _09701_ ;
wire _09702_ ;
wire _09703_ ;
wire _09704_ ;
wire _09705_ ;
wire _09706_ ;
wire _09707_ ;
wire _09708_ ;
wire _09709_ ;
wire _09710_ ;
wire _09711_ ;
wire _09712_ ;
wire _09713_ ;
wire _09714_ ;
wire _09715_ ;
wire _09716_ ;
wire _09717_ ;
wire _09718_ ;
wire _09719_ ;
wire _09720_ ;
wire _09721_ ;
wire _09722_ ;
wire _09723_ ;
wire _09724_ ;
wire _09725_ ;
wire _09726_ ;
wire _09727_ ;
wire _09728_ ;
wire _09729_ ;
wire _09730_ ;
wire _09731_ ;
wire _09732_ ;
wire _09733_ ;
wire _09734_ ;
wire _09735_ ;
wire _09736_ ;
wire _09737_ ;
wire _09738_ ;
wire _09739_ ;
wire _09740_ ;
wire _09741_ ;
wire _09742_ ;
wire _09743_ ;
wire _09744_ ;
wire _09745_ ;
wire _09746_ ;
wire _09747_ ;
wire _09748_ ;
wire _09749_ ;
wire _09750_ ;
wire _09751_ ;
wire _09752_ ;
wire _09753_ ;
wire _09754_ ;
wire _09755_ ;
wire _09756_ ;
wire _09757_ ;
wire _09758_ ;
wire _09759_ ;
wire _09760_ ;
wire _09761_ ;
wire _09762_ ;
wire _09763_ ;
wire _09764_ ;
wire _09765_ ;
wire _09766_ ;
wire _09767_ ;
wire _09768_ ;
wire _09769_ ;
wire _09770_ ;
wire _09771_ ;
wire _09772_ ;
wire _09773_ ;
wire _09774_ ;
wire _09775_ ;
wire _09776_ ;
wire _09777_ ;
wire _09778_ ;
wire _09779_ ;
wire _09780_ ;
wire _09781_ ;
wire _09782_ ;
wire _09783_ ;
wire _09784_ ;
wire _09785_ ;
wire _09786_ ;
wire _09787_ ;
wire _09788_ ;
wire _09789_ ;
wire _09790_ ;
wire _09791_ ;
wire _09792_ ;
wire _09793_ ;
wire _09794_ ;
wire _09795_ ;
wire _09796_ ;
wire _09797_ ;
wire _09798_ ;
wire _09799_ ;
wire _09800_ ;
wire _09801_ ;
wire _09802_ ;
wire _09803_ ;
wire _09804_ ;
wire _09805_ ;
wire _09806_ ;
wire _09807_ ;
wire _09808_ ;
wire _09809_ ;
wire _09810_ ;
wire _09811_ ;
wire _09812_ ;
wire _09813_ ;
wire _09814_ ;
wire _09815_ ;
wire _09816_ ;
wire _09817_ ;
wire _09818_ ;
wire _09819_ ;
wire _09820_ ;
wire _09821_ ;
wire _09822_ ;
wire _09823_ ;
wire _09824_ ;
wire _09825_ ;
wire _09826_ ;
wire _09827_ ;
wire _09828_ ;
wire _09829_ ;
wire _09830_ ;
wire _09831_ ;
wire _09832_ ;
wire _09833_ ;
wire _09834_ ;
wire _09835_ ;
wire _09836_ ;
wire _09837_ ;
wire _09838_ ;
wire _09839_ ;
wire _09840_ ;
wire _09841_ ;
wire _09842_ ;
wire _09843_ ;
wire _09844_ ;
wire _09845_ ;
wire _09846_ ;
wire _09847_ ;
wire _09848_ ;
wire _09849_ ;
wire _09850_ ;
wire _09851_ ;
wire _09852_ ;
wire _09853_ ;
wire _09854_ ;
wire _09855_ ;
wire _09856_ ;
wire _09857_ ;
wire _09858_ ;
wire _09859_ ;
wire _09860_ ;
wire _09861_ ;
wire _09862_ ;
wire _09863_ ;
wire _09864_ ;
wire _09865_ ;
wire _09866_ ;
wire _09867_ ;
wire _09868_ ;
wire _09869_ ;
wire _09870_ ;
wire _09871_ ;
wire _09872_ ;
wire _09873_ ;
wire _09874_ ;
wire _09875_ ;
wire _09876_ ;
wire _09877_ ;
wire _09878_ ;
wire _09879_ ;
wire _09880_ ;
wire _09881_ ;
wire _09882_ ;
wire _09883_ ;
wire _09884_ ;
wire _09885_ ;
wire _09886_ ;
wire _09887_ ;
wire _09888_ ;
wire _09889_ ;
wire _09890_ ;
wire _09891_ ;
wire _09892_ ;
wire _09893_ ;
wire _09894_ ;
wire _09895_ ;
wire _09896_ ;
wire _09897_ ;
wire _09898_ ;
wire _09899_ ;
wire _09900_ ;
wire _09901_ ;
wire _09902_ ;
wire _09903_ ;
wire _09904_ ;
wire _09905_ ;
wire _09906_ ;
wire _09907_ ;
wire _09908_ ;
wire _09909_ ;
wire _09910_ ;
wire _09911_ ;
wire _09912_ ;
wire _09913_ ;
wire _09914_ ;
wire _09915_ ;
wire _09916_ ;
wire _09917_ ;
wire _09918_ ;
wire _09919_ ;
wire _09920_ ;
wire _09921_ ;
wire _09922_ ;
wire _09923_ ;
wire _09924_ ;
wire _09925_ ;
wire _09926_ ;
wire _09927_ ;
wire _09928_ ;
wire _09929_ ;
wire _09930_ ;
wire _09931_ ;
wire _09932_ ;
wire _09933_ ;
wire _09934_ ;
wire _09935_ ;
wire _09936_ ;
wire _09937_ ;
wire _09938_ ;
wire _09939_ ;
wire _09940_ ;
wire _09941_ ;
wire _09942_ ;
wire _09943_ ;
wire _09944_ ;
wire _09945_ ;
wire _09946_ ;
wire _09947_ ;
wire _09948_ ;
wire _09949_ ;
wire _09950_ ;
wire _09951_ ;
wire _09952_ ;
wire _09953_ ;
wire _09954_ ;
wire _09955_ ;
wire _09956_ ;
wire _09957_ ;
wire _09958_ ;
wire _09959_ ;
wire _09960_ ;
wire _09961_ ;
wire _09962_ ;
wire _09963_ ;
wire _09964_ ;
wire _09965_ ;
wire _09966_ ;
wire _09967_ ;
wire _09968_ ;
wire _09969_ ;
wire _09970_ ;
wire _09971_ ;
wire _09972_ ;
wire _09973_ ;
wire _09974_ ;
wire _09975_ ;
wire _09976_ ;
wire _09977_ ;
wire _09978_ ;
wire _09979_ ;
wire _09980_ ;
wire _09981_ ;
wire _09982_ ;
wire _09983_ ;
wire _09984_ ;
wire _09985_ ;
wire _09986_ ;
wire _09987_ ;
wire _09988_ ;
wire _09989_ ;
wire _09990_ ;
wire _09991_ ;
wire _09992_ ;
wire _09993_ ;
wire _09994_ ;
wire _09995_ ;
wire _09996_ ;
wire _09997_ ;
wire _09998_ ;
wire _09999_ ;
wire _10000_ ;
wire _10001_ ;
wire _10002_ ;
wire _10003_ ;
wire _10004_ ;
wire _10005_ ;
wire _10006_ ;
wire _10007_ ;
wire _10008_ ;
wire _10009_ ;
wire _10010_ ;
wire _10011_ ;
wire _10012_ ;
wire _10013_ ;
wire _10014_ ;
wire _10015_ ;
wire _10016_ ;
wire _10017_ ;
wire _10018_ ;
wire _10019_ ;
wire _10020_ ;
wire _10021_ ;
wire _10022_ ;
wire _10023_ ;
wire _10024_ ;
wire _10025_ ;
wire _10026_ ;
wire _10027_ ;
wire _10028_ ;
wire _10029_ ;
wire _10030_ ;
wire _10031_ ;
wire _10032_ ;
wire _10033_ ;
wire _10034_ ;
wire _10035_ ;
wire _10036_ ;
wire _10037_ ;
wire _10038_ ;
wire _10039_ ;
wire _10040_ ;
wire _10041_ ;
wire _10042_ ;
wire _10043_ ;
wire _10044_ ;
wire _10045_ ;
wire _10046_ ;
wire _10047_ ;
wire _10048_ ;
wire _10049_ ;
wire _10050_ ;
wire _10051_ ;
wire _10052_ ;
wire _10053_ ;
wire _10054_ ;
wire _10055_ ;
wire _10056_ ;
wire _10057_ ;
wire _10058_ ;
wire _10059_ ;
wire _10060_ ;
wire _10061_ ;
wire _10062_ ;
wire _10063_ ;
wire _10064_ ;
wire _10065_ ;
wire _10066_ ;
wire _10067_ ;
wire _10068_ ;
wire _10069_ ;
wire _10070_ ;
wire _10071_ ;
wire _10072_ ;
wire _10073_ ;
wire _10074_ ;
wire _10075_ ;
wire _10076_ ;
wire _10077_ ;
wire _10078_ ;
wire _10079_ ;
wire _10080_ ;
wire _10081_ ;
wire _10082_ ;
wire _10083_ ;
wire _10084_ ;
wire _10085_ ;
wire _10086_ ;
wire _10087_ ;
wire _10088_ ;
wire _10089_ ;
wire _10090_ ;
wire _10091_ ;
wire _10092_ ;
wire _10093_ ;
wire _10094_ ;
wire _10095_ ;
wire _10096_ ;
wire _10097_ ;
wire _10098_ ;
wire _10099_ ;
wire _10100_ ;
wire _10101_ ;
wire _10102_ ;
wire _10103_ ;
wire _10104_ ;
wire _10105_ ;
wire _10106_ ;
wire _10107_ ;
wire _10108_ ;
wire _10109_ ;
wire _10110_ ;
wire _10111_ ;
wire _10112_ ;
wire _10113_ ;
wire _10114_ ;
wire _10115_ ;
wire _10116_ ;
wire _10117_ ;
wire _10118_ ;
wire _10119_ ;
wire _10120_ ;
wire _10121_ ;
wire _10122_ ;
wire _10123_ ;
wire _10124_ ;
wire _10125_ ;
wire _10126_ ;
wire _10127_ ;
wire _10128_ ;
wire _10129_ ;
wire _10130_ ;
wire _10131_ ;
wire _10132_ ;
wire _10133_ ;
wire _10134_ ;
wire _10135_ ;
wire _10136_ ;
wire _10137_ ;
wire _10138_ ;
wire _10139_ ;
wire _10140_ ;
wire _10141_ ;
wire _10142_ ;
wire _10143_ ;
wire _10144_ ;
wire _10145_ ;
wire _10146_ ;
wire _10147_ ;
wire _10148_ ;
wire _10149_ ;
wire _10150_ ;
wire _10151_ ;
wire _10152_ ;
wire _10153_ ;
wire _10154_ ;
wire _10155_ ;
wire _10156_ ;
wire _10157_ ;
wire _10158_ ;
wire _10159_ ;
wire _10160_ ;
wire _10161_ ;
wire _10162_ ;
wire _10163_ ;
wire _10164_ ;
wire _10165_ ;
wire _10166_ ;
wire _10167_ ;
wire _10168_ ;
wire _10169_ ;
wire _10170_ ;
wire _10171_ ;
wire _10172_ ;
wire _10173_ ;
wire _10174_ ;
wire _10175_ ;
wire _10176_ ;
wire _10177_ ;
wire _10178_ ;
wire _10179_ ;
wire _10180_ ;
wire _10181_ ;
wire _10182_ ;
wire _10183_ ;
wire _10184_ ;
wire _10185_ ;
wire _10186_ ;
wire _10187_ ;
wire _10188_ ;
wire _10189_ ;
wire _10190_ ;
wire _10191_ ;
wire _10192_ ;
wire _10193_ ;
wire _10194_ ;
wire _10195_ ;
wire _10196_ ;
wire _10197_ ;
wire _10198_ ;
wire _10199_ ;
wire _10200_ ;
wire _10201_ ;
wire _10202_ ;
wire _10203_ ;
wire _10204_ ;
wire _10205_ ;
wire _10206_ ;
wire _10207_ ;
wire _10208_ ;
wire _10209_ ;
wire _10210_ ;
wire _10211_ ;
wire _10212_ ;
wire _10213_ ;
wire _10214_ ;
wire _10215_ ;
wire _10216_ ;
wire _10217_ ;
wire _10218_ ;
wire _10219_ ;
wire _10220_ ;
wire _10221_ ;
wire _10222_ ;
wire _10223_ ;
wire _10224_ ;
wire _10225_ ;
wire _10226_ ;
wire _10227_ ;
wire _10228_ ;
wire _10229_ ;
wire _10230_ ;
wire _10231_ ;
wire _10232_ ;
wire _10233_ ;
wire _10234_ ;
wire _10235_ ;
wire _10236_ ;
wire _10237_ ;
wire _10238_ ;
wire _10239_ ;
wire _10240_ ;
wire _10241_ ;
wire _10242_ ;
wire _10243_ ;
wire _10244_ ;
wire _10245_ ;
wire _10246_ ;
wire _10247_ ;
wire _10248_ ;
wire _10249_ ;
wire _10250_ ;
wire _10251_ ;
wire _10252_ ;
wire _10253_ ;
wire _10254_ ;
wire _10255_ ;
wire _10256_ ;
wire _10257_ ;
wire _10258_ ;
wire _10259_ ;
wire _10260_ ;
wire _10261_ ;
wire _10262_ ;
wire _10263_ ;
wire _10264_ ;
wire _10265_ ;
wire _10266_ ;
wire _10267_ ;
wire _10268_ ;
wire _10269_ ;
wire _10270_ ;
wire _10271_ ;
wire _10272_ ;
wire _10273_ ;
wire _10274_ ;
wire _10275_ ;
wire _10276_ ;
wire _10277_ ;
wire _10278_ ;
wire _10279_ ;
wire _10280_ ;
wire _10281_ ;
wire _10282_ ;
wire _10283_ ;
wire _10284_ ;
wire _10285_ ;
wire _10286_ ;
wire _10287_ ;
wire _10288_ ;
wire _10289_ ;
wire _10290_ ;
wire _10291_ ;
wire _10292_ ;
wire _10293_ ;
wire _10294_ ;
wire _10295_ ;
wire _10296_ ;
wire _10297_ ;
wire _10298_ ;
wire _10299_ ;
wire _10300_ ;
wire _10301_ ;
wire _10302_ ;
wire _10303_ ;
wire _10304_ ;
wire _10305_ ;
wire _10306_ ;
wire _10307_ ;
wire _10308_ ;
wire _10309_ ;
wire _10310_ ;
wire _10311_ ;
wire _10312_ ;
wire _10313_ ;
wire _10314_ ;
wire _10315_ ;
wire _10316_ ;
wire _10317_ ;
wire _10318_ ;
wire _10319_ ;
wire _10320_ ;
wire _10321_ ;
wire _10322_ ;
wire _10323_ ;
wire _10324_ ;
wire _10325_ ;
wire _10326_ ;
wire _10327_ ;
wire _10328_ ;
wire _10329_ ;
wire _10330_ ;
wire _10331_ ;
wire _10332_ ;
wire _10333_ ;
wire _10334_ ;
wire _10335_ ;
wire _10336_ ;
wire _10337_ ;
wire _10338_ ;
wire _10339_ ;
wire _10340_ ;
wire _10341_ ;
wire _10342_ ;
wire _10343_ ;
wire _10344_ ;
wire _10345_ ;
wire _10346_ ;
wire _10347_ ;
wire _10348_ ;
wire _10349_ ;
wire _10350_ ;
wire _10351_ ;
wire _10352_ ;
wire _10353_ ;
wire _10354_ ;
wire _10355_ ;
wire _10356_ ;
wire _10357_ ;
wire _10358_ ;
wire _10359_ ;
wire _10360_ ;
wire _10361_ ;
wire _10362_ ;
wire _10363_ ;
wire _10364_ ;
wire _10365_ ;
wire _10366_ ;
wire _10367_ ;
wire _10368_ ;
wire _10369_ ;
wire _10370_ ;
wire _10371_ ;
wire _10372_ ;
wire _10373_ ;
wire _10374_ ;
wire _10375_ ;
wire _10376_ ;
wire _10377_ ;
wire _10378_ ;
wire _10379_ ;
wire _10380_ ;
wire _10381_ ;
wire _10382_ ;
wire _10383_ ;
wire _10384_ ;
wire _10385_ ;
wire _10386_ ;
wire _10387_ ;
wire _10388_ ;
wire _10389_ ;
wire _10390_ ;
wire _10391_ ;
wire _10392_ ;
wire _10393_ ;
wire _10394_ ;
wire _10395_ ;
wire _10396_ ;
wire _10397_ ;
wire _10398_ ;
wire _10399_ ;
wire _10400_ ;
wire _10401_ ;
wire _10402_ ;
wire _10403_ ;
wire _10404_ ;
wire _10405_ ;
wire _10406_ ;
wire _10407_ ;
wire _10408_ ;
wire _10409_ ;
wire _10410_ ;
wire _10411_ ;
wire _10412_ ;
wire _10413_ ;
wire _10414_ ;
wire _10415_ ;
wire _10416_ ;
wire _10417_ ;
wire _10418_ ;
wire _10419_ ;
wire _10420_ ;
wire _10421_ ;
wire _10422_ ;
wire _10423_ ;
wire _10424_ ;
wire _10425_ ;
wire _10426_ ;
wire _10427_ ;
wire _10428_ ;
wire _10429_ ;
wire _10430_ ;
wire _10431_ ;
wire _10432_ ;
wire _10433_ ;
wire _10434_ ;
wire _10435_ ;
wire _10436_ ;
wire _10437_ ;
wire _10438_ ;
wire _10439_ ;
wire _10440_ ;
wire _10441_ ;
wire _10442_ ;
wire _10443_ ;
wire _10444_ ;
wire _10445_ ;
wire _10446_ ;
wire _10447_ ;
wire _10448_ ;
wire _10449_ ;
wire _10450_ ;
wire _10451_ ;
wire _10452_ ;
wire _10453_ ;
wire _10454_ ;
wire _10455_ ;
wire _10456_ ;
wire _10457_ ;
wire _10458_ ;
wire _10459_ ;
wire _10460_ ;
wire _10461_ ;
wire _10462_ ;
wire _10463_ ;
wire _10464_ ;
wire _10465_ ;
wire _10466_ ;
wire _10467_ ;
wire _10468_ ;
wire _10469_ ;
wire _10470_ ;
wire _10471_ ;
wire _10472_ ;
wire _10473_ ;
wire _10474_ ;
wire _10475_ ;
wire _10476_ ;
wire _10477_ ;
wire _10478_ ;
wire _10479_ ;
wire _10480_ ;
wire _10481_ ;
wire _10482_ ;
wire _10483_ ;
wire _10484_ ;
wire _10485_ ;
wire _10486_ ;
wire _10487_ ;
wire _10488_ ;
wire _10489_ ;
wire _10490_ ;
wire _10491_ ;
wire _10492_ ;
wire _10493_ ;
wire _10494_ ;
wire _10495_ ;
wire _10496_ ;
wire _10497_ ;
wire _10498_ ;
wire _10499_ ;
wire _10500_ ;
wire _10501_ ;
wire _10502_ ;
wire _10503_ ;
wire _10504_ ;
wire _10505_ ;
wire _10506_ ;
wire _10507_ ;
wire _10508_ ;
wire _10509_ ;
wire _10510_ ;
wire _10511_ ;
wire _10512_ ;
wire _10513_ ;
wire _10514_ ;
wire _10515_ ;
wire _10516_ ;
wire _10517_ ;
wire _10518_ ;
wire _10519_ ;
wire _10520_ ;
wire _10521_ ;
wire _10522_ ;
wire _10523_ ;
wire _10524_ ;
wire _10525_ ;
wire _10526_ ;
wire _10527_ ;
wire _10528_ ;
wire _10529_ ;
wire _10530_ ;
wire _10531_ ;
wire _10532_ ;
wire _10533_ ;
wire _10534_ ;
wire _10535_ ;
wire _10536_ ;
wire _10537_ ;
wire _10538_ ;
wire _10539_ ;
wire _10540_ ;
wire _10541_ ;
wire _10542_ ;
wire _10543_ ;
wire _10544_ ;
wire _10545_ ;
wire _10546_ ;
wire _10547_ ;
wire _10548_ ;
wire _10549_ ;
wire _10550_ ;
wire _10551_ ;
wire _10552_ ;
wire _10553_ ;
wire _10554_ ;
wire _10555_ ;
wire _10556_ ;
wire _10557_ ;
wire _10558_ ;
wire _10559_ ;
wire _10560_ ;
wire _10561_ ;
wire _10562_ ;
wire _10563_ ;
wire _10564_ ;
wire _10565_ ;
wire _10566_ ;
wire _10567_ ;
wire _10568_ ;
wire _10569_ ;
wire _10570_ ;
wire _10571_ ;
wire _10572_ ;
wire _10573_ ;
wire _10574_ ;
wire _10575_ ;
wire _10576_ ;
wire _10577_ ;
wire _10578_ ;
wire _10579_ ;
wire _10580_ ;
wire _10581_ ;
wire _10582_ ;
wire _10583_ ;
wire _10584_ ;
wire _10585_ ;
wire _10586_ ;
wire _10587_ ;
wire _10588_ ;
wire _10589_ ;
wire _10590_ ;
wire _10591_ ;
wire _10592_ ;
wire _10593_ ;
wire _10594_ ;
wire _10595_ ;
wire _10596_ ;
wire _10597_ ;
wire _10598_ ;
wire _10599_ ;
wire _10600_ ;
wire _10601_ ;
wire _10602_ ;
wire _10603_ ;
wire _10604_ ;
wire _10605_ ;
wire _10606_ ;
wire _10607_ ;
wire _10608_ ;
wire _10609_ ;
wire _10610_ ;
wire _10611_ ;
wire _10612_ ;
wire _10613_ ;
wire _10614_ ;
wire _10615_ ;
wire _10616_ ;
wire _10617_ ;
wire _10618_ ;
wire _10619_ ;
wire _10620_ ;
wire _10621_ ;
wire _10622_ ;
wire _10623_ ;
wire _10624_ ;
wire _10625_ ;
wire _10626_ ;
wire _10627_ ;
wire _10628_ ;
wire _10629_ ;
wire _10630_ ;
wire _10631_ ;
wire _10632_ ;
wire _10633_ ;
wire _10634_ ;
wire _10635_ ;
wire _10636_ ;
wire _10637_ ;
wire _10638_ ;
wire _10639_ ;
wire _10640_ ;
wire _10641_ ;
wire _10642_ ;
wire _10643_ ;
wire _10644_ ;
wire _10645_ ;
wire _10646_ ;
wire _10647_ ;
wire _10648_ ;
wire _10649_ ;
wire _10650_ ;
wire _10651_ ;
wire _10652_ ;
wire _10653_ ;
wire _10654_ ;
wire _10655_ ;
wire _10656_ ;
wire _10657_ ;
wire _10658_ ;
wire _10659_ ;
wire _10660_ ;
wire _10661_ ;
wire _10662_ ;
wire _10663_ ;
wire _10664_ ;
wire _10665_ ;
wire _10666_ ;
wire _10667_ ;
wire _10668_ ;
wire _10669_ ;
wire _10670_ ;
wire _10671_ ;
wire _10672_ ;
wire _10673_ ;
wire _10674_ ;
wire _10675_ ;
wire _10676_ ;
wire _10677_ ;
wire _10678_ ;
wire _10679_ ;
wire _10680_ ;
wire _10681_ ;
wire _10682_ ;
wire _10683_ ;
wire _10684_ ;
wire _10685_ ;
wire _10686_ ;
wire _10687_ ;
wire _10688_ ;
wire _10689_ ;
wire _10690_ ;
wire _10691_ ;
wire _10692_ ;
wire _10693_ ;
wire _10694_ ;
wire _10695_ ;
wire _10696_ ;
wire _10697_ ;
wire _10698_ ;
wire _10699_ ;
wire _10700_ ;
wire _10701_ ;
wire _10702_ ;
wire _10703_ ;
wire _10704_ ;
wire _10705_ ;
wire _10706_ ;
wire _10707_ ;
wire _10708_ ;
wire _10709_ ;
wire _10710_ ;
wire _10711_ ;
wire _10712_ ;
wire _10713_ ;
wire _10714_ ;
wire _10715_ ;
wire _10716_ ;
wire _10717_ ;
wire _10718_ ;
wire _10719_ ;
wire _10720_ ;
wire _10721_ ;
wire _10722_ ;
wire _10723_ ;
wire _10724_ ;
wire _10725_ ;
wire _10726_ ;
wire _10727_ ;
wire _10728_ ;
wire _10729_ ;
wire _10730_ ;
wire _10731_ ;
wire _10732_ ;
wire _10733_ ;
wire _10734_ ;
wire _10735_ ;
wire _10736_ ;
wire _10737_ ;
wire _10738_ ;
wire _10739_ ;
wire _10740_ ;
wire _10741_ ;
wire _10742_ ;
wire _10743_ ;
wire _10744_ ;
wire _10745_ ;
wire _10746_ ;
wire _10747_ ;
wire _10748_ ;
wire _10749_ ;
wire _10750_ ;
wire _10751_ ;
wire _10752_ ;
wire _10753_ ;
wire _10754_ ;
wire _10755_ ;
wire _10756_ ;
wire _10757_ ;
wire _10758_ ;
wire _10759_ ;
wire _10760_ ;
wire _10761_ ;
wire _10762_ ;
wire _10763_ ;
wire _10764_ ;
wire _10765_ ;
wire _10766_ ;
wire _10767_ ;
wire _10768_ ;
wire _10769_ ;
wire _10770_ ;
wire _10771_ ;
wire _10772_ ;
wire _10773_ ;
wire _10774_ ;
wire _10775_ ;
wire _10776_ ;
wire _10777_ ;
wire _10778_ ;
wire _10779_ ;
wire _10780_ ;
wire _10781_ ;
wire _10782_ ;
wire _10783_ ;
wire _10784_ ;
wire _10785_ ;
wire _10786_ ;
wire _10787_ ;
wire _10788_ ;
wire _10789_ ;
wire _10790_ ;
wire _10791_ ;
wire _10792_ ;
wire _10793_ ;
wire _10794_ ;
wire _10795_ ;
wire _10796_ ;
wire _10797_ ;
wire _10798_ ;
wire _10799_ ;
wire _10800_ ;
wire _10801_ ;
wire _10802_ ;
wire _10803_ ;
wire _10804_ ;
wire _10805_ ;
wire _10806_ ;
wire _10807_ ;
wire _10808_ ;
wire _10809_ ;
wire _10810_ ;
wire _10811_ ;
wire _10812_ ;
wire _10813_ ;
wire _10814_ ;
wire _10815_ ;
wire _10816_ ;
wire _10817_ ;
wire _10818_ ;
wire _10819_ ;
wire _10820_ ;
wire _10821_ ;
wire _10822_ ;
wire _10823_ ;
wire _10824_ ;
wire _10825_ ;
wire _10826_ ;
wire _10827_ ;
wire _10828_ ;
wire _10829_ ;
wire _10830_ ;
wire _10831_ ;
wire _10832_ ;
wire _10833_ ;
wire _10834_ ;
wire _10835_ ;
wire _10836_ ;
wire _10837_ ;
wire _10838_ ;
wire _10839_ ;
wire _10840_ ;
wire _10841_ ;
wire _10842_ ;
wire _10843_ ;
wire _10844_ ;
wire _10845_ ;
wire _10846_ ;
wire _10847_ ;
wire _10848_ ;
wire _10849_ ;
wire _10850_ ;
wire _10851_ ;
wire _10852_ ;
wire _10853_ ;
wire _10854_ ;
wire _10855_ ;
wire _10856_ ;
wire _10857_ ;
wire _10858_ ;
wire _10859_ ;
wire _10860_ ;
wire _10861_ ;
wire _10862_ ;
wire _10863_ ;
wire _10864_ ;
wire _10865_ ;
wire _10866_ ;
wire _10867_ ;
wire _10868_ ;
wire _10869_ ;
wire _10870_ ;
wire _10871_ ;
wire _10872_ ;
wire _10873_ ;
wire _10874_ ;
wire _10875_ ;
wire _10876_ ;
wire _10877_ ;
wire _10878_ ;
wire _10879_ ;
wire _10880_ ;
wire _10881_ ;
wire _10882_ ;
wire _10883_ ;
wire _10884_ ;
wire _10885_ ;
wire _10886_ ;
wire _10887_ ;
wire _10888_ ;
wire _10889_ ;
wire _10890_ ;
wire _10891_ ;
wire _10892_ ;
wire _10893_ ;
wire _10894_ ;
wire _10895_ ;
wire _10896_ ;
wire _10897_ ;
wire _10898_ ;
wire _10899_ ;
wire _10900_ ;
wire _10901_ ;
wire _10902_ ;
wire _10903_ ;
wire _10904_ ;
wire _10905_ ;
wire _10906_ ;
wire _10907_ ;
wire _10908_ ;
wire _10909_ ;
wire _10910_ ;
wire _10911_ ;
wire _10912_ ;
wire _10913_ ;
wire _10914_ ;
wire _10915_ ;
wire _10916_ ;
wire _10917_ ;
wire _10918_ ;
wire _10919_ ;
wire _10920_ ;
wire _10921_ ;
wire _10922_ ;
wire _10923_ ;
wire _10924_ ;
wire _10925_ ;
wire _10926_ ;
wire _10927_ ;
wire _10928_ ;
wire _10929_ ;
wire _10930_ ;
wire _10931_ ;
wire _10932_ ;
wire _10933_ ;
wire _10934_ ;
wire _10935_ ;
wire _10936_ ;
wire _10937_ ;
wire _10938_ ;
wire _10939_ ;
wire _10940_ ;
wire _10941_ ;
wire _10942_ ;
wire _10943_ ;
wire _10944_ ;
wire _10945_ ;
wire _10946_ ;
wire _10947_ ;
wire _10948_ ;
wire _10949_ ;
wire _10950_ ;
wire _10951_ ;
wire _10952_ ;
wire _10953_ ;
wire _10954_ ;
wire _10955_ ;
wire _10956_ ;
wire _10957_ ;
wire _10958_ ;
wire _10959_ ;
wire _10960_ ;
wire _10961_ ;
wire _10962_ ;
wire _10963_ ;
wire _10964_ ;
wire _10965_ ;
wire _10966_ ;
wire _10967_ ;
wire _10968_ ;
wire _10969_ ;
wire _10970_ ;
wire _10971_ ;
wire _10972_ ;
wire _10973_ ;
wire _10974_ ;
wire _10975_ ;
wire _10976_ ;
wire _10977_ ;
wire _10978_ ;
wire _10979_ ;
wire _10980_ ;
wire _10981_ ;
wire _10982_ ;
wire _10983_ ;
wire _10984_ ;
wire _10985_ ;
wire _10986_ ;
wire _10987_ ;
wire _10988_ ;
wire _10989_ ;
wire _10990_ ;
wire _10991_ ;
wire _10992_ ;
wire _10993_ ;
wire _10994_ ;
wire _10995_ ;
wire _10996_ ;
wire _10997_ ;
wire _10998_ ;
wire _10999_ ;
wire _11000_ ;
wire _11001_ ;
wire _11002_ ;
wire _11003_ ;
wire _11004_ ;
wire _11005_ ;
wire _11006_ ;
wire _11007_ ;
wire _11008_ ;
wire _11009_ ;
wire _11010_ ;
wire _11011_ ;
wire _11012_ ;
wire _11013_ ;
wire _11014_ ;
wire _11015_ ;
wire _11016_ ;
wire _11017_ ;
wire _11018_ ;
wire _11019_ ;
wire _11020_ ;
wire _11021_ ;
wire _11022_ ;
wire _11023_ ;
wire _11024_ ;
wire _11025_ ;
wire _11026_ ;
wire _11027_ ;
wire _11028_ ;
wire _11029_ ;
wire _11030_ ;
wire _11031_ ;
wire _11032_ ;
wire _11033_ ;
wire _11034_ ;
wire _11035_ ;
wire _11036_ ;
wire _11037_ ;
wire _11038_ ;
wire _11039_ ;
wire _11040_ ;
wire _11041_ ;
wire _11042_ ;
wire _11043_ ;
wire _11044_ ;
wire _11045_ ;
wire _11046_ ;
wire _11047_ ;
wire _11048_ ;
wire _11049_ ;
wire _11050_ ;
wire _11051_ ;
wire _11052_ ;
wire _11053_ ;
wire _11054_ ;
wire _11055_ ;
wire _11056_ ;
wire _11057_ ;
wire _11058_ ;
wire _11059_ ;
wire _11060_ ;
wire _11061_ ;
wire _11062_ ;
wire _11063_ ;
wire _11064_ ;
wire _11065_ ;
wire _11066_ ;
wire _11067_ ;
wire _11068_ ;
wire _11069_ ;
wire _11070_ ;
wire _11071_ ;
wire _11072_ ;
wire _11073_ ;
wire _11074_ ;
wire _11075_ ;
wire _11076_ ;
wire _11077_ ;
wire _11078_ ;
wire _11079_ ;
wire _11080_ ;
wire _11081_ ;
wire _11082_ ;
wire _11083_ ;
wire _11084_ ;
wire _11085_ ;
wire _11086_ ;
wire _11087_ ;
wire _11088_ ;
wire _11089_ ;
wire _11090_ ;
wire _11091_ ;
wire _11092_ ;
wire _11093_ ;
wire _11094_ ;
wire _11095_ ;
wire _11096_ ;
wire _11097_ ;
wire _11098_ ;
wire _11099_ ;
wire _11100_ ;
wire _11101_ ;
wire _11102_ ;
wire _11103_ ;
wire _11104_ ;
wire _11105_ ;
wire _11106_ ;
wire _11107_ ;
wire _11108_ ;
wire _11109_ ;
wire _11110_ ;
wire _11111_ ;
wire _11112_ ;
wire _11113_ ;
wire _11114_ ;
wire _11115_ ;
wire _11116_ ;
wire _11117_ ;
wire _11118_ ;
wire _11119_ ;
wire _11120_ ;
wire _11121_ ;
wire _11122_ ;
wire _11123_ ;
wire _11124_ ;
wire _11125_ ;
wire _11126_ ;
wire _11127_ ;
wire _11128_ ;
wire _11129_ ;
wire _11130_ ;
wire _11131_ ;
wire _11132_ ;
wire _11133_ ;
wire _11134_ ;
wire _11135_ ;
wire _11136_ ;
wire _11137_ ;
wire _11138_ ;
wire _11139_ ;
wire _11140_ ;
wire _11141_ ;
wire _11142_ ;
wire _11143_ ;
wire _11144_ ;
wire _11145_ ;
wire _11146_ ;
wire _11147_ ;
wire _11148_ ;
wire _11149_ ;
wire _11150_ ;
wire _11151_ ;
wire _11152_ ;
wire _11153_ ;
wire _11154_ ;
wire _11155_ ;
wire _11156_ ;
wire _11157_ ;
wire _11158_ ;
wire _11159_ ;
wire _11160_ ;
wire _11161_ ;
wire _11162_ ;
wire _11163_ ;
wire _11164_ ;
wire _11165_ ;
wire _11166_ ;
wire _11167_ ;
wire _11168_ ;
wire _11169_ ;
wire _11170_ ;
wire _11171_ ;
wire _11172_ ;
wire _11173_ ;
wire _11174_ ;
wire _11175_ ;
wire _11176_ ;
wire _11177_ ;
wire _11178_ ;
wire _11179_ ;
wire _11180_ ;
wire _11181_ ;
wire _11182_ ;
wire _11183_ ;
wire _11184_ ;
wire _11185_ ;
wire _11186_ ;
wire _11187_ ;
wire _11188_ ;
wire _11189_ ;
wire _11190_ ;
wire _11191_ ;
wire _11192_ ;
wire _11193_ ;
wire _11194_ ;
wire _11195_ ;
wire _11196_ ;
wire _11197_ ;
wire _11198_ ;
wire _11199_ ;
wire _11200_ ;
wire _11201_ ;
wire _11202_ ;
wire _11203_ ;
wire _11204_ ;
wire _11205_ ;
wire _11206_ ;
wire _11207_ ;
wire _11208_ ;
wire _11209_ ;
wire _11210_ ;
wire _11211_ ;
wire _11212_ ;
wire _11213_ ;
wire _11214_ ;
wire _11215_ ;
wire _11216_ ;
wire _11217_ ;
wire _11218_ ;
wire _11219_ ;
wire _11220_ ;
wire _11221_ ;
wire _11222_ ;
wire _11223_ ;
wire _11224_ ;
wire _11225_ ;
wire _11226_ ;
wire _11227_ ;
wire _11228_ ;
wire _11229_ ;
wire _11230_ ;
wire _11231_ ;
wire _11232_ ;
wire _11233_ ;
wire _11234_ ;
wire _11235_ ;
wire _11236_ ;
wire _11237_ ;
wire _11238_ ;
wire _11239_ ;
wire _11240_ ;
wire _11241_ ;
wire _11242_ ;
wire _11243_ ;
wire _11244_ ;
wire _11245_ ;
wire _11246_ ;
wire _11247_ ;
wire _11248_ ;
wire _11249_ ;
wire _11250_ ;
wire _11251_ ;
wire _11252_ ;
wire _11253_ ;
wire _11254_ ;
wire _11255_ ;
wire _11256_ ;
wire _11257_ ;
wire _11258_ ;
wire _11259_ ;
wire _11260_ ;
wire _11261_ ;
wire _11262_ ;
wire _11263_ ;
wire _11264_ ;
wire _11265_ ;
wire _11266_ ;
wire _11267_ ;
wire _11268_ ;
wire _11269_ ;
wire _11270_ ;
wire _11271_ ;
wire _11272_ ;
wire _11273_ ;
wire _11274_ ;
wire _11275_ ;
wire _11276_ ;
wire _11277_ ;
wire _11278_ ;
wire _11279_ ;
wire _11280_ ;
wire _11281_ ;
wire _11282_ ;
wire _11283_ ;
wire _11284_ ;
wire _11285_ ;
wire _11286_ ;
wire _11287_ ;
wire _11288_ ;
wire _11289_ ;
wire _11290_ ;
wire _11291_ ;
wire _11292_ ;
wire _11293_ ;
wire _11294_ ;
wire _11295_ ;
wire _11296_ ;
wire _11297_ ;
wire _11298_ ;
wire _11299_ ;
wire _11300_ ;
wire _11301_ ;
wire _11302_ ;
wire _11303_ ;
wire _11304_ ;
wire _11305_ ;
wire _11306_ ;
wire _11307_ ;
wire _11308_ ;
wire _11309_ ;
wire _11310_ ;
wire _11311_ ;
wire _11312_ ;
wire _11313_ ;
wire _11314_ ;
wire _11315_ ;
wire _11316_ ;
wire _11317_ ;
wire _11318_ ;
wire _11319_ ;
wire _11320_ ;
wire _11321_ ;
wire _11322_ ;
wire _11323_ ;
wire _11324_ ;
wire _11325_ ;
wire _11326_ ;
wire _11327_ ;
wire _11328_ ;
wire _11329_ ;
wire _11330_ ;
wire _11331_ ;
wire _11332_ ;
wire _11333_ ;
wire _11334_ ;
wire _11335_ ;
wire _11336_ ;
wire _11337_ ;
wire _11338_ ;
wire _11339_ ;
wire _11340_ ;
wire _11341_ ;
wire _11342_ ;
wire _11343_ ;
wire _11344_ ;
wire _11345_ ;
wire _11346_ ;
wire _11347_ ;
wire _11348_ ;
wire _11349_ ;
wire _11350_ ;
wire _11351_ ;
wire _11352_ ;
wire _11353_ ;
wire _11354_ ;
wire _11355_ ;
wire _11356_ ;
wire _11357_ ;
wire _11358_ ;
wire _11359_ ;
wire _11360_ ;
wire _11361_ ;
wire _11362_ ;
wire _11363_ ;
wire _11364_ ;
wire _11365_ ;
wire _11366_ ;
wire _11367_ ;
wire _11368_ ;
wire _11369_ ;
wire _11370_ ;
wire _11371_ ;
wire _11372_ ;
wire _11373_ ;
wire _11374_ ;
wire _11375_ ;
wire _11376_ ;
wire _11377_ ;
wire _11378_ ;
wire _11379_ ;
wire _11380_ ;
wire _11381_ ;
wire _11382_ ;
wire _11383_ ;
wire _11384_ ;
wire _11385_ ;
wire _11386_ ;
wire _11387_ ;
wire _11388_ ;
wire _11389_ ;
wire _11390_ ;
wire _11391_ ;
wire _11392_ ;
wire _11393_ ;
wire _11394_ ;
wire _11395_ ;
wire _11396_ ;
wire _11397_ ;
wire _11398_ ;
wire _11399_ ;
wire _11400_ ;
wire _11401_ ;
wire _11402_ ;
wire _11403_ ;
wire _11404_ ;
wire _11405_ ;
wire _11406_ ;
wire _11407_ ;
wire _11408_ ;
wire _11409_ ;
wire _11410_ ;
wire _11411_ ;
wire _11412_ ;
wire _11413_ ;
wire _11414_ ;
wire _11415_ ;
wire _11416_ ;
wire _11417_ ;
wire _11418_ ;
wire _11419_ ;
wire _11420_ ;
wire _11421_ ;
wire _11422_ ;
wire _11423_ ;
wire _11424_ ;
wire _11425_ ;
wire _11426_ ;
wire _11427_ ;
wire _11428_ ;
wire _11429_ ;
wire _11430_ ;
wire _11431_ ;
wire _11432_ ;
wire _11433_ ;
wire _11434_ ;
wire _11435_ ;
wire _11436_ ;
wire _11437_ ;
wire _11438_ ;
wire _11439_ ;
wire _11440_ ;
wire _11441_ ;
wire _11442_ ;
wire _11443_ ;
wire _11444_ ;
wire _11445_ ;
wire _11446_ ;
wire _11447_ ;
wire _11448_ ;
wire _11449_ ;
wire _11450_ ;
wire _11451_ ;
wire _11452_ ;
wire _11453_ ;
wire _11454_ ;
wire _11455_ ;
wire _11456_ ;
wire _11457_ ;
wire _11458_ ;
wire _11459_ ;
wire _11460_ ;
wire _11461_ ;
wire _11462_ ;
wire _11463_ ;
wire _11464_ ;
wire _11465_ ;
wire _11466_ ;
wire _11467_ ;
wire _11468_ ;
wire _11469_ ;
wire _11470_ ;
wire _11471_ ;
wire _11472_ ;
wire _11473_ ;
wire _11474_ ;
wire _11475_ ;
wire _11476_ ;
wire _11477_ ;
wire _11478_ ;
wire _11479_ ;
wire _11480_ ;
wire _11481_ ;
wire _11482_ ;
wire _11483_ ;
wire _11484_ ;
wire _11485_ ;
wire _11486_ ;
wire _11487_ ;
wire _11488_ ;
wire _11489_ ;
wire _11490_ ;
wire _11491_ ;
wire _11492_ ;
wire _11493_ ;
wire _11494_ ;
wire _11495_ ;
wire _11496_ ;
wire _11497_ ;
wire _11498_ ;
wire _11499_ ;
wire _11500_ ;
wire _11501_ ;
wire _11502_ ;
wire _11503_ ;
wire _11504_ ;
wire _11505_ ;
wire _11506_ ;
wire _11507_ ;
wire _11508_ ;
wire _11509_ ;
wire _11510_ ;
wire _11511_ ;
wire _11512_ ;
wire _11513_ ;
wire _11514_ ;
wire _11515_ ;
wire _11516_ ;
wire _11517_ ;
wire _11518_ ;
wire _11519_ ;
wire _11520_ ;
wire _11521_ ;
wire _11522_ ;
wire _11523_ ;
wire _11524_ ;
wire _11525_ ;
wire _11526_ ;
wire _11527_ ;
wire _11528_ ;
wire _11529_ ;
wire _11530_ ;
wire _11531_ ;
wire _11532_ ;
wire _11533_ ;
wire _11534_ ;
wire _11535_ ;
wire _11536_ ;
wire _11537_ ;
wire _11538_ ;
wire _11539_ ;
wire _11540_ ;
wire _11541_ ;
wire _11542_ ;
wire _11543_ ;
wire _11544_ ;
wire _11545_ ;
wire _11546_ ;
wire _11547_ ;
wire _11548_ ;
wire _11549_ ;
wire _11550_ ;
wire _11551_ ;
wire _11552_ ;
wire _11553_ ;
wire _11554_ ;
wire _11555_ ;
wire _11556_ ;
wire _11557_ ;
wire _11558_ ;
wire _11559_ ;
wire _11560_ ;
wire _11561_ ;
wire _11562_ ;
wire _11563_ ;
wire _11564_ ;
wire _11565_ ;
wire _11566_ ;
wire _11567_ ;
wire _11568_ ;
wire _11569_ ;
wire _11570_ ;
wire _11571_ ;
wire _11572_ ;
wire _11573_ ;
wire _11574_ ;
wire _11575_ ;
wire _11576_ ;
wire _11577_ ;
wire _11578_ ;
wire _11579_ ;
wire _11580_ ;
wire _11581_ ;
wire _11582_ ;
wire _11583_ ;
wire _11584_ ;
wire _11585_ ;
wire _11586_ ;
wire _11587_ ;
wire _11588_ ;
wire _11589_ ;
wire _11590_ ;
wire _11591_ ;
wire _11592_ ;
wire _11593_ ;
wire _11594_ ;
wire _11595_ ;
wire _11596_ ;
wire _11597_ ;
wire _11598_ ;
wire _11599_ ;
wire _11600_ ;
wire _11601_ ;
wire _11602_ ;
wire _11603_ ;
wire _11604_ ;
wire _11605_ ;
wire _11606_ ;
wire _11607_ ;
wire _11608_ ;
wire _11609_ ;
wire _11610_ ;
wire _11611_ ;
wire _11612_ ;
wire _11613_ ;
wire _11614_ ;
wire _11615_ ;
wire _11616_ ;
wire _11617_ ;
wire _11618_ ;
wire _11619_ ;
wire _11620_ ;
wire _11621_ ;
wire _11622_ ;
wire _11623_ ;
wire _11624_ ;
wire _11625_ ;
wire _11626_ ;
wire _11627_ ;
wire _11628_ ;
wire _11629_ ;
wire _11630_ ;
wire _11631_ ;
wire _11632_ ;
wire _11633_ ;
wire _11634_ ;
wire _11635_ ;
wire _11636_ ;
wire _11637_ ;
wire _11638_ ;
wire _11639_ ;
wire _11640_ ;
wire _11641_ ;
wire _11642_ ;
wire _11643_ ;
wire _11644_ ;
wire _11645_ ;
wire _11646_ ;
wire _11647_ ;
wire _11648_ ;
wire _11649_ ;
wire _11650_ ;
wire _11651_ ;
wire _11652_ ;
wire _11653_ ;
wire _11654_ ;
wire _11655_ ;
wire _11656_ ;
wire _11657_ ;
wire _11658_ ;
wire _11659_ ;
wire _11660_ ;
wire _11661_ ;
wire _11662_ ;
wire _11663_ ;
wire _11664_ ;
wire _11665_ ;
wire _11666_ ;
wire _11667_ ;
wire _11668_ ;
wire _11669_ ;
wire _11670_ ;
wire _11671_ ;
wire _11672_ ;
wire _11673_ ;
wire _11674_ ;
wire _11675_ ;
wire _11676_ ;
wire _11677_ ;
wire _11678_ ;
wire _11679_ ;
wire _11680_ ;
wire _11681_ ;
wire _11682_ ;
wire _11683_ ;
wire _11684_ ;
wire _11685_ ;
wire _11686_ ;
wire _11687_ ;
wire _11688_ ;
wire _11689_ ;
wire _11690_ ;
wire _11691_ ;
wire _11692_ ;
wire _11693_ ;
wire _11694_ ;
wire _11695_ ;
wire _11696_ ;
wire _11697_ ;
wire _11698_ ;
wire _11699_ ;
wire _11700_ ;
wire _11701_ ;
wire _11702_ ;
wire _11703_ ;
wire _11704_ ;
wire _11705_ ;
wire _11706_ ;
wire _11707_ ;
wire _11708_ ;
wire _11709_ ;
wire _11710_ ;
wire _11711_ ;
wire _11712_ ;
wire _11713_ ;
wire _11714_ ;
wire _11715_ ;
wire _11716_ ;
wire _11717_ ;
wire _11718_ ;
wire _11719_ ;
wire _11720_ ;
wire _11721_ ;
wire _11722_ ;
wire _11723_ ;
wire _11724_ ;
wire _11725_ ;
wire _11726_ ;
wire _11727_ ;
wire _11728_ ;
wire _11729_ ;
wire _11730_ ;
wire _11731_ ;
wire _11732_ ;
wire _11733_ ;
wire _11734_ ;
wire _11735_ ;
wire _11736_ ;
wire _11737_ ;
wire _11738_ ;
wire _11739_ ;
wire _11740_ ;
wire _11741_ ;
wire _11742_ ;
wire _11743_ ;
wire _11744_ ;
wire _11745_ ;
wire _11746_ ;
wire _11747_ ;
wire _11748_ ;
wire _11749_ ;
wire _11750_ ;
wire _11751_ ;
wire _11752_ ;
wire _11753_ ;
wire _11754_ ;
wire _11755_ ;
wire _11756_ ;
wire _11757_ ;
wire _11758_ ;
wire _11759_ ;
wire _11760_ ;
wire _11761_ ;
wire _11762_ ;
wire _11763_ ;
wire _11764_ ;
wire _11765_ ;
wire _11766_ ;
wire _11767_ ;
wire _11768_ ;
wire _11769_ ;
wire _11770_ ;
wire _11771_ ;
wire _11772_ ;
wire _11773_ ;
wire _11774_ ;
wire _11775_ ;
wire _11776_ ;
wire _11777_ ;
wire _11778_ ;
wire _11779_ ;
wire _11780_ ;
wire _11781_ ;
wire _11782_ ;
wire _11783_ ;
wire _11784_ ;
wire _11785_ ;
wire _11786_ ;
wire _11787_ ;
wire _11788_ ;
wire _11789_ ;
wire _11790_ ;
wire _11791_ ;
wire _11792_ ;
wire _11793_ ;
wire _11794_ ;
wire _11795_ ;
wire _11796_ ;
wire _11797_ ;
wire _11798_ ;
wire _11799_ ;
wire _11800_ ;
wire _11801_ ;
wire _11802_ ;
wire _11803_ ;
wire _11804_ ;
wire _11805_ ;
wire _11806_ ;
wire _11807_ ;
wire _11808_ ;
wire _11809_ ;
wire _11810_ ;
wire _11811_ ;
wire _11812_ ;
wire _11813_ ;
wire _11814_ ;
wire _11815_ ;
wire _11816_ ;
wire _11817_ ;
wire _11818_ ;
wire _11819_ ;
wire _11820_ ;
wire _11821_ ;
wire _11822_ ;
wire _11823_ ;
wire _11824_ ;
wire _11825_ ;
wire _11826_ ;
wire _11827_ ;
wire _11828_ ;
wire _11829_ ;
wire _11830_ ;
wire _11831_ ;
wire _11832_ ;
wire _11833_ ;
wire _11834_ ;
wire _11835_ ;
wire _11836_ ;
wire _11837_ ;
wire _11838_ ;
wire _11839_ ;
wire _11840_ ;
wire _11841_ ;
wire _11842_ ;
wire _11843_ ;
wire _11844_ ;
wire _11845_ ;
wire _11846_ ;
wire _11847_ ;
wire _11848_ ;
wire _11849_ ;
wire _11850_ ;
wire _11851_ ;
wire _11852_ ;
wire _11853_ ;
wire _11854_ ;
wire _11855_ ;
wire _11856_ ;
wire _11857_ ;
wire _11858_ ;
wire _11859_ ;
wire _11860_ ;
wire _11861_ ;
wire _11862_ ;
wire _11863_ ;
wire _11864_ ;
wire _11865_ ;
wire _11866_ ;
wire _11867_ ;
wire _11868_ ;
wire _11869_ ;
wire _11870_ ;
wire _11871_ ;
wire _11872_ ;
wire _11873_ ;
wire _11874_ ;
wire _11875_ ;
wire _11876_ ;
wire _11877_ ;
wire _11878_ ;
wire _11879_ ;
wire _11880_ ;
wire _11881_ ;
wire _11882_ ;
wire _11883_ ;
wire _11884_ ;
wire _11885_ ;
wire _11886_ ;
wire _11887_ ;
wire _11888_ ;
wire _11889_ ;
wire _11890_ ;
wire _11891_ ;
wire _11892_ ;
wire _11893_ ;
wire _11894_ ;
wire _11895_ ;
wire _11896_ ;
wire _11897_ ;
wire _11898_ ;
wire _11899_ ;
wire _11900_ ;
wire _11901_ ;
wire _11902_ ;
wire _11903_ ;
wire _11904_ ;
wire _11905_ ;
wire _11906_ ;
wire _11907_ ;
wire _11908_ ;
wire _11909_ ;
wire _11910_ ;
wire _11911_ ;
wire _11912_ ;
wire _11913_ ;
wire _11914_ ;
wire _11915_ ;
wire _11916_ ;
wire _11917_ ;
wire _11918_ ;
wire _11919_ ;
wire _11920_ ;
wire _11921_ ;
wire _11922_ ;
wire _11923_ ;
wire _11924_ ;
wire _11925_ ;
wire _11926_ ;
wire _11927_ ;
wire _11928_ ;
wire _11929_ ;
wire _11930_ ;
wire _11931_ ;
wire _11932_ ;
wire _11933_ ;
wire _11934_ ;
wire _11935_ ;
wire _11936_ ;
wire _11937_ ;
wire _11938_ ;
wire _11939_ ;
wire _11940_ ;
wire _11941_ ;
wire _11942_ ;
wire _11943_ ;
wire _11944_ ;
wire _11945_ ;
wire _11946_ ;
wire _11947_ ;
wire _11948_ ;
wire _11949_ ;
wire _11950_ ;
wire _11951_ ;
wire _11952_ ;
wire _11953_ ;
wire _11954_ ;
wire _11955_ ;
wire _11956_ ;
wire _11957_ ;
wire _11958_ ;
wire _11959_ ;
wire _11960_ ;
wire _11961_ ;
wire _11962_ ;
wire _11963_ ;
wire _11964_ ;
wire _11965_ ;
wire _11966_ ;
wire _11967_ ;
wire _11968_ ;
wire _11969_ ;
wire _11970_ ;
wire _11971_ ;
wire _11972_ ;
wire _11973_ ;
wire _11974_ ;
wire _11975_ ;
wire _11976_ ;
wire _11977_ ;
wire _11978_ ;
wire _11979_ ;
wire _11980_ ;
wire _11981_ ;
wire _11982_ ;
wire _11983_ ;
wire _11984_ ;
wire _11985_ ;
wire _11986_ ;
wire _11987_ ;
wire _11988_ ;
wire _11989_ ;
wire _11990_ ;
wire _11991_ ;
wire _11992_ ;
wire _11993_ ;
wire _11994_ ;
wire _11995_ ;
wire _11996_ ;
wire _11997_ ;
wire _11998_ ;
wire _11999_ ;
wire _12000_ ;
wire _12001_ ;
wire _12002_ ;
wire _12003_ ;
wire _12004_ ;
wire _12005_ ;
wire _12006_ ;
wire _12007_ ;
wire _12008_ ;
wire _12009_ ;
wire _12010_ ;
wire _12011_ ;
wire _12012_ ;
wire _12013_ ;
wire _12014_ ;
wire _12015_ ;
wire _12016_ ;
wire _12017_ ;
wire _12018_ ;
wire _12019_ ;
wire _12020_ ;
wire _12021_ ;
wire _12022_ ;
wire _12023_ ;
wire _12024_ ;
wire _12025_ ;
wire _12026_ ;
wire _12027_ ;
wire _12028_ ;
wire _12029_ ;
wire _12030_ ;
wire _12031_ ;
wire _12032_ ;
wire _12033_ ;
wire _12034_ ;
wire _12035_ ;
wire _12036_ ;
wire _12037_ ;
wire _12038_ ;
wire _12039_ ;
wire _12040_ ;
wire _12041_ ;
wire _12042_ ;
wire _12043_ ;
wire _12044_ ;
wire _12045_ ;
wire _12046_ ;
wire _12047_ ;
wire _12048_ ;
wire _12049_ ;
wire _12050_ ;
wire _12051_ ;
wire _12052_ ;
wire _12053_ ;
wire _12054_ ;
wire _12055_ ;
wire _12056_ ;
wire _12057_ ;
wire _12058_ ;
wire _12059_ ;
wire _12060_ ;
wire _12061_ ;
wire _12062_ ;
wire _12063_ ;
wire _12064_ ;
wire _12065_ ;
wire _12066_ ;
wire _12067_ ;
wire _12068_ ;
wire _12069_ ;
wire _12070_ ;
wire _12071_ ;
wire _12072_ ;
wire _12073_ ;
wire _12074_ ;
wire _12075_ ;
wire _12076_ ;
wire _12077_ ;
wire _12078_ ;
wire _12079_ ;
wire _12080_ ;
wire _12081_ ;
wire _12082_ ;
wire _12083_ ;
wire _12084_ ;
wire _12085_ ;
wire _12086_ ;
wire _12087_ ;
wire _12088_ ;
wire _12089_ ;
wire _12090_ ;
wire _12091_ ;
wire _12092_ ;
wire _12093_ ;
wire _12094_ ;
wire _12095_ ;
wire _12096_ ;
wire _12097_ ;
wire _12098_ ;
wire _12099_ ;
wire _12100_ ;
wire _12101_ ;
wire _12102_ ;
wire _12103_ ;
wire _12104_ ;
wire _12105_ ;
wire _12106_ ;
wire _12107_ ;
wire _12108_ ;
wire _12109_ ;
wire _12110_ ;
wire _12111_ ;
wire _12112_ ;
wire _12113_ ;
wire _12114_ ;
wire _12115_ ;
wire _12116_ ;
wire _12117_ ;
wire _12118_ ;
wire _12119_ ;
wire _12120_ ;
wire _12121_ ;
wire _12122_ ;
wire _12123_ ;
wire _12124_ ;
wire _12125_ ;
wire _12126_ ;
wire _12127_ ;
wire _12128_ ;
wire _12129_ ;
wire _12130_ ;
wire _12131_ ;
wire _12132_ ;
wire _12133_ ;
wire _12134_ ;
wire _12135_ ;
wire _12136_ ;
wire _12137_ ;
wire _12138_ ;
wire _12139_ ;
wire _12140_ ;
wire _12141_ ;
wire _12142_ ;
wire _12143_ ;
wire _12144_ ;
wire _12145_ ;
wire _12146_ ;
wire _12147_ ;
wire _12148_ ;
wire _12149_ ;
wire _12150_ ;
wire _12151_ ;
wire _12152_ ;
wire _12153_ ;
wire _12154_ ;
wire _12155_ ;
wire _12156_ ;
wire _12157_ ;
wire _12158_ ;
wire _12159_ ;
wire _12160_ ;
wire _12161_ ;
wire _12162_ ;
wire _12163_ ;
wire _12164_ ;
wire _12165_ ;
wire _12166_ ;
wire _12167_ ;
wire _12168_ ;
wire _12169_ ;
wire _12170_ ;
wire _12171_ ;
wire _12172_ ;
wire _12173_ ;
wire _12174_ ;
wire _12175_ ;
wire _12176_ ;
wire _12177_ ;
wire _12178_ ;
wire _12179_ ;
wire _12180_ ;
wire _12181_ ;
wire _12182_ ;
wire _12183_ ;
wire _12184_ ;
wire _12185_ ;
wire _12186_ ;
wire _12187_ ;
wire _12188_ ;
wire _12189_ ;
wire _12190_ ;
wire _12191_ ;
wire _12192_ ;
wire _12193_ ;
wire _12194_ ;
wire _12195_ ;
wire _12196_ ;
wire _12197_ ;
wire _12198_ ;
wire _12199_ ;
wire _12200_ ;
wire _12201_ ;
wire _12202_ ;
wire _12203_ ;
wire _12204_ ;
wire _12205_ ;
wire _12206_ ;
wire _12207_ ;
wire _12208_ ;
wire _12209_ ;
wire _12210_ ;
wire _12211_ ;
wire _12212_ ;
wire _12213_ ;
wire _12214_ ;
wire _12215_ ;
wire _12216_ ;
wire _12217_ ;
wire _12218_ ;
wire _12219_ ;
wire _12220_ ;
wire _12221_ ;
wire _12222_ ;
wire _12223_ ;
wire _12224_ ;
wire _12225_ ;
wire _12226_ ;
wire _12227_ ;
wire _12228_ ;
wire _12229_ ;
wire _12230_ ;
wire _12231_ ;
wire _12232_ ;
wire _12233_ ;
wire _12234_ ;
wire _12235_ ;
wire _12236_ ;
wire _12237_ ;
wire _12238_ ;
wire _12239_ ;
wire _12240_ ;
wire _12241_ ;
wire _12242_ ;
wire _12243_ ;
wire _12244_ ;
wire _12245_ ;
wire _12246_ ;
wire _12247_ ;
wire _12248_ ;
wire _12249_ ;
wire _12250_ ;
wire _12251_ ;
wire _12252_ ;
wire _12253_ ;
wire _12254_ ;
wire _12255_ ;
wire _12256_ ;
wire _12257_ ;
wire _12258_ ;
wire _12259_ ;
wire _12260_ ;
wire _12261_ ;
wire _12262_ ;
wire _12263_ ;
wire _12264_ ;
wire _12265_ ;
wire _12266_ ;
wire _12267_ ;
wire _12268_ ;
wire _12269_ ;
wire _12270_ ;
wire _12271_ ;
wire _12272_ ;
wire _12273_ ;
wire _12274_ ;
wire _12275_ ;
wire _12276_ ;
wire _12277_ ;
wire _12278_ ;
wire _12279_ ;
wire _12280_ ;
wire _12281_ ;
wire _12282_ ;
wire _12283_ ;
wire _12284_ ;
wire _12285_ ;
wire _12286_ ;
wire _12287_ ;
wire _12288_ ;
wire _12289_ ;
wire _12290_ ;
wire _12291_ ;
wire _12292_ ;
wire _12293_ ;
wire _12294_ ;
wire _12295_ ;
wire _12296_ ;
wire _12297_ ;
wire _12298_ ;
wire _12299_ ;
wire _12300_ ;
wire _12301_ ;
wire _12302_ ;
wire _12303_ ;
wire _12304_ ;
wire _12305_ ;
wire _12306_ ;
wire _12307_ ;
wire _12308_ ;
wire _12309_ ;
wire _12310_ ;
wire _12311_ ;
wire _12312_ ;
wire _12313_ ;
wire _12314_ ;
wire _12315_ ;
wire _12316_ ;
wire _12317_ ;
wire _12318_ ;
wire _12319_ ;
wire _12320_ ;
wire _12321_ ;
wire _12322_ ;
wire _12323_ ;
wire _12324_ ;
wire _12325_ ;
wire _12326_ ;
wire _12327_ ;
wire _12328_ ;
wire _12329_ ;
wire _12330_ ;
wire _12331_ ;
wire _12332_ ;
wire _12333_ ;
wire _12334_ ;
wire _12335_ ;
wire _12336_ ;
wire _12337_ ;
wire _12338_ ;
wire _12339_ ;
wire _12340_ ;
wire _12341_ ;
wire _12342_ ;
wire _12343_ ;
wire _12344_ ;
wire _12345_ ;
wire _12346_ ;
wire _12347_ ;
wire _12348_ ;
wire _12349_ ;
wire _12350_ ;
wire _12351_ ;
wire _12352_ ;
wire _12353_ ;
wire _12354_ ;
wire _12355_ ;
wire _12356_ ;
wire _12357_ ;
wire _12358_ ;
wire _12359_ ;
wire _12360_ ;
wire _12361_ ;
wire _12362_ ;
wire _12363_ ;
wire _12364_ ;
wire _12365_ ;
wire _12366_ ;
wire _12367_ ;
wire _12368_ ;
wire _12369_ ;
wire _12370_ ;
wire _12371_ ;
wire _12372_ ;
wire _12373_ ;
wire _12374_ ;
wire _12375_ ;
wire _12376_ ;
wire _12377_ ;
wire _12378_ ;
wire _12379_ ;
wire _12380_ ;
wire _12381_ ;
wire _12382_ ;
wire _12383_ ;
wire _12384_ ;
wire _12385_ ;
wire _12386_ ;
wire _12387_ ;
wire _12388_ ;
wire _12389_ ;
wire _12390_ ;
wire _12391_ ;
wire _12392_ ;
wire _12393_ ;
wire _12394_ ;
wire _12395_ ;
wire _12396_ ;
wire _12397_ ;
wire _12398_ ;
wire _12399_ ;
wire _12400_ ;
wire _12401_ ;
wire _12402_ ;
wire _12403_ ;
wire _12404_ ;
wire _12405_ ;
wire _12406_ ;
wire _12407_ ;
wire _12408_ ;
wire _12409_ ;
wire _12410_ ;
wire _12411_ ;
wire _12412_ ;
wire _12413_ ;
wire _12414_ ;
wire _12415_ ;
wire _12416_ ;
wire _12417_ ;
wire _12418_ ;
wire _12419_ ;
wire _12420_ ;
wire _12421_ ;
wire _12422_ ;
wire _12423_ ;
wire _12424_ ;
wire _12425_ ;
wire _12426_ ;
wire _12427_ ;
wire _12428_ ;
wire _12429_ ;
wire _12430_ ;
wire _12431_ ;
wire _12432_ ;
wire _12433_ ;
wire _12434_ ;
wire _12435_ ;
wire _12436_ ;
wire _12437_ ;
wire _12438_ ;
wire _12439_ ;
wire _12440_ ;
wire _12441_ ;
wire _12442_ ;
wire _12443_ ;
wire _12444_ ;
wire _12445_ ;
wire _12446_ ;
wire _12447_ ;
wire _12448_ ;
wire _12449_ ;
wire _12450_ ;
wire _12451_ ;
wire _12452_ ;
wire _12453_ ;
wire _12454_ ;
wire _12455_ ;
wire _12456_ ;
wire _12457_ ;
wire _12458_ ;
wire _12459_ ;
wire _12460_ ;
wire _12461_ ;
wire _12462_ ;
wire _12463_ ;
wire _12464_ ;
wire _12465_ ;
wire _12466_ ;
wire _12467_ ;
wire _12468_ ;
wire _12469_ ;
wire _12470_ ;
wire _12471_ ;
wire _12472_ ;
wire _12473_ ;
wire _12474_ ;
wire _12475_ ;
wire _12476_ ;
wire _12477_ ;
wire _12478_ ;
wire _12479_ ;
wire _12480_ ;
wire _12481_ ;
wire _12482_ ;
wire _12483_ ;
wire _12484_ ;
wire _12485_ ;
wire _12486_ ;
wire _12487_ ;
wire _12488_ ;
wire _12489_ ;
wire _12490_ ;
wire _12491_ ;
wire _12492_ ;
wire _12493_ ;
wire _12494_ ;
wire _12495_ ;
wire _12496_ ;
wire _12497_ ;
wire _12498_ ;
wire _12499_ ;
wire _12500_ ;
wire _12501_ ;
wire _12502_ ;
wire _12503_ ;
wire _12504_ ;
wire _12505_ ;
wire _12506_ ;
wire _12507_ ;
wire _12508_ ;
wire _12509_ ;
wire _12510_ ;
wire _12511_ ;
wire _12512_ ;
wire _12513_ ;
wire _12514_ ;
wire _12515_ ;
wire _12516_ ;
wire _12517_ ;
wire _12518_ ;
wire _12519_ ;
wire _12520_ ;
wire _12521_ ;
wire _12522_ ;
wire _12523_ ;
wire _12524_ ;
wire _12525_ ;
wire _12526_ ;
wire _12527_ ;
wire _12528_ ;
wire _12529_ ;
wire _12530_ ;
wire _12531_ ;
wire _12532_ ;
wire _12533_ ;
wire _12534_ ;
wire _12535_ ;
wire _12536_ ;
wire _12537_ ;
wire _12538_ ;
wire _12539_ ;
wire _12540_ ;
wire _12541_ ;
wire _12542_ ;
wire _12543_ ;
wire _12544_ ;
wire _12545_ ;
wire _12546_ ;
wire _12547_ ;
wire _12548_ ;
wire _12549_ ;
wire _12550_ ;
wire _12551_ ;
wire _12552_ ;
wire _12553_ ;
wire _12554_ ;
wire _12555_ ;
wire _12556_ ;
wire _12557_ ;
wire _12558_ ;
wire _12559_ ;
wire _12560_ ;
wire _12561_ ;
wire _12562_ ;
wire _12563_ ;
wire _12564_ ;
wire _12565_ ;
wire _12566_ ;
wire _12567_ ;
wire _12568_ ;
wire _12569_ ;
wire _12570_ ;
wire _12571_ ;
wire _12572_ ;
wire _12573_ ;
wire _12574_ ;
wire _12575_ ;
wire _12576_ ;
wire _12577_ ;
wire _12578_ ;
wire _12579_ ;
wire _12580_ ;
wire _12581_ ;
wire _12582_ ;
wire _12583_ ;
wire _12584_ ;
wire _12585_ ;
wire _12586_ ;
wire _12587_ ;
wire _12588_ ;
wire _12589_ ;
wire _12590_ ;
wire _12591_ ;
wire _12592_ ;
wire _12593_ ;
wire _12594_ ;
wire _12595_ ;
wire _12596_ ;
wire _12597_ ;
wire _12598_ ;
wire _12599_ ;
wire _12600_ ;
wire _12601_ ;
wire _12602_ ;
wire _12603_ ;
wire _12604_ ;
wire _12605_ ;
wire _12606_ ;
wire _12607_ ;
wire _12608_ ;
wire _12609_ ;
wire _12610_ ;
wire _12611_ ;
wire _12612_ ;
wire _12613_ ;
wire _12614_ ;
wire _12615_ ;
wire _12616_ ;
wire _12617_ ;
wire _12618_ ;
wire _12619_ ;
wire _12620_ ;
wire _12621_ ;
wire _12622_ ;
wire _12623_ ;
wire _12624_ ;
wire _12625_ ;
wire _12626_ ;
wire _12627_ ;
wire _12628_ ;
wire _12629_ ;
wire _12630_ ;
wire _12631_ ;
wire _12632_ ;
wire _12633_ ;
wire _12634_ ;
wire _12635_ ;
wire _12636_ ;
wire _12637_ ;
wire _12638_ ;
wire _12639_ ;
wire _12640_ ;
wire _12641_ ;
wire _12642_ ;
wire _12643_ ;
wire _12644_ ;
wire _12645_ ;
wire _12646_ ;
wire _12647_ ;
wire _12648_ ;
wire _12649_ ;
wire _12650_ ;
wire _12651_ ;
wire _12652_ ;
wire _12653_ ;
wire _12654_ ;
wire _12655_ ;
wire _12656_ ;
wire _12657_ ;
wire _12658_ ;
wire _12659_ ;
wire _12660_ ;
wire _12661_ ;
wire _12662_ ;
wire _12663_ ;
wire _12664_ ;
wire _12665_ ;
wire _12666_ ;
wire _12667_ ;
wire _12668_ ;
wire _12669_ ;
wire _12670_ ;
wire _12671_ ;
wire _12672_ ;
wire _12673_ ;
wire _12674_ ;
wire _12675_ ;
wire _12676_ ;
wire _12677_ ;
wire _12678_ ;
wire _12679_ ;
wire _12680_ ;
wire _12681_ ;
wire _12682_ ;
wire _12683_ ;
wire _12684_ ;
wire _12685_ ;
wire _12686_ ;
wire _12687_ ;
wire _12688_ ;
wire _12689_ ;
wire _12690_ ;
wire _12691_ ;
wire _12692_ ;
wire _12693_ ;
wire _12694_ ;
wire _12695_ ;
wire _12696_ ;
wire _12697_ ;
wire _12698_ ;
wire _12699_ ;
wire _12700_ ;
wire _12701_ ;
wire _12702_ ;
wire _12703_ ;
wire _12704_ ;
wire _12705_ ;
wire _12706_ ;
wire _12707_ ;
wire _12708_ ;
wire _12709_ ;
wire _12710_ ;
wire _12711_ ;
wire _12712_ ;
wire _12713_ ;
wire _12714_ ;
wire _12715_ ;
wire _12716_ ;
wire _12717_ ;
wire _12718_ ;
wire _12719_ ;
wire _12720_ ;
wire _12721_ ;
wire _12722_ ;
wire _12723_ ;
wire _12724_ ;
wire _12725_ ;
wire _12726_ ;
wire _12727_ ;
wire _12728_ ;
wire _12729_ ;
wire _12730_ ;
wire _12731_ ;
wire _12732_ ;
wire _12733_ ;
wire _12734_ ;
wire _12735_ ;
wire _12736_ ;
wire _12737_ ;
wire _12738_ ;
wire _12739_ ;
wire _12740_ ;
wire _12741_ ;
wire _12742_ ;
wire _12743_ ;
wire _12744_ ;
wire _12745_ ;
wire _12746_ ;
wire _12747_ ;
wire _12748_ ;
wire _12749_ ;
wire _12750_ ;
wire _12751_ ;
wire _12752_ ;
wire _12753_ ;
wire _12754_ ;
wire _12755_ ;
wire _12756_ ;
wire _12757_ ;
wire _12758_ ;
wire _12759_ ;
wire _12760_ ;
wire _12761_ ;
wire _12762_ ;
wire _12763_ ;
wire _12764_ ;
wire _12765_ ;
wire _12766_ ;
wire _12767_ ;
wire _12768_ ;
wire _12769_ ;
wire _12770_ ;
wire _12771_ ;
wire _12772_ ;
wire _12773_ ;
wire _12774_ ;
wire _12775_ ;
wire _12776_ ;
wire _12777_ ;
wire _12778_ ;
wire _12779_ ;
wire _12780_ ;
wire _12781_ ;
wire _12782_ ;
wire _12783_ ;
wire _12784_ ;
wire _12785_ ;
wire _12786_ ;
wire _12787_ ;
wire _12788_ ;
wire _12789_ ;
wire _12790_ ;
wire _12791_ ;
wire _12792_ ;
wire _12793_ ;
wire _12794_ ;
wire _12795_ ;
wire _12796_ ;
wire _12797_ ;
wire _12798_ ;
wire _12799_ ;
wire _12800_ ;
wire _12801_ ;
wire _12802_ ;
wire _12803_ ;
wire _12804_ ;
wire _12805_ ;
wire _12806_ ;
wire _12807_ ;
wire _12808_ ;
wire _12809_ ;
wire _12810_ ;
wire _12811_ ;
wire _12812_ ;
wire _12813_ ;
wire _12814_ ;
wire _12815_ ;
wire _12816_ ;
wire _12817_ ;
wire _12818_ ;
wire _12819_ ;
wire _12820_ ;
wire _12821_ ;
wire _12822_ ;
wire _12823_ ;
wire _12824_ ;
wire _12825_ ;
wire _12826_ ;
wire _12827_ ;
wire _12828_ ;
wire _12829_ ;
wire _12830_ ;
wire _12831_ ;
wire _12832_ ;
wire _12833_ ;
wire _12834_ ;
wire _12835_ ;
wire _12836_ ;
wire _12837_ ;
wire _12838_ ;
wire _12839_ ;
wire _12840_ ;
wire _12841_ ;
wire _12842_ ;
wire _12843_ ;
wire _12844_ ;
wire _12845_ ;
wire _12846_ ;
wire _12847_ ;
wire _12848_ ;
wire _12849_ ;
wire _12850_ ;
wire _12851_ ;
wire _12852_ ;
wire _12853_ ;
wire _12854_ ;
wire _12855_ ;
wire _12856_ ;
wire _12857_ ;
wire _12858_ ;
wire _12859_ ;
wire _12860_ ;
wire _12861_ ;
wire _12862_ ;
wire _12863_ ;
wire _12864_ ;
wire _12865_ ;
wire _12866_ ;
wire _12867_ ;
wire _12868_ ;
wire _12869_ ;
wire _12870_ ;
wire _12871_ ;
wire _12872_ ;
wire _12873_ ;
wire _12874_ ;
wire _12875_ ;
wire _12876_ ;
wire _12877_ ;
wire _12878_ ;
wire _12879_ ;
wire _12880_ ;
wire _12881_ ;
wire _12882_ ;
wire _12883_ ;
wire _12884_ ;
wire _12885_ ;
wire _12886_ ;
wire _12887_ ;
wire _12888_ ;
wire _12889_ ;
wire _12890_ ;
wire _12891_ ;
wire _12892_ ;
wire _12893_ ;
wire _12894_ ;
wire _12895_ ;
wire _12896_ ;
wire _12897_ ;
wire _12898_ ;
wire _12899_ ;
wire _12900_ ;
wire _12901_ ;
wire _12902_ ;
wire _12903_ ;
wire _12904_ ;
wire _12905_ ;
wire _12906_ ;
wire _12907_ ;
wire _12908_ ;
wire _12909_ ;
wire _12910_ ;
wire _12911_ ;
wire _12912_ ;
wire _12913_ ;
wire _12914_ ;
wire _12915_ ;
wire _12916_ ;
wire _12917_ ;
wire _12918_ ;
wire _12919_ ;
wire _12920_ ;
wire _12921_ ;
wire _12922_ ;
wire _12923_ ;
wire _12924_ ;
wire _12925_ ;
wire _12926_ ;
wire _12927_ ;
wire _12928_ ;
wire _12929_ ;
wire _12930_ ;
wire _12931_ ;
wire _12932_ ;
wire _12933_ ;
wire _12934_ ;
wire _12935_ ;
wire _12936_ ;
wire _12937_ ;
wire _12938_ ;
wire _12939_ ;
wire _12940_ ;
wire _12941_ ;
wire _12942_ ;
wire _12943_ ;
wire _12944_ ;
wire _12945_ ;
wire _12946_ ;
wire _12947_ ;
wire _12948_ ;
wire _12949_ ;
wire _12950_ ;
wire _12951_ ;
wire _12952_ ;
wire _12953_ ;
wire _12954_ ;
wire _12955_ ;
wire _12956_ ;
wire _12957_ ;
wire _12958_ ;
wire _12959_ ;
wire _12960_ ;
wire _12961_ ;
wire _12962_ ;
wire _12963_ ;
wire _12964_ ;
wire _12965_ ;
wire _12966_ ;
wire _12967_ ;
wire _12968_ ;
wire _12969_ ;
wire _12970_ ;
wire _12971_ ;
wire _12972_ ;
wire _12973_ ;
wire _12974_ ;
wire _12975_ ;
wire _12976_ ;
wire _12977_ ;
wire _12978_ ;
wire _12979_ ;
wire _12980_ ;
wire _12981_ ;
wire _12982_ ;
wire _12983_ ;
wire _12984_ ;
wire _12985_ ;
wire _12986_ ;
wire _12987_ ;
wire _12988_ ;
wire _12989_ ;
wire _12990_ ;
wire _12991_ ;
wire _12992_ ;
wire _12993_ ;
wire _12994_ ;
wire _12995_ ;
wire _12996_ ;
wire _12997_ ;
wire _12998_ ;
wire _12999_ ;
wire _13000_ ;
wire _13001_ ;
wire _13002_ ;
wire _13003_ ;
wire _13004_ ;
wire _13005_ ;
wire _13006_ ;
wire _13007_ ;
wire _13008_ ;
wire _13009_ ;
wire _13010_ ;
wire _13011_ ;
wire _13012_ ;
wire _13013_ ;
wire _13014_ ;
wire _13015_ ;
wire _13016_ ;
wire _13017_ ;
wire _13018_ ;
wire _13019_ ;
wire _13020_ ;
wire _13021_ ;
wire _13022_ ;
wire _13023_ ;
wire _13024_ ;
wire _13025_ ;
wire _13026_ ;
wire _13027_ ;
wire _13028_ ;
wire _13029_ ;
wire _13030_ ;
wire _13031_ ;
wire _13032_ ;
wire _13033_ ;
wire _13034_ ;
wire _13035_ ;
wire _13036_ ;
wire _13037_ ;
wire _13038_ ;
wire _13039_ ;
wire _13040_ ;
wire _13041_ ;
wire _13042_ ;
wire _13043_ ;
wire _13044_ ;
wire _13045_ ;
wire _13046_ ;
wire _13047_ ;
wire _13048_ ;
wire _13049_ ;
wire _13050_ ;
wire _13051_ ;
wire _13052_ ;
wire _13053_ ;
wire _13054_ ;
wire _13055_ ;
wire _13056_ ;
wire _13057_ ;
wire _13058_ ;
wire _13059_ ;
wire _13060_ ;
wire _13061_ ;
wire _13062_ ;
wire _13063_ ;
wire _13064_ ;
wire _13065_ ;
wire _13066_ ;
wire _13067_ ;
wire _13068_ ;
wire _13069_ ;
wire _13070_ ;
wire _13071_ ;
wire _13072_ ;
wire _13073_ ;
wire _13074_ ;
wire _13075_ ;
wire _13076_ ;
wire _13077_ ;
wire _13078_ ;
wire _13079_ ;
wire _13080_ ;
wire _13081_ ;
wire _13082_ ;
wire _13083_ ;
wire _13084_ ;
wire _13085_ ;
wire _13086_ ;
wire _13087_ ;
wire _13088_ ;
wire _13089_ ;
wire _13090_ ;
wire _13091_ ;
wire _13092_ ;
wire _13093_ ;
wire _13094_ ;
wire _13095_ ;
wire _13096_ ;
wire _13097_ ;
wire _13098_ ;
wire _13099_ ;
wire _13100_ ;
wire _13101_ ;
wire _13102_ ;
wire _13103_ ;
wire _13104_ ;
wire _13105_ ;
wire _13106_ ;
wire _13107_ ;
wire _13108_ ;
wire _13109_ ;
wire _13110_ ;
wire _13111_ ;
wire _13112_ ;
wire _13113_ ;
wire _13114_ ;
wire _13115_ ;
wire _13116_ ;
wire _13117_ ;
wire _13118_ ;
wire _13119_ ;
wire _13120_ ;
wire _13121_ ;
wire _13122_ ;
wire _13123_ ;
wire _13124_ ;
wire _13125_ ;
wire _13126_ ;
wire _13127_ ;
wire _13128_ ;
wire _13129_ ;
wire _13130_ ;
wire _13131_ ;
wire _13132_ ;
wire _13133_ ;
wire _13134_ ;
wire _13135_ ;
wire _13136_ ;
wire _13137_ ;
wire _13138_ ;
wire _13139_ ;
wire _13140_ ;
wire _13141_ ;
wire _13142_ ;
wire _13143_ ;
wire _13144_ ;
wire _13145_ ;
wire _13146_ ;
wire _13147_ ;
wire _13148_ ;
wire _13149_ ;
wire _13150_ ;
wire _13151_ ;
wire _13152_ ;
wire _13153_ ;
wire _13154_ ;
wire _13155_ ;
wire _13156_ ;
wire _13157_ ;
wire _13158_ ;
wire _13159_ ;
wire _13160_ ;
wire _13161_ ;
wire _13162_ ;
wire _13163_ ;
wire _13164_ ;
wire _13165_ ;
wire _13166_ ;
wire _13167_ ;
wire _13168_ ;
wire _13169_ ;
wire _13170_ ;
wire _13171_ ;
wire _13172_ ;
wire _13173_ ;
wire _13174_ ;
wire _13175_ ;
wire _13176_ ;
wire _13177_ ;
wire _13178_ ;
wire _13179_ ;
wire _13180_ ;
wire _13181_ ;
wire _13182_ ;
wire _13183_ ;
wire _13184_ ;
wire _13185_ ;
wire _13186_ ;
wire _13187_ ;
wire _13188_ ;
wire _13189_ ;
wire _13190_ ;
wire _13191_ ;
wire _13192_ ;
wire _13193_ ;
wire _13194_ ;
wire _13195_ ;
wire _13196_ ;
wire _13197_ ;
wire _13198_ ;
wire _13199_ ;
wire _13200_ ;
wire _13201_ ;
wire _13202_ ;
wire _13203_ ;
wire _13204_ ;
wire _13205_ ;
wire _13206_ ;
wire _13207_ ;
wire _13208_ ;
wire _13209_ ;
wire _13210_ ;
wire _13211_ ;
wire _13212_ ;
wire _13213_ ;
wire _13214_ ;
wire _13215_ ;
wire _13216_ ;
wire _13217_ ;
wire _13218_ ;
wire _13219_ ;
wire _13220_ ;
wire _13221_ ;
wire _13222_ ;
wire _13223_ ;
wire _13224_ ;
wire _13225_ ;
wire _13226_ ;
wire _13227_ ;
wire _13228_ ;
wire _13229_ ;
wire _13230_ ;
wire _13231_ ;
wire _13232_ ;
wire _13233_ ;
wire _13234_ ;
wire _13235_ ;
wire _13236_ ;
wire _13237_ ;
wire _13238_ ;
wire _13239_ ;
wire _13240_ ;
wire _13241_ ;
wire _13242_ ;
wire _13243_ ;
wire _13244_ ;
wire _13245_ ;
wire _13246_ ;
wire _13247_ ;
wire _13248_ ;
wire _13249_ ;
wire _13250_ ;
wire _13251_ ;
wire _13252_ ;
wire _13253_ ;
wire _13254_ ;
wire _13255_ ;
wire _13256_ ;
wire _13257_ ;
wire _13258_ ;
wire _13259_ ;
wire _13260_ ;
wire _13261_ ;
wire _13262_ ;
wire _13263_ ;
wire _13264_ ;
wire _13265_ ;
wire _13266_ ;
wire _13267_ ;
wire _13268_ ;
wire _13269_ ;
wire _13270_ ;
wire _13271_ ;
wire _13272_ ;
wire _13273_ ;
wire _13274_ ;
wire _13275_ ;
wire _13276_ ;
wire _13277_ ;
wire _13278_ ;
wire _13279_ ;
wire _13280_ ;
wire _13281_ ;
wire _13282_ ;
wire _13283_ ;
wire _13284_ ;
wire _13285_ ;
wire _13286_ ;
wire _13287_ ;
wire _13288_ ;
wire _13289_ ;
wire _13290_ ;
wire _13291_ ;
wire _13292_ ;
wire _13293_ ;
wire _13294_ ;
wire _13295_ ;
wire _13296_ ;
wire _13297_ ;
wire _13298_ ;
wire _13299_ ;
wire _13300_ ;
wire _13301_ ;
wire _13302_ ;
wire _13303_ ;
wire _13304_ ;
wire _13305_ ;
wire _13306_ ;
wire _13307_ ;
wire _13308_ ;
wire _13309_ ;
wire _13310_ ;
wire _13311_ ;
wire _13312_ ;
wire _13313_ ;
wire _13314_ ;
wire _13315_ ;
wire _13316_ ;
wire _13317_ ;
wire _13318_ ;
wire _13319_ ;
wire _13320_ ;
wire _13321_ ;
wire _13322_ ;
wire _13323_ ;
wire _13324_ ;
wire _13325_ ;
wire _13326_ ;
wire _13327_ ;
wire _13328_ ;
wire _13329_ ;
wire _13330_ ;
wire _13331_ ;
wire _13332_ ;
wire _13333_ ;
wire _13334_ ;
wire _13335_ ;
wire _13336_ ;
wire _13337_ ;
wire _13338_ ;
wire _13339_ ;
wire _13340_ ;
wire _13341_ ;
wire _13342_ ;
wire _13343_ ;
wire _13344_ ;
wire _13345_ ;
wire _13346_ ;
wire _13347_ ;
wire _13348_ ;
wire _13349_ ;
wire _13350_ ;
wire _13351_ ;
wire _13352_ ;
wire _13353_ ;
wire _13354_ ;
wire _13355_ ;
wire _13356_ ;
wire _13357_ ;
wire _13358_ ;
wire _13359_ ;
wire _13360_ ;
wire _13361_ ;
wire _13362_ ;
wire _13363_ ;
wire _13364_ ;
wire _13365_ ;
wire _13366_ ;
wire _13367_ ;
wire _13368_ ;
wire _13369_ ;
wire _13370_ ;
wire _13371_ ;
wire _13372_ ;
wire _13373_ ;
wire _13374_ ;
wire _13375_ ;
wire _13376_ ;
wire _13377_ ;
wire _13378_ ;
wire _13379_ ;
wire _13380_ ;
wire _13381_ ;
wire _13382_ ;
wire _13383_ ;
wire _13384_ ;
wire _13385_ ;
wire _13386_ ;
wire _13387_ ;
wire _13388_ ;
wire _13389_ ;
wire _13390_ ;
wire _13391_ ;
wire _13392_ ;
wire _13393_ ;
wire _13394_ ;
wire _13395_ ;
wire _13396_ ;
wire _13397_ ;
wire _13398_ ;
wire _13399_ ;
wire _13400_ ;
wire _13401_ ;
wire _13402_ ;
wire _13403_ ;
wire _13404_ ;
wire _13405_ ;
wire _13406_ ;
wire _13407_ ;
wire _13408_ ;
wire _13409_ ;
wire _13410_ ;
wire _13411_ ;
wire _13412_ ;
wire _13413_ ;
wire _13414_ ;
wire _13415_ ;
wire _13416_ ;
wire _13417_ ;
wire _13418_ ;
wire _13419_ ;
wire _13420_ ;
wire _13421_ ;
wire _13422_ ;
wire _13423_ ;
wire _13424_ ;
wire _13425_ ;
wire _13426_ ;
wire _13427_ ;
wire _13428_ ;
wire _13429_ ;
wire _13430_ ;
wire _13431_ ;
wire _13432_ ;
wire _13433_ ;
wire _13434_ ;
wire _13435_ ;
wire _13436_ ;
wire _13437_ ;
wire _13438_ ;
wire _13439_ ;
wire _13440_ ;
wire _13441_ ;
wire _13442_ ;
wire _13443_ ;
wire _13444_ ;
wire _13445_ ;
wire _13446_ ;
wire _13447_ ;
wire _13448_ ;
wire _13449_ ;
wire _13450_ ;
wire _13451_ ;
wire _13452_ ;
wire _13453_ ;
wire _13454_ ;
wire _13455_ ;
wire _13456_ ;
wire _13457_ ;
wire _13458_ ;
wire _13459_ ;
wire _13460_ ;
wire _13461_ ;
wire _13462_ ;
wire _13463_ ;
wire _13464_ ;
wire _13465_ ;
wire _13466_ ;
wire _13467_ ;
wire _13468_ ;
wire _13469_ ;
wire _13470_ ;
wire _13471_ ;
wire _13472_ ;
wire _13473_ ;
wire _13474_ ;
wire _13475_ ;
wire _13476_ ;
wire _13477_ ;
wire _13478_ ;
wire _13479_ ;
wire _13480_ ;
wire _13481_ ;
wire _13482_ ;
wire _13483_ ;
wire _13484_ ;
wire _13485_ ;
wire _13486_ ;
wire _13487_ ;
wire _13488_ ;
wire _13489_ ;
wire _13490_ ;
wire _13491_ ;
wire _13492_ ;
wire _13493_ ;
wire _13494_ ;
wire _13495_ ;
wire _13496_ ;
wire _13497_ ;
wire _13498_ ;
wire _13499_ ;
wire _13500_ ;
wire _13501_ ;
wire _13502_ ;
wire _13503_ ;
wire _13504_ ;
wire _13505_ ;
wire _13506_ ;
wire _13507_ ;
wire _13508_ ;
wire _13509_ ;
wire _13510_ ;
wire _13511_ ;
wire _13512_ ;
wire _13513_ ;
wire _13514_ ;
wire _13515_ ;
wire _13516_ ;
wire _13517_ ;
wire _13518_ ;
wire _13519_ ;
wire _13520_ ;
wire _13521_ ;
wire _13522_ ;
wire _13523_ ;
wire _13524_ ;
wire _13525_ ;
wire _13526_ ;
wire _13527_ ;
wire _13528_ ;
wire _13529_ ;
wire _13530_ ;
wire _13531_ ;
wire _13532_ ;
wire _13533_ ;
wire _13534_ ;
wire _13535_ ;
wire _13536_ ;
wire _13537_ ;
wire _13538_ ;
wire _13539_ ;
wire _13540_ ;
wire _13541_ ;
wire _13542_ ;
wire _13543_ ;
wire _13544_ ;
wire _13545_ ;
wire _13546_ ;
wire _13547_ ;
wire _13548_ ;
wire _13549_ ;
wire _13550_ ;
wire _13551_ ;
wire _13552_ ;
wire _13553_ ;
wire _13554_ ;
wire _13555_ ;
wire _13556_ ;
wire _13557_ ;
wire _13558_ ;
wire _13559_ ;
wire _13560_ ;
wire _13561_ ;
wire _13562_ ;
wire _13563_ ;
wire _13564_ ;
wire _13565_ ;
wire _13566_ ;
wire _13567_ ;
wire _13568_ ;
wire _13569_ ;
wire _13570_ ;
wire _13571_ ;
wire _13572_ ;
wire _13573_ ;
wire _13574_ ;
wire _13575_ ;
wire _13576_ ;
wire _13577_ ;
wire _13578_ ;
wire _13579_ ;
wire _13580_ ;
wire _13581_ ;
wire _13582_ ;
wire _13583_ ;
wire _13584_ ;
wire _13585_ ;
wire _13586_ ;
wire _13587_ ;
wire _13588_ ;
wire _13589_ ;
wire _13590_ ;
wire _13591_ ;
wire _13592_ ;
wire _13593_ ;
wire _13594_ ;
wire _13595_ ;
wire _13596_ ;
wire _13597_ ;
wire _13598_ ;
wire _13599_ ;
wire _13600_ ;
wire _13601_ ;
wire _13602_ ;
wire _13603_ ;
wire _13604_ ;
wire _13605_ ;
wire _13606_ ;
wire _13607_ ;
wire _13608_ ;
wire _13609_ ;
wire _13610_ ;
wire _13611_ ;
wire _13612_ ;
wire _13613_ ;
wire _13614_ ;
wire _13615_ ;
wire _13616_ ;
wire _13617_ ;
wire _13618_ ;
wire _13619_ ;
wire _13620_ ;
wire _13621_ ;
wire _13622_ ;
wire _13623_ ;
wire _13624_ ;
wire _13625_ ;
wire _13626_ ;
wire _13627_ ;
wire _13628_ ;
wire _13629_ ;
wire _13630_ ;
wire _13631_ ;
wire _13632_ ;
wire _13633_ ;
wire _13634_ ;
wire _13635_ ;
wire _13636_ ;
wire _13637_ ;
wire _13638_ ;
wire _13639_ ;
wire _13640_ ;
wire _13641_ ;
wire _13642_ ;
wire _13643_ ;
wire _13644_ ;
wire _13645_ ;
wire _13646_ ;
wire _13647_ ;
wire _13648_ ;
wire _13649_ ;
wire _13650_ ;
wire _13651_ ;
wire _13652_ ;
wire _13653_ ;
wire _13654_ ;
wire _13655_ ;
wire _13656_ ;
wire _13657_ ;
wire _13658_ ;
wire _13659_ ;
wire _13660_ ;
wire _13661_ ;
wire _13662_ ;
wire _13663_ ;
wire _13664_ ;
wire _13665_ ;
wire _13666_ ;
wire _13667_ ;
wire _13668_ ;
wire _13669_ ;
wire _13670_ ;
wire _13671_ ;
wire _13672_ ;
wire _13673_ ;
wire _13674_ ;
wire _13675_ ;
wire _13676_ ;
wire _13677_ ;
wire _13678_ ;
wire _13679_ ;
wire _13680_ ;
wire _13681_ ;
wire _13682_ ;
wire _13683_ ;
wire _13684_ ;
wire _13685_ ;
wire _13686_ ;
wire _13687_ ;
wire _13688_ ;
wire _13689_ ;
wire _13690_ ;
wire _13691_ ;
wire _13692_ ;
wire _13693_ ;
wire _13694_ ;
wire _13695_ ;
wire _13696_ ;
wire _13697_ ;
wire _13698_ ;
wire _13699_ ;
wire _13700_ ;
wire _13701_ ;
wire _13702_ ;
wire _13703_ ;
wire _13704_ ;
wire _13705_ ;
wire _13706_ ;
wire _13707_ ;
wire _13708_ ;
wire _13709_ ;
wire _13710_ ;
wire _13711_ ;
wire _13712_ ;
wire _13713_ ;
wire _13714_ ;
wire _13715_ ;
wire _13716_ ;
wire _13717_ ;
wire _13718_ ;
wire _13719_ ;
wire _13720_ ;
wire _13721_ ;
wire _13722_ ;
wire _13723_ ;
wire _13724_ ;
wire _13725_ ;
wire _13726_ ;
wire _13727_ ;
wire _13728_ ;
wire _13729_ ;
wire _13730_ ;
wire _13731_ ;
wire _13732_ ;
wire _13733_ ;
wire _13734_ ;
wire _13735_ ;
wire _13736_ ;
wire _13737_ ;
wire _13738_ ;
wire _13739_ ;
wire _13740_ ;
wire _13741_ ;
wire _13742_ ;
wire _13743_ ;
wire _13744_ ;
wire _13745_ ;
wire _13746_ ;
wire _13747_ ;
wire _13748_ ;
wire _13749_ ;
wire _13750_ ;
wire _13751_ ;
wire _13752_ ;
wire _13753_ ;
wire _13754_ ;
wire _13755_ ;
wire _13756_ ;
wire _13757_ ;
wire _13758_ ;
wire _13759_ ;
wire _13760_ ;
wire _13761_ ;
wire _13762_ ;
wire _13763_ ;
wire _13764_ ;
wire _13765_ ;
wire _13766_ ;
wire _13767_ ;
wire _13768_ ;
wire _13769_ ;
wire _13770_ ;
wire _13771_ ;
wire _13772_ ;
wire _13773_ ;
wire _13774_ ;
wire _13775_ ;
wire _13776_ ;
wire _13777_ ;
wire _13778_ ;
wire _13779_ ;
wire _13780_ ;
wire _13781_ ;
wire _13782_ ;
wire _13783_ ;
wire _13784_ ;
wire _13785_ ;
wire _13786_ ;
wire _13787_ ;
wire _13788_ ;
wire _13789_ ;
wire _13790_ ;
wire _13791_ ;
wire _13792_ ;
wire _13793_ ;
wire _13794_ ;
wire _13795_ ;
wire _13796_ ;
wire _13797_ ;
wire _13798_ ;
wire _13799_ ;
wire _13800_ ;
wire _13801_ ;
wire _13802_ ;
wire _13803_ ;
wire _13804_ ;
wire _13805_ ;
wire _13806_ ;
wire _13807_ ;
wire _13808_ ;
wire _13809_ ;
wire _13810_ ;
wire _13811_ ;
wire _13812_ ;
wire _13813_ ;
wire _13814_ ;
wire _13815_ ;
wire _13816_ ;
wire _13817_ ;
wire _13818_ ;
wire _13819_ ;
wire _13820_ ;
wire _13821_ ;
wire _13822_ ;
wire _13823_ ;
wire _13824_ ;
wire _13825_ ;
wire _13826_ ;
wire _13827_ ;
wire _13828_ ;
wire _13829_ ;
wire _13830_ ;
wire _13831_ ;
wire _13832_ ;
wire _13833_ ;
wire _13834_ ;
wire _13835_ ;
wire _13836_ ;
wire _13837_ ;
wire _13838_ ;
wire _13839_ ;
wire _13840_ ;
wire _13841_ ;
wire _13842_ ;
wire _13843_ ;
wire _13844_ ;
wire _13845_ ;
wire _13846_ ;
wire _13847_ ;
wire _13848_ ;
wire _13849_ ;
wire _13850_ ;
wire _13851_ ;
wire _13852_ ;
wire _13853_ ;
wire _13854_ ;
wire _13855_ ;
wire _13856_ ;
wire _13857_ ;
wire _13858_ ;
wire _13859_ ;
wire _13860_ ;
wire _13861_ ;
wire _13862_ ;
wire _13863_ ;
wire _13864_ ;
wire _13865_ ;
wire _13866_ ;
wire _13867_ ;
wire _13868_ ;
wire _13869_ ;
wire _13870_ ;
wire _13871_ ;
wire _13872_ ;
wire _13873_ ;
wire _13874_ ;
wire _13875_ ;
wire _13876_ ;
wire _13877_ ;
wire _13878_ ;
wire _13879_ ;
wire _13880_ ;
wire _13881_ ;
wire _13882_ ;
wire _13883_ ;
wire _13884_ ;
wire _13885_ ;
wire _13886_ ;
wire _13887_ ;
wire _13888_ ;
wire _13889_ ;
wire _13890_ ;
wire _13891_ ;
wire _13892_ ;
wire _13893_ ;
wire _13894_ ;
wire _13895_ ;
wire _13896_ ;
wire _13897_ ;
wire _13898_ ;
wire _13899_ ;
wire _13900_ ;
wire _13901_ ;
wire _13902_ ;
wire _13903_ ;
wire _13904_ ;
wire _13905_ ;
wire _13906_ ;
wire _13907_ ;
wire _13908_ ;
wire _13909_ ;
wire _13910_ ;
wire _13911_ ;
wire _13912_ ;
wire _13913_ ;
wire _13914_ ;
wire _13915_ ;
wire _13916_ ;
wire _13917_ ;
wire _13918_ ;
wire _13919_ ;
wire _13920_ ;
wire _13921_ ;
wire _13922_ ;
wire _13923_ ;
wire _13924_ ;
wire _13925_ ;
wire _13926_ ;
wire _13927_ ;
wire _13928_ ;
wire _13929_ ;
wire _13930_ ;
wire _13931_ ;
wire _13932_ ;
wire _13933_ ;
wire _13934_ ;
wire _13935_ ;
wire _13936_ ;
wire _13937_ ;
wire _13938_ ;
wire _13939_ ;
wire _13940_ ;
wire _13941_ ;
wire _13942_ ;
wire _13943_ ;
wire _13944_ ;
wire _13945_ ;
wire _13946_ ;
wire _13947_ ;
wire _13948_ ;
wire _13949_ ;
wire _13950_ ;
wire _13951_ ;
wire _13952_ ;
wire _13953_ ;
wire _13954_ ;
wire _13955_ ;
wire _13956_ ;
wire _13957_ ;
wire _13958_ ;
wire _13959_ ;
wire _13960_ ;
wire _13961_ ;
wire _13962_ ;
wire _13963_ ;
wire _13964_ ;
wire _13965_ ;
wire _13966_ ;
wire _13967_ ;
wire _13968_ ;
wire _13969_ ;
wire _13970_ ;
wire _13971_ ;
wire _13972_ ;
wire _13973_ ;
wire _13974_ ;
wire _13975_ ;
wire _13976_ ;
wire _13977_ ;
wire _13978_ ;
wire _13979_ ;
wire _13980_ ;
wire _13981_ ;
wire _13982_ ;
wire _13983_ ;
wire _13984_ ;
wire _13985_ ;
wire _13986_ ;
wire _13987_ ;
wire _13988_ ;
wire _13989_ ;
wire _13990_ ;
wire _13991_ ;
wire _13992_ ;
wire _13993_ ;
wire _13994_ ;
wire _13995_ ;
wire _13996_ ;
wire _13997_ ;
wire _13998_ ;
wire _13999_ ;
wire _14000_ ;
wire _14001_ ;
wire _14002_ ;
wire _14003_ ;
wire _14004_ ;
wire _14005_ ;
wire _14006_ ;
wire _14007_ ;
wire _14008_ ;
wire _14009_ ;
wire _14010_ ;
wire _14011_ ;
wire _14012_ ;
wire _14013_ ;
wire _14014_ ;
wire _14015_ ;
wire _14016_ ;
wire _14017_ ;
wire _14018_ ;
wire _14019_ ;
wire _14020_ ;
wire _14021_ ;
wire _14022_ ;
wire _14023_ ;
wire _14024_ ;
wire _14025_ ;
wire _14026_ ;
wire _14027_ ;
wire _14028_ ;
wire _14029_ ;
wire _14030_ ;
wire _14031_ ;
wire _14032_ ;
wire _14033_ ;
wire _14034_ ;
wire _14035_ ;
wire _14036_ ;
wire _14037_ ;
wire _14038_ ;
wire _14039_ ;
wire _14040_ ;
wire _14041_ ;
wire _14042_ ;
wire _14043_ ;
wire _14044_ ;
wire _14045_ ;
wire _14046_ ;
wire _14047_ ;
wire _14048_ ;
wire _14049_ ;
wire _14050_ ;
wire _14051_ ;
wire _14052_ ;
wire _14053_ ;
wire _14054_ ;
wire _14055_ ;
wire _14056_ ;
wire _14057_ ;
wire _14058_ ;
wire _14059_ ;
wire _14060_ ;
wire _14061_ ;
wire _14062_ ;
wire _14063_ ;
wire _14064_ ;
wire _14065_ ;
wire _14066_ ;
wire _14067_ ;
wire _14068_ ;
wire _14069_ ;
wire _14070_ ;
wire _14071_ ;
wire _14072_ ;
wire _14073_ ;
wire _14074_ ;
wire _14075_ ;
wire _14076_ ;
wire _14077_ ;
wire _14078_ ;
wire _14079_ ;
wire _14080_ ;
wire _14081_ ;
wire _14082_ ;
wire _14083_ ;
wire _14084_ ;
wire _14085_ ;
wire _14086_ ;
wire _14087_ ;
wire _14088_ ;
wire _14089_ ;
wire _14090_ ;
wire _14091_ ;
wire _14092_ ;
wire _14093_ ;
wire _14094_ ;
wire _14095_ ;
wire _14096_ ;
wire _14097_ ;
wire _14098_ ;
wire _14099_ ;
wire _14100_ ;
wire _14101_ ;
wire _14102_ ;
wire _14103_ ;
wire _14104_ ;
wire _14105_ ;
wire _14106_ ;
wire _14107_ ;
wire _14108_ ;
wire _14109_ ;
wire _14110_ ;
wire _14111_ ;
wire _14112_ ;
wire _14113_ ;
wire _14114_ ;
wire _14115_ ;
wire _14116_ ;
wire _14117_ ;
wire _14118_ ;
wire _14119_ ;
wire _14120_ ;
wire _14121_ ;
wire _14122_ ;
wire _14123_ ;
wire _14124_ ;
wire _14125_ ;
wire _14126_ ;
wire _14127_ ;
wire _14128_ ;
wire _14129_ ;
wire _14130_ ;
wire _14131_ ;
wire _14132_ ;
wire _14133_ ;
wire _14134_ ;
wire _14135_ ;
wire _14136_ ;
wire _14137_ ;
wire _14138_ ;
wire _14139_ ;
wire _14140_ ;
wire _14141_ ;
wire _14142_ ;
wire _14143_ ;
wire _14144_ ;
wire _14145_ ;
wire _14146_ ;
wire _14147_ ;
wire _14148_ ;
wire _14149_ ;
wire _14150_ ;
wire _14151_ ;
wire _14152_ ;
wire _14153_ ;
wire _14154_ ;
wire _14155_ ;
wire _14156_ ;
wire _14157_ ;
wire _14158_ ;
wire _14159_ ;
wire _14160_ ;
wire _14161_ ;
wire _14162_ ;
wire _14163_ ;
wire _14164_ ;
wire _14165_ ;
wire _14166_ ;
wire _14167_ ;
wire _14168_ ;
wire _14169_ ;
wire _14170_ ;
wire _14171_ ;
wire _14172_ ;
wire _14173_ ;
wire _14174_ ;
wire _14175_ ;
wire _14176_ ;
wire _14177_ ;
wire _14178_ ;
wire _14179_ ;
wire _14180_ ;
wire _14181_ ;
wire _14182_ ;
wire _14183_ ;
wire _14184_ ;
wire _14185_ ;
wire _14186_ ;
wire _14187_ ;
wire _14188_ ;
wire _14189_ ;
wire _14190_ ;
wire _14191_ ;
wire _14192_ ;
wire _14193_ ;
wire _14194_ ;
wire _14195_ ;
wire _14196_ ;
wire _14197_ ;
wire _14198_ ;
wire _14199_ ;
wire _14200_ ;
wire _14201_ ;
wire _14202_ ;
wire _14203_ ;
wire _14204_ ;
wire _14205_ ;
wire _14206_ ;
wire _14207_ ;
wire _14208_ ;
wire _14209_ ;
wire _14210_ ;
wire _14211_ ;
wire _14212_ ;
wire _14213_ ;
wire _14214_ ;
wire _14215_ ;
wire _14216_ ;
wire _14217_ ;
wire _14218_ ;
wire _14219_ ;
wire _14220_ ;
wire _14221_ ;
wire _14222_ ;
wire _14223_ ;
wire _14224_ ;
wire _14225_ ;
wire _14226_ ;
wire _14227_ ;
wire _14228_ ;
wire _14229_ ;
wire _14230_ ;
wire _14231_ ;
wire _14232_ ;
wire _14233_ ;
wire _14234_ ;
wire _14235_ ;
wire _14236_ ;
wire _14237_ ;
wire _14238_ ;
wire _14239_ ;
wire _14240_ ;
wire _14241_ ;
wire _14242_ ;
wire _14243_ ;
wire _14244_ ;
wire _14245_ ;
wire _14246_ ;
wire _14247_ ;
wire _14248_ ;
wire _14249_ ;
wire _14250_ ;
wire _14251_ ;
wire _14252_ ;
wire _14253_ ;
wire _14254_ ;
wire _14255_ ;
wire _14256_ ;
wire _14257_ ;
wire _14258_ ;
wire _14259_ ;
wire _14260_ ;
wire _14261_ ;
wire _14262_ ;
wire _14263_ ;
wire _14264_ ;
wire _14265_ ;
wire _14266_ ;
wire _14267_ ;
wire _14268_ ;
wire _14269_ ;
wire _14270_ ;
wire _14271_ ;
wire _14272_ ;
wire _14273_ ;
wire _14274_ ;
wire _14275_ ;
wire _14276_ ;
wire _14277_ ;
wire _14278_ ;
wire _14279_ ;
wire _14280_ ;
wire _14281_ ;
wire _14282_ ;
wire _14283_ ;
wire _14284_ ;
wire _14285_ ;
wire _14286_ ;
wire _14287_ ;
wire _14288_ ;
wire _14289_ ;
wire _14290_ ;
wire _14291_ ;
wire _14292_ ;
wire _14293_ ;
wire _14294_ ;
wire _14295_ ;
wire _14296_ ;
wire _14297_ ;
wire _14298_ ;
wire _14299_ ;
wire _14300_ ;
wire _14301_ ;
wire _14302_ ;
wire _14303_ ;
wire _14304_ ;
wire _14305_ ;
wire _14306_ ;
wire _14307_ ;
wire _14308_ ;
wire _14309_ ;
wire _14310_ ;
wire _14311_ ;
wire _14312_ ;
wire _14313_ ;
wire _14314_ ;
wire _14315_ ;
wire _14316_ ;
wire _14317_ ;
wire _14318_ ;
wire _14319_ ;
wire _14320_ ;
wire _14321_ ;
wire _14322_ ;
wire _14323_ ;
wire _14324_ ;
wire _14325_ ;
wire _14326_ ;
wire _14327_ ;
wire _14328_ ;
wire _14329_ ;
wire _14330_ ;
wire _14331_ ;
wire _14332_ ;
wire _14333_ ;
wire _14334_ ;
wire _14335_ ;
wire _14336_ ;
wire _14337_ ;
wire _14338_ ;
wire _14339_ ;
wire _14340_ ;
wire _14341_ ;
wire _14342_ ;
wire _14343_ ;
wire _14344_ ;
wire _14345_ ;
wire _14346_ ;
wire _14347_ ;
wire _14348_ ;
wire _14349_ ;
wire _14350_ ;
wire _14351_ ;
wire _14352_ ;
wire _14353_ ;
wire _14354_ ;
wire _14355_ ;
wire _14356_ ;
wire _14357_ ;
wire _14358_ ;
wire _14359_ ;
wire _14360_ ;
wire _14361_ ;
wire _14362_ ;
wire _14363_ ;
wire _14364_ ;
wire _14365_ ;
wire _14366_ ;
wire _14367_ ;
wire _14368_ ;
wire _14369_ ;
wire _14370_ ;
wire _14371_ ;
wire _14372_ ;
wire _14373_ ;
wire _14374_ ;
wire _14375_ ;
wire _14376_ ;
wire _14377_ ;
wire _14378_ ;
wire _14379_ ;
wire _14380_ ;
wire _14381_ ;
wire _14382_ ;
wire _14383_ ;
wire _14384_ ;
wire _14385_ ;
wire _14386_ ;
wire _14387_ ;
wire _14388_ ;
wire _14389_ ;
wire _14390_ ;
wire _14391_ ;
wire _14392_ ;
wire _14393_ ;
wire _14394_ ;
wire _14395_ ;
wire _14396_ ;
wire _14397_ ;
wire _14398_ ;
wire _14399_ ;
wire _14400_ ;
wire _14401_ ;
wire _14402_ ;
wire _14403_ ;
wire _14404_ ;
wire _14405_ ;
wire _14406_ ;
wire _14407_ ;
wire _14408_ ;
wire _14409_ ;
wire _14410_ ;
wire _14411_ ;
wire _14412_ ;
wire _14413_ ;
wire _14414_ ;
wire _14415_ ;
wire _14416_ ;
wire _14417_ ;
wire _14418_ ;
wire _14419_ ;
wire _14420_ ;
wire _14421_ ;
wire _14422_ ;
wire _14423_ ;
wire _14424_ ;
wire _14425_ ;
wire _14426_ ;
wire _14427_ ;
wire _14428_ ;
wire _14429_ ;
wire _14430_ ;
wire _14431_ ;
wire _14432_ ;
wire _14433_ ;
wire _14434_ ;
wire _14435_ ;
wire _14436_ ;
wire _14437_ ;
wire _14438_ ;
wire _14439_ ;
wire _14440_ ;
wire _14441_ ;
wire _14442_ ;
wire _14443_ ;
wire _14444_ ;
wire _14445_ ;
wire _14446_ ;
wire _14447_ ;
wire _14448_ ;
wire _14449_ ;
wire _14450_ ;
wire _14451_ ;
wire _14452_ ;
wire _14453_ ;
wire _14454_ ;
wire _14455_ ;
wire _14456_ ;
wire _14457_ ;
wire _14458_ ;
wire _14459_ ;
wire _14460_ ;
wire _14461_ ;
wire _14462_ ;
wire _14463_ ;
wire _14464_ ;
wire _14465_ ;
wire _14466_ ;
wire _14467_ ;
wire _14468_ ;
wire _14469_ ;
wire _14470_ ;
wire _14471_ ;
wire _14472_ ;
wire _14473_ ;
wire _14474_ ;
wire _14475_ ;
wire _14476_ ;
wire _14477_ ;
wire _14478_ ;
wire _14479_ ;
wire _14480_ ;
wire _14481_ ;
wire _14482_ ;
wire _14483_ ;
wire _14484_ ;
wire _14485_ ;
wire _14486_ ;
wire _14487_ ;
wire _14488_ ;
wire _14489_ ;
wire _14490_ ;
wire _14491_ ;
wire _14492_ ;
wire _14493_ ;
wire _14494_ ;
wire _14495_ ;
wire _14496_ ;
wire _14497_ ;
wire _14498_ ;
wire _14499_ ;
wire _14500_ ;
wire _14501_ ;
wire _14502_ ;
wire _14503_ ;
wire _14504_ ;
wire _14505_ ;
wire _14506_ ;
wire _14507_ ;
wire _14508_ ;
wire _14509_ ;
wire _14510_ ;
wire _14511_ ;
wire _14512_ ;
wire _14513_ ;
wire _14514_ ;
wire _14515_ ;
wire _14516_ ;
wire _14517_ ;
wire _14518_ ;
wire _14519_ ;
wire _14520_ ;
wire _14521_ ;
wire _14522_ ;
wire _14523_ ;
wire _14524_ ;
wire _14525_ ;
wire _14526_ ;
wire _14527_ ;
wire _14528_ ;
wire _14529_ ;
wire _14530_ ;
wire _14531_ ;
wire _14532_ ;
wire _14533_ ;
wire _14534_ ;
wire _14535_ ;
wire _14536_ ;
wire _14537_ ;
wire _14538_ ;
wire _14539_ ;
wire _14540_ ;
wire _14541_ ;
wire _14542_ ;
wire _14543_ ;
wire _14544_ ;
wire _14545_ ;
wire _14546_ ;
wire _14547_ ;
wire _14548_ ;
wire _14549_ ;
wire _14550_ ;
wire _14551_ ;
wire _14552_ ;
wire _14553_ ;
wire _14554_ ;
wire _14555_ ;
wire _14556_ ;
wire _14557_ ;
wire _14558_ ;
wire _14559_ ;
wire _14560_ ;
wire _14561_ ;
wire _14562_ ;
wire _14563_ ;
wire _14564_ ;
wire _14565_ ;
wire _14566_ ;
wire _14567_ ;
wire _14568_ ;
wire _14569_ ;
wire _14570_ ;
wire _14571_ ;
wire _14572_ ;
wire _14573_ ;
wire _14574_ ;
wire _14575_ ;
wire _14576_ ;
wire _14577_ ;
wire _14578_ ;
wire _14579_ ;
wire _14580_ ;
wire _14581_ ;
wire _14582_ ;
wire _14583_ ;
wire _14584_ ;
wire _14585_ ;
wire _14586_ ;
wire _14587_ ;
wire _14588_ ;
wire _14589_ ;
wire _14590_ ;
wire _14591_ ;
wire _14592_ ;
wire _14593_ ;
wire _14594_ ;
wire _14595_ ;
wire _14596_ ;
wire _14597_ ;
wire _14598_ ;
wire _14599_ ;
wire _14600_ ;
wire _14601_ ;
wire _14602_ ;
wire _14603_ ;
wire _14604_ ;
wire _14605_ ;
wire _14606_ ;
wire _14607_ ;
wire _14608_ ;
wire _14609_ ;
wire _14610_ ;
wire _14611_ ;
wire _14612_ ;
wire _14613_ ;
wire _14614_ ;
wire _14615_ ;
wire _14616_ ;
wire _14617_ ;
wire _14618_ ;
wire _14619_ ;
wire _14620_ ;
wire _14621_ ;
wire _14622_ ;
wire _14623_ ;
wire _14624_ ;
wire _14625_ ;
wire _14626_ ;
wire _14627_ ;
wire _14628_ ;
wire _14629_ ;
wire _14630_ ;
wire _14631_ ;
wire _14632_ ;
wire _14633_ ;
wire _14634_ ;
wire _14635_ ;
wire _14636_ ;
wire _14637_ ;
wire _14638_ ;
wire _14639_ ;
wire _14640_ ;
wire _14641_ ;
wire _14642_ ;
wire _14643_ ;
wire _14644_ ;
wire _14645_ ;
wire _14646_ ;
wire _14647_ ;
wire _14648_ ;
wire _14649_ ;
wire _14650_ ;
wire _14651_ ;
wire _14652_ ;
wire _14653_ ;
wire _14654_ ;
wire _14655_ ;
wire _14656_ ;
wire _14657_ ;
wire _14658_ ;
wire _14659_ ;
wire _14660_ ;
wire _14661_ ;
wire _14662_ ;
wire _14663_ ;
wire _14664_ ;
wire _14665_ ;
wire _14666_ ;
wire _14667_ ;
wire _14668_ ;
wire _14669_ ;
wire _14670_ ;
wire _14671_ ;
wire _14672_ ;
wire _14673_ ;
wire _14674_ ;
wire _14675_ ;
wire _14676_ ;
wire _14677_ ;
wire _14678_ ;
wire _14679_ ;
wire _14680_ ;
wire _14681_ ;
wire _14682_ ;
wire _14683_ ;
wire _14684_ ;
wire _14685_ ;
wire _14686_ ;
wire _14687_ ;
wire _14688_ ;
wire _14689_ ;
wire _14690_ ;
wire _14691_ ;
wire _14692_ ;
wire _14693_ ;
wire _14694_ ;
wire _14695_ ;
wire _14696_ ;
wire _14697_ ;
wire _14698_ ;
wire _14699_ ;
wire _14700_ ;
wire _14701_ ;
wire _14702_ ;
wire _14703_ ;
wire _14704_ ;
wire _14705_ ;
wire _14706_ ;
wire _14707_ ;
wire _14708_ ;
wire _14709_ ;
wire _14710_ ;
wire _14711_ ;
wire _14712_ ;
wire _14713_ ;
wire _14714_ ;
wire _14715_ ;
wire _14716_ ;
wire _14717_ ;
wire _14718_ ;
wire _14719_ ;
wire _14720_ ;
wire _14721_ ;
wire _14722_ ;
wire _14723_ ;
wire _14724_ ;
wire _14725_ ;
wire _14726_ ;
wire _14727_ ;
wire _14728_ ;
wire _14729_ ;
wire _14730_ ;
wire _14731_ ;
wire _14732_ ;
wire _14733_ ;
wire _14734_ ;
wire _14735_ ;
wire _14736_ ;
wire _14737_ ;
wire _14738_ ;
wire _14739_ ;
wire _14740_ ;
wire _14741_ ;
wire _14742_ ;
wire _14743_ ;
wire _14744_ ;
wire _14745_ ;
wire _14746_ ;
wire _14747_ ;
wire _14748_ ;
wire _14749_ ;
wire _14750_ ;
wire _14751_ ;
wire _14752_ ;
wire _14753_ ;
wire _14754_ ;
wire _14755_ ;
wire _14756_ ;
wire _14757_ ;
wire _14758_ ;
wire _14759_ ;
wire _14760_ ;
wire _14761_ ;
wire _14762_ ;
wire _14763_ ;
wire _14764_ ;
wire _14765_ ;
wire _14766_ ;
wire _14767_ ;
wire _14768_ ;
wire _14769_ ;
wire _14770_ ;
wire _14771_ ;
wire _14772_ ;
wire _14773_ ;
wire _14774_ ;
wire _14775_ ;
wire _14776_ ;
wire _14777_ ;
wire _14778_ ;
wire _14779_ ;
wire _14780_ ;
wire _14781_ ;
wire _14782_ ;
wire _14783_ ;
wire _14784_ ;
wire _14785_ ;
wire _14786_ ;
wire _14787_ ;
wire _14788_ ;
wire _14789_ ;
wire _14790_ ;
wire _14791_ ;
wire _14792_ ;
wire _14793_ ;
wire _14794_ ;
wire _14795_ ;
wire _14796_ ;
wire _14797_ ;
wire _14798_ ;
wire _14799_ ;
wire _14800_ ;
wire _14801_ ;
wire _14802_ ;
wire _14803_ ;
wire _14804_ ;
wire _14805_ ;
wire _14806_ ;
wire _14807_ ;
wire _14808_ ;
wire _14809_ ;
wire _14810_ ;
wire _14811_ ;
wire _14812_ ;
wire _14813_ ;
wire _14814_ ;
wire _14815_ ;
wire _14816_ ;
wire _14817_ ;
wire _14818_ ;
wire _14819_ ;
wire _14820_ ;
wire _14821_ ;
wire _14822_ ;
wire _14823_ ;
wire _14824_ ;
wire _14825_ ;
wire _14826_ ;
wire _14827_ ;
wire _14828_ ;
wire _14829_ ;
wire _14830_ ;
wire _14831_ ;
wire _14832_ ;
wire _14833_ ;
wire _14834_ ;
wire _14835_ ;
wire _14836_ ;
wire _14837_ ;
wire _14838_ ;
wire _14839_ ;
wire _14840_ ;
wire _14841_ ;
wire _14842_ ;
wire _14843_ ;
wire _14844_ ;
wire _14845_ ;
wire _14846_ ;
wire _14847_ ;
wire _14848_ ;
wire _14849_ ;
wire _14850_ ;
wire _14851_ ;
wire _14852_ ;
wire _14853_ ;
wire _14854_ ;
wire _14855_ ;
wire _14856_ ;
wire _14857_ ;
wire _14858_ ;
wire _14859_ ;
wire _14860_ ;
wire _14861_ ;
wire _14862_ ;
wire _14863_ ;
wire _14864_ ;
wire _14865_ ;
wire _14866_ ;
wire _14867_ ;
wire _14868_ ;
wire _14869_ ;
wire _14870_ ;
wire _14871_ ;
wire _14872_ ;
wire _14873_ ;
wire _14874_ ;
wire _14875_ ;
wire _14876_ ;
wire _14877_ ;
wire _14878_ ;
wire _14879_ ;
wire _14880_ ;
wire _14881_ ;
wire _14882_ ;
wire _14883_ ;
wire _14884_ ;
wire _14885_ ;
wire _14886_ ;
wire _14887_ ;
wire _14888_ ;
wire _14889_ ;
wire _14890_ ;
wire _14891_ ;
wire _14892_ ;
wire _14893_ ;
wire _14894_ ;
wire _14895_ ;
wire _14896_ ;
wire _14897_ ;
wire _14898_ ;
wire _14899_ ;
wire _14900_ ;
wire _14901_ ;
wire _14902_ ;
wire _14903_ ;
wire _14904_ ;
wire _14905_ ;
wire _14906_ ;
wire _14907_ ;
wire _14908_ ;
wire _14909_ ;
wire _14910_ ;
wire _14911_ ;
wire _14912_ ;
wire _14913_ ;
wire _14914_ ;
wire _14915_ ;
wire _14916_ ;
wire _14917_ ;
wire _14918_ ;
wire _14919_ ;
wire _14920_ ;
wire _14921_ ;
wire _14922_ ;
wire _14923_ ;
wire _14924_ ;
wire _14925_ ;
wire _14926_ ;
wire _14927_ ;
wire _14928_ ;
wire _14929_ ;
wire _14930_ ;
wire _14931_ ;
wire _14932_ ;
wire _14933_ ;
wire _14934_ ;
wire _14935_ ;
wire _14936_ ;
wire _14937_ ;
wire _14938_ ;
wire _14939_ ;
wire _14940_ ;
wire _14941_ ;
wire _14942_ ;
wire _14943_ ;
wire _14944_ ;
wire _14945_ ;
wire _14946_ ;
wire _14947_ ;
wire _14948_ ;
wire _14949_ ;
wire _14950_ ;
wire _14951_ ;
wire _14952_ ;
wire _14953_ ;
wire _14954_ ;
wire _14955_ ;
wire _14956_ ;
wire _14957_ ;
wire _14958_ ;
wire _14959_ ;
wire _14960_ ;
wire _14961_ ;
wire _14962_ ;
wire _14963_ ;
wire _14964_ ;
wire _14965_ ;
wire _14966_ ;
wire _14967_ ;
wire _14968_ ;
wire _14969_ ;
wire _14970_ ;
wire _14971_ ;
wire _14972_ ;
wire _14973_ ;
wire _14974_ ;
wire _14975_ ;
wire _14976_ ;
wire _14977_ ;
wire _14978_ ;
wire _14979_ ;
wire _14980_ ;
wire _14981_ ;
wire _14982_ ;
wire _14983_ ;
wire _14984_ ;
wire _14985_ ;
wire _14986_ ;
wire _14987_ ;
wire _14988_ ;
wire _14989_ ;
wire _14990_ ;
wire _14991_ ;
wire _14992_ ;
wire _14993_ ;
wire _14994_ ;
wire _14995_ ;
wire _14996_ ;
wire _14997_ ;
wire _14998_ ;
wire _14999_ ;
wire _15000_ ;
wire _15001_ ;
wire _15002_ ;
wire _15003_ ;
wire _15004_ ;
wire _15005_ ;
wire _15006_ ;
wire _15007_ ;
wire _15008_ ;
wire _15009_ ;
wire _15010_ ;
wire _15011_ ;
wire _15012_ ;
wire _15013_ ;
wire _15014_ ;
wire _15015_ ;
wire _15016_ ;
wire _15017_ ;
wire _15018_ ;
wire _15019_ ;
wire _15020_ ;
wire _15021_ ;
wire _15022_ ;
wire _15023_ ;
wire _15024_ ;
wire _15025_ ;
wire _15026_ ;
wire _15027_ ;
wire _15028_ ;
wire _15029_ ;
wire _15030_ ;
wire _15031_ ;
wire _15032_ ;
wire _15033_ ;
wire _15034_ ;
wire _15035_ ;
wire _15036_ ;
wire _15037_ ;
wire _15038_ ;
wire _exu_io_in_bits_T ;
wire _idu_io_in_bits_T ;
wire _lsu_io_in_bits_T ;
wire _wbu_io_in_bits_T ;
wire \arbiter._clink_io_axi_araddr_T ;
wire \arbiter._io_axi_araddr_T ;
wire \arbiter._io_axi_araddr_T_6 ;
wire \arbiter.clink.io_axi_arvalid ;
wire \arbiter.clink.io_axi_rvalid ;
wire \arbiter.clink.io_axi_rvalid_REG_$_NOT__A_Y ;
wire \arbiter.ifu_end ;
wire \arbiter.lsu_end ;
wire \arbiter.state_$_DFF_P__Q_1_D ;
wire \arbiter.state_$_DFF_P__Q_2_D ;
wire \arbiter.state_$_DFF_P__Q_D ;
wire clock ;
wire \exu.add.io_is ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_10_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_11_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_12_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_13_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_14_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_15_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_16_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_17_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_17_A_$_MUX__A_B_$_MUX__B_1_A_$_XOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_NOR__B_Y_$_XOR__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_18_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_19_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_1_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_20_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_21_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_22_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_23_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_24_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_25_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_26_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_27_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_28_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_29_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_2_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_3_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_4_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_5_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_6_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_7_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_8_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_9_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_9_A_$_MUX__A_B_$_MUX__B_1_A_$_XOR__Y_A_$_NOR__A_Y_$_XOR__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_A_$_MUX__A_B ;
wire \exu.addi._io_rd_T_4_$_NOT__Y_A_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \exu.addi._io_rd_T_4_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_B ;
wire \exu.addi.io_is ;
wire \exu.and_.io_is ;
wire \exu.andi.io_is ;
wire \exu.auipc.io_is ;
wire \exu.beq.io_is ;
wire \exu.bge.io_is ;
wire \exu.bgeu.io_is ;
wire \exu.blt.io_is ;
wire \exu.bltu.io_is ;
wire \exu.bne.io_is ;
wire \exu.csrrs.io_is ;
wire \exu.csrrw.io_is ;
wire \exu.ecall.io_is ;
wire \exu.io_in_bits_en_dnpc ;
wire \exu.io_in_bits_fencei ;
wire \exu.io_in_bits_jal ;
wire \exu.io_in_bits_jalr ;
wire \exu.io_in_bits_lb ;
wire \exu.io_in_bits_lbu ;
wire \exu.io_in_bits_lh ;
wire \exu.io_in_bits_lhu ;
wire \exu.io_in_bits_lui ;
wire \exu.io_in_bits_lw ;
wire \exu.io_in_bits_mret ;
wire \exu.io_in_bits_or ;
wire \exu.io_in_bits_ori ;
wire \exu.io_in_bits_sb ;
wire \exu.io_in_bits_sh ;
wire \exu.io_in_bits_sll ;
wire \exu.io_in_bits_slli ;
wire \exu.io_in_bits_slt ;
wire \exu.io_in_bits_slti ;
wire \exu.io_in_bits_sltiu ;
wire \exu.io_in_bits_sltu ;
wire \exu.io_in_bits_sra ;
wire \exu.io_in_bits_srai ;
wire \exu.io_in_bits_srl ;
wire \exu.io_in_bits_srli ;
wire \exu.io_in_bits_sub ;
wire \exu.io_in_bits_sw ;
wire \exu.io_in_bits_wen_csr ;
wire \exu.io_in_bits_wen_rd ;
wire \exu.io_in_bits_xor ;
wire \exu.io_in_bits_xori ;
wire \exu.io_in_valid ;
wire \exu.io_out_bits_ren ;
wire \exu.io_out_bits_wdata_$_MUX__Y_11_B_$_ANDNOT__Y_B ;
wire \exu.io_out_bits_wdata_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__A_B ;
wire \exu.io_out_bits_wdata_$_MUX__Y_12_B_$_ANDNOT__Y_B ;
wire \exu.io_out_bits_wdata_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__A_B ;
wire \exu.io_out_bits_wdata_$_MUX__Y_13_B_$_ANDNOT__Y_B ;
wire \exu.io_out_bits_wdata_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__A_B ;
wire \exu.io_out_bits_wdata_$_MUX__Y_14_B_$_ANDNOT__Y_B ;
wire \exu.io_out_bits_wdata_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__A_B ;
wire \exu.io_out_bits_wen ;
wire \exu.state ;
wire exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ;
wire exu_io_in_bits_r_lui_$_NOT__A_Y ;
wire exu_io_in_bits_r_slti_$_NOT__A_Y ;
wire exu_io_in_valid_REG_$_NOT__A_Y ;
wire \icache._icache_reg_T ;
wire \icache._io_out_arvalid_T ;
wire \icache._io_out_arvalid_T_2 ;
wire \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_E ;
wire \icache.offset_buf_$_NAND__A_Y_$_ANDNOT__B_Y ;
wire \icache.offset_buf_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \icache.offset_buf_$_OR__A_Y_$_NOR__A_Y ;
wire \icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_ANDNOT__B_Y ;
wire \icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_NOR__A_Y ;
wire \icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_ANDNOT__B_Y ;
wire \icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_NOR__A_Y ;
wire \icache.offset_buf_$_SDFFE_PP0P__Q_E ;
wire \icache.state_$_DFF_P__Q_1_D ;
wire \icache.state_$_DFF_P__Q_2_D ;
wire \icache.state_$_DFF_P__Q_D ;
wire \icache.valid_reg_0 ;
wire \icache.valid_reg_1 ;
wire \icache.valid_reg_1_$_MUX__A_Y_$_OR__B_A_$_ANDNOT__A_1_Y ;
wire \icache.valid_reg_1_$_MUX__A_Y_$_OR__B_A_$_ANDNOT__A_Y ;
wire \idu.io_in_valid ;
wire \idu.io_out_bits_add ;
wire \idu.io_out_bits_addi ;
wire \idu.io_out_bits_and ;
wire \idu.io_out_bits_andi ;
wire \idu.io_out_bits_auipc ;
wire \idu.io_out_bits_beq ;
wire \idu.io_out_bits_bge ;
wire \idu.io_out_bits_bgeu ;
wire \idu.io_out_bits_blt ;
wire \idu.io_out_bits_bltu ;
wire \idu.io_out_bits_bne ;
wire \idu.io_out_bits_csrrs ;
wire \idu.io_out_bits_csrrw ;
wire \idu.io_out_bits_en_dnpc ;
wire \idu.io_out_bits_fencei ;
wire \idu.io_out_bits_jal ;
wire \idu.io_out_bits_jalr ;
wire \idu.io_out_bits_lb ;
wire \idu.io_out_bits_lbu ;
wire \idu.io_out_bits_lh ;
wire \idu.io_out_bits_lhu ;
wire \idu.io_out_bits_lui ;
wire \idu.io_out_bits_lw ;
wire \idu.io_out_bits_or ;
wire \idu.io_out_bits_ori ;
wire \idu.io_out_bits_sb ;
wire \idu.io_out_bits_sh ;
wire \idu.io_out_bits_sll ;
wire \idu.io_out_bits_slli ;
wire \idu.io_out_bits_slt ;
wire \idu.io_out_bits_slti ;
wire \idu.io_out_bits_sltiu ;
wire \idu.io_out_bits_sltu ;
wire \idu.io_out_bits_sra ;
wire \idu.io_out_bits_srai ;
wire \idu.io_out_bits_srl ;
wire \idu.io_out_bits_srli ;
wire \idu.io_out_bits_sub ;
wire \idu.io_out_bits_sw ;
wire \idu.io_out_bits_wen_csr ;
wire \idu.io_out_bits_wen_rd ;
wire \idu.io_out_bits_xor ;
wire \idu.io_out_bits_xori ;
wire \idu.io_out_valid_REG ;
wire \idu.io_raw ;
wire \idu.io_raw_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \idu.rs_reg ;
wire \idu.rs_reg_$_DFF_P__Q_D ;
wire \idu.state ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \ifu._start_T ;
wire \ifu.io_out_bits_pc_$_MUX__Y_13_A_$_MUX__Y_A_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ;
wire \ifu.io_out_bits_pc_$_MUX__Y_9_A_$_MUX__Y_A_$_OR__Y_B_$_ANDNOT__Y_A ;
wire \ifu.io_out_bits_pc_$_NOT__Y_10_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_11_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_11_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_12_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__A_Y ;
wire \ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_14_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_15_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_1_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_2_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_3_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_4_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_5_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_6_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_7_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_8_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_9_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_9_A_$_MUX__Y_B ;
wire \ifu.io_out_bits_pc_$_NOT__Y_A_$_MUX__Y_B ;
wire \ifu.io_valid ;
wire \ifu.pc_$_SDFFE_PP0P__Q_E ;
wire \ifu.ren_REG ;
wire \ifu.ren_REG_$_DFF_P__Q_D ;
wire \ifu.ren_REG_$_DFF_P__Q_D_$_NAND__Y_B ;
wire \ifu.state_$_DFF_P__Q_1_D ;
wire \ifu.state_$_DFF_P__Q_2_D ;
wire \ifu.state_$_DFF_P__Q_D ;
wire io_interrupt ;
wire io_master_arready ;
wire io_master_arvalid ;
wire fanout_net_16 ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_rlast ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_wlast ;
wire io_master_wready ;
wire io_master_wready_$_ANDNOT__B_Y_$_OR__A_B ;
wire io_master_wstrb_$_ANDNOT__Y_A ;
wire io_master_wvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_rlast ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_wlast ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire \lsu._io_axi_awvalid_T_1 ;
wire \lsu._io_in_ready_T ;
wire \lsu.io_in_bits_ecall ;
wire \lsu.io_in_bits_lb ;
wire \lsu.io_in_bits_lbu ;
wire \lsu.io_in_bits_lh ;
wire \lsu.io_in_bits_lhu ;
wire \lsu.io_in_bits_ren ;
wire \lsu.io_in_bits_wen ;
wire \lsu.io_in_bits_wen_csr ;
wire \lsu.io_in_bits_wen_rd ;
wire \lsu.io_in_valid ;
wire \lsu.state_$_DFF_P__Q_1_D ;
wire \lsu.state_$_DFF_P__Q_2_D ;
wire \lsu.state_$_DFF_P__Q_3_D ;
wire \lsu.state_$_DFF_P__Q_D ;
wire lsu_io_in_bits_r_sb_$_ANDNOT__B_Y_$_ANDNOT__B_A ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_10_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_10_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_11_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_11_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_12_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_12_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_13_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_13_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_14_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_14_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_15_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_15_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_16_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_17_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_18_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_19_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_1_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_20_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_21_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_22_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_23_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_2_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_3_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_4_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_5_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_6_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_7_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_8_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_8_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_9_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_9_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ;
wire lsu_io_out_bits_rd_wdata_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ;
wire reset ;
wire \wbu.csr_0_$_SDFFE_PP0P__Q_E ;
wire \wbu.io_in_bits_ecall ;
wire \wbu.io_in_bits_wen_csr ;
wire \wbu.io_in_bits_wen_rd ;
wire \wbu.rf_31_$_SDFFE_PP0P__Q_E ;
wire wbu_io_in_bits_csr_waddr_$_ANDNOT__A_Y ;
wire wbu_io_in_bits_csr_waddr_$_AND__A_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_1_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_1_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_1_Y ;
wire wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ;
wire wbu_io_in_valid_REG_$_NOT__A_Y ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire [0:0] \arbiter.clink._mtime_T_1 ;
wire [31:0] \arbiter.clink.io_axi_rdata ;
wire [63:0] \arbiter.clink.mtime ;
wire [4:0] \arbiter.io_ifu_araddr ;
wire [1:0] \arbiter.io_lsu_arsize ;
wire [31:0] \exu._GEN_0 ;
wire [4:0] \exu._io_out_bits_wdata_T_1 ;
wire [31:0] \exu._io_out_bits_wdata_T_2 ;
wire [31:0] \exu.add.io_rs1_data ;
wire [31:0] \exu.addi._io_rd_T_4 ;
wire [31:0] \exu.addi.io_imm ;
wire [31:0] \exu.auipc.io_rs1_data ;
wire [31:0] \exu.csrrs.io_csr_rdata ;
wire [1:0] \exu.io_in_bits_csr_waddr ;
wire [4:0] \exu.io_in_bits_rd ;
wire [5:0] \exu.io_in_bits_shamt ;
wire [31:0] \exu.io_out_bits_csr_wdata ;
wire [31:0] \exu.io_out_bits_rd_wdata ;
wire [31:0] \icache.icache_reg_0_0 ;
wire [31:0] \icache.icache_reg_0_1 ;
wire [31:0] \icache.icache_reg_0_2 ;
wire [31:0] \icache.icache_reg_0_3 ;
wire [31:0] \icache.icache_reg_1_0 ;
wire [31:0] \icache.icache_reg_1_1 ;
wire [31:0] \icache.icache_reg_1_2 ;
wire [31:0] \icache.icache_reg_1_3 ;
wire [1:0] \icache.offset_buf ;
wire [26:0] \icache.tag_reg_0 ;
wire [26:0] \icache.tag_reg_1 ;
wire [0:0] \idu._io_csr_raddr_T_14 ;
wire [1:0] \idu._io_csr_raddr_T_15 ;
wire [1:0] \idu._io_out_bits_csr_waddr_T_16 ;
wire [0:0] \idu.funct7 ;
wire [11:0] \idu.immB ;
wire [4:0] \idu.immI ;
wire [31:0] \idu.io_in_bits_inst ;
wire [31:0] \idu.io_in_bits_pc ;
wire [31:0] \idu.io_out_bits_imm ;
wire [31:0] \idu.io_out_bits_rs1_data ;
wire [31:0] \idu.io_out_bits_rs2_data ;
wire [1:0] \ifu._pc_T_8 ;
wire [0:0] \ifu._start_T_2 ;
wire [31:0] \ifu.inst ;
wire [31:0] \ifu.io_out_bits_inst ;
wire [31:0] \ifu.io_out_bits_pc ;
wire [31:0] \ifu.pc ;
wire [1:0] \ifu.start ;
wire [2:0] \ifu.state ;
wire [31:0] io_master_araddr ;
wire [1:0] io_master_arburst ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [31:0] io_master_awaddr ;
wire [1:0] io_master_awburst ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [3:0] io_master_bid ;
wire [1:0] io_master_bresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [31:0] io_slave_araddr ;
wire [1:0] io_slave_arburst ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [31:0] io_slave_awaddr ;
wire [1:0] io_slave_awburst ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [3:0] io_slave_bid ;
wire [1:0] io_slave_bresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [0:0] \lsu._GEN_1 ;
wire [1:0] \lsu.io_in_bits_csr_waddr ;
wire [31:0] \lsu.io_in_bits_csr_wdata ;
wire [31:0] \lsu.io_in_bits_pc ;
wire [4:0] \lsu.io_in_bits_rd ;
wire [31:0] \lsu.io_in_bits_rd_wdata ;
wire [31:0] \lsu.io_out_bits_rd_wdata ;
wire [1:0] \lsu.state ;
wire [31:0] \wbu._GEN_135 ;
wire [31:0] \wbu._GEN_71 ;
wire [0:0] \wbu.csr_0 ;
wire [31:0] \wbu.csr_2 ;
wire [31:0] \wbu.csr_3 ;
wire [1:0] \wbu.io_in_bits_csr_waddr ;
wire [31:0] \wbu.io_in_bits_csr_wdata ;
wire [31:0] \wbu.io_in_bits_pc ;
wire [4:0] \wbu.io_in_bits_rd ;
wire [31:0] \wbu.io_in_bits_rd_wdata ;
wire [31:0] \wbu.rf_10 ;
wire [31:0] \wbu.rf_11 ;
wire [31:0] \wbu.rf_12 ;
wire [31:0] \wbu.rf_13 ;
wire [31:0] \wbu.rf_14 ;
wire [31:0] \wbu.rf_15 ;
wire [31:0] \wbu.rf_16 ;
wire [31:0] \wbu.rf_17 ;
wire [31:0] \wbu.rf_18 ;
wire [31:0] \wbu.rf_19 ;
wire [31:0] \wbu.rf_20 ;
wire [31:0] \wbu.rf_21 ;
wire [31:0] \wbu.rf_22 ;
wire [31:0] \wbu.rf_23 ;
wire [31:0] \wbu.rf_24 ;
wire [31:0] \wbu.rf_25 ;
wire [31:0] \wbu.rf_26 ;
wire [31:0] \wbu.rf_27 ;
wire [31:0] \wbu.rf_28 ;
wire [31:0] \wbu.rf_29 ;
wire [31:0] \wbu.rf_2 ;
wire [31:0] \wbu.rf_30 ;
wire [31:0] \wbu.rf_31 ;
wire [31:0] \wbu.rf_3 ;
wire [31:0] \wbu.rf_4 ;
wire [31:0] \wbu.rf_5 ;
wire [31:0] \wbu.rf_6 ;
wire [31:0] \wbu.rf_7 ;
wire [31:0] \wbu.rf_8 ;
wire [31:0] \wbu.rf_9 ;

assign \io_master_arid [0] = \io_master_arburst [1] ;
assign \io_master_arid [1] = \io_master_arburst [1] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [1] = \io_master_arlen [0] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign \io_master_arsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign \io_master_awid [0] = \io_master_arburst [1] ;
assign \io_master_awid [1] = \io_master_arburst [1] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awburst [0] ;
assign io_master_wvalid = io_master_awvalid ;
assign io_slave_arready = \io_master_awburst [0] ;
assign io_slave_awready = \io_master_awburst [0] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_awburst [0] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_awburst [0] ;

NOR2_X1 _15039_ ( .A1(\io_master_awaddr [28] ), .A2(\io_master_awaddr [27] ), .ZN(_08532_ ) );
INV_X1 _15040_ ( .A(\io_master_awaddr [26] ), .ZN(_08533_ ) );
INV_X1 _15041_ ( .A(\io_master_awaddr [24] ), .ZN(_08534_ ) );
AND3_X1 _15042_ ( .A1(_08532_ ), .A2(_08533_ ), .A3(_08534_ ), .ZN(_08535_ ) );
INV_X1 _15043_ ( .A(\io_master_awaddr [5] ), .ZN(_08536_ ) );
INV_X1 _15044_ ( .A(\io_master_awaddr [4] ), .ZN(_08537_ ) );
INV_X1 _15045_ ( .A(\io_master_awaddr [3] ), .ZN(_08538_ ) );
AND4_X1 _15046_ ( .A1(_08536_ ), .A2(_08537_ ), .A3(_08538_ ), .A4(\io_master_awaddr [25] ), .ZN(_08539_ ) );
AND2_X1 _15047_ ( .A1(_08535_ ), .A2(_08539_ ), .ZN(_08540_ ) );
INV_X1 _15048_ ( .A(\io_master_awaddr [29] ), .ZN(_08541_ ) );
NOR2_X1 _15049_ ( .A1(\io_master_awaddr [31] ), .A2(\io_master_awaddr [30] ), .ZN(_08542_ ) );
NOR2_X1 _15050_ ( .A1(\io_master_awaddr [14] ), .A2(\io_master_awaddr [13] ), .ZN(_08543_ ) );
NOR2_X1 _15051_ ( .A1(\io_master_awaddr [15] ), .A2(\io_master_awaddr [12] ), .ZN(_08544_ ) );
AND2_X1 _15052_ ( .A1(_08543_ ), .A2(_08544_ ), .ZN(_08545_ ) );
NAND4_X1 _15053_ ( .A1(_08540_ ), .A2(_08541_ ), .A3(_08542_ ), .A4(_08545_ ), .ZN(_08546_ ) );
BUF_X2 _15054_ ( .A(_08546_ ), .Z(_08547_ ) );
NOR2_X1 _15055_ ( .A1(\io_master_awaddr [23] ), .A2(\io_master_awaddr [22] ), .ZN(_08548_ ) );
INV_X1 _15056_ ( .A(\io_master_awaddr [21] ), .ZN(_08549_ ) );
INV_X1 _15057_ ( .A(\io_master_awaddr [20] ), .ZN(_08550_ ) );
NAND3_X1 _15058_ ( .A1(_08548_ ), .A2(_08549_ ), .A3(_08550_ ), .ZN(_08551_ ) );
NOR2_X1 _15059_ ( .A1(\io_master_awaddr [17] ), .A2(\io_master_awaddr [16] ), .ZN(_08552_ ) );
INV_X1 _15060_ ( .A(\io_master_awaddr [19] ), .ZN(_08553_ ) );
INV_X1 _15061_ ( .A(\io_master_awaddr [18] ), .ZN(_08554_ ) );
NAND3_X1 _15062_ ( .A1(_08552_ ), .A2(_08553_ ), .A3(_08554_ ), .ZN(_08555_ ) );
NOR2_X1 _15063_ ( .A1(_08551_ ), .A2(_08555_ ), .ZN(_08556_ ) );
NOR4_X1 _15064_ ( .A1(\io_master_awaddr [9] ), .A2(\io_master_awaddr [8] ), .A3(\io_master_awaddr [7] ), .A4(\io_master_awaddr [6] ), .ZN(_08557_ ) );
NOR4_X1 _15065_ ( .A1(\io_master_awaddr [11] ), .A2(\io_master_awaddr [10] ), .A3(\io_master_awaddr [1] ), .A4(\io_master_awaddr [0] ), .ZN(_08558_ ) );
NAND3_X1 _15066_ ( .A1(_08556_ ), .A2(_08557_ ), .A3(_08558_ ), .ZN(_08559_ ) );
BUF_X2 _15067_ ( .A(_08559_ ), .Z(_08560_ ) );
NOR3_X1 _15068_ ( .A1(_08547_ ), .A2(\arbiter.clink.io_axi_rvalid_REG_$_NOT__A_Y ), .A3(_08560_ ), .ZN(_08561_ ) );
NOR2_X2 _15069_ ( .A1(_08546_ ), .A2(_08559_ ), .ZN(_08562_ ) );
INV_X1 _15070_ ( .A(_08562_ ), .ZN(_08563_ ) );
AOI21_X1 _15071_ ( .A(_08561_ ), .B1(_08563_ ), .B2(io_master_rvalid ), .ZN(_08564_ ) );
INV_X1 _15072_ ( .A(io_master_bvalid ), .ZN(_08565_ ) );
NAND2_X1 _15073_ ( .A1(_08564_ ), .A2(_08565_ ), .ZN(_08566_ ) );
NAND3_X1 _15074_ ( .A1(_08566_ ), .A2(io_master_bready ), .A3(fanout_net_1 ), .ZN(_08567_ ) );
NOR2_X1 _15075_ ( .A1(\lsu.io_in_bits_ren ), .A2(\lsu.io_in_bits_wen ), .ZN(_08568_ ) );
NAND3_X1 _15076_ ( .A1(_08568_ ), .A2(\lsu.io_in_valid ), .A3(\lsu._io_in_ready_T ), .ZN(_08569_ ) );
AND2_X2 _15077_ ( .A1(_08567_ ), .A2(_08569_ ), .ZN(_08570_ ) );
INV_X1 _15078_ ( .A(_08570_ ), .ZN(_wbu_io_in_bits_T ) );
INV_X1 _15079_ ( .A(fanout_net_29 ), .ZN(_08571_ ) );
NOR2_X1 _15080_ ( .A1(\wbu.io_in_bits_rd [3] ), .A2(\wbu.io_in_bits_rd [2] ), .ZN(_08572_ ) );
BUF_X2 _15081_ ( .A(_08572_ ), .Z(_08573_ ) );
BUF_X2 _15082_ ( .A(_08573_ ), .Z(_08574_ ) );
BUF_X2 _15083_ ( .A(_08574_ ), .Z(_08575_ ) );
INV_X1 _15084_ ( .A(\wbu.io_in_bits_rd [1] ), .ZN(_08576_ ) );
AND4_X1 _15085_ ( .A1(_08571_ ), .A2(_08575_ ), .A3(\wbu.io_in_bits_rd [0] ), .A4(_08576_ ), .ZN(_00000_ ) );
INV_X1 _15086_ ( .A(\wbu.io_in_bits_csr_waddr [0] ), .ZN(_08577_ ) );
BUF_X4 _15087_ ( .A(_08577_ ), .Z(_08578_ ) );
NOR2_X1 _15088_ ( .A1(_08578_ ), .A2(fanout_net_28 ), .ZN(_00001_ ) );
XOR2_X1 _15089_ ( .A(\exu.addi.io_imm [16] ), .B(\exu.auipc.io_rs1_data [16] ), .Z(_08579_ ) );
XOR2_X1 _15090_ ( .A(\exu.addi.io_imm [17] ), .B(\exu.auipc.io_rs1_data [17] ), .Z(_08580_ ) );
AND2_X1 _15091_ ( .A1(_08579_ ), .A2(_08580_ ), .ZN(_08581_ ) );
XOR2_X1 _15092_ ( .A(\exu.auipc.io_rs1_data [19] ), .B(\exu.addi.io_imm [19] ), .Z(_08582_ ) );
XOR2_X1 _15093_ ( .A(\exu.auipc.io_rs1_data [18] ), .B(\exu.addi.io_imm [18] ), .Z(_08583_ ) );
AND3_X1 _15094_ ( .A1(_08581_ ), .A2(_08582_ ), .A3(_08583_ ), .ZN(_08584_ ) );
XOR2_X1 _15095_ ( .A(\exu.addi.io_imm [4] ), .B(\exu.auipc.io_rs1_data [4] ), .Z(_08585_ ) );
NOR2_X1 _15096_ ( .A1(\exu.auipc.io_rs1_data [3] ), .A2(\exu.addi.io_imm [3] ), .ZN(_08586_ ) );
XOR2_X1 _15097_ ( .A(\exu.addi.io_imm [1] ), .B(\exu.auipc.io_rs1_data [1] ), .Z(_08587_ ) );
AND2_X1 _15098_ ( .A1(\exu.addi.io_imm [0] ), .A2(\exu.auipc.io_rs1_data [0] ), .ZN(_08588_ ) );
NAND2_X1 _15099_ ( .A1(_08587_ ), .A2(_08588_ ), .ZN(_08589_ ) );
INV_X1 _15100_ ( .A(\exu.addi.io_imm [1] ), .ZN(_08590_ ) );
INV_X1 _15101_ ( .A(\exu.auipc.io_rs1_data [1] ), .ZN(_08591_ ) );
OAI21_X1 _15102_ ( .A(_08589_ ), .B1(_08590_ ), .B2(_08591_ ), .ZN(_08592_ ) );
XOR2_X1 _15103_ ( .A(\exu.auipc.io_rs1_data [2] ), .B(\exu.addi.io_imm [2] ), .Z(_08593_ ) );
NAND2_X1 _15104_ ( .A1(_08592_ ), .A2(_08593_ ), .ZN(_08594_ ) );
NAND2_X1 _15105_ ( .A1(\exu.auipc.io_rs1_data [2] ), .A2(\exu.addi.io_imm [2] ), .ZN(_08595_ ) );
AOI21_X1 _15106_ ( .A(_08586_ ), .B1(_08594_ ), .B2(_08595_ ), .ZN(_08596_ ) );
AND2_X1 _15107_ ( .A1(\exu.auipc.io_rs1_data [3] ), .A2(\exu.addi.io_imm [3] ), .ZN(_08597_ ) );
OR2_X1 _15108_ ( .A1(_08596_ ), .A2(_08597_ ), .ZN(_08598_ ) );
XOR2_X1 _15109_ ( .A(\exu.auipc.io_rs1_data [7] ), .B(\exu.addi.io_imm [7] ), .Z(_08599_ ) );
XOR2_X1 _15110_ ( .A(\exu.auipc.io_rs1_data [6] ), .B(\exu.addi.io_imm [6] ), .Z(_08600_ ) );
AND2_X1 _15111_ ( .A1(_08599_ ), .A2(_08600_ ), .ZN(_08601_ ) );
XOR2_X1 _15112_ ( .A(\exu.addi.io_imm [5] ), .B(\exu.auipc.io_rs1_data [5] ), .Z(_08602_ ) );
AND4_X1 _15113_ ( .A1(_08585_ ), .A2(_08598_ ), .A3(_08601_ ), .A4(_08602_ ), .ZN(_08603_ ) );
AND2_X1 _15114_ ( .A1(\exu.auipc.io_rs1_data [6] ), .A2(\exu.addi.io_imm [6] ), .ZN(_08604_ ) );
AND2_X1 _15115_ ( .A1(_08599_ ), .A2(_08604_ ), .ZN(_08605_ ) );
NAND2_X1 _15116_ ( .A1(\exu.addi.io_imm [4] ), .A2(\exu.auipc.io_rs1_data [4] ), .ZN(_08606_ ) );
INV_X1 _15117_ ( .A(\exu.addi.io_imm [5] ), .ZN(_08607_ ) );
INV_X1 _15118_ ( .A(\exu.auipc.io_rs1_data [5] ), .ZN(_08608_ ) );
OAI21_X1 _15119_ ( .A(_08606_ ), .B1(_08607_ ), .B2(_08608_ ), .ZN(_08609_ ) );
NOR2_X1 _15120_ ( .A1(\exu.addi.io_imm [5] ), .A2(\exu.auipc.io_rs1_data [5] ), .ZN(_08610_ ) );
INV_X1 _15121_ ( .A(_08610_ ), .ZN(_08611_ ) );
AND2_X1 _15122_ ( .A1(_08609_ ), .A2(_08611_ ), .ZN(_08612_ ) );
AOI221_X4 _15123_ ( .A(_08605_ ), .B1(\exu.auipc.io_rs1_data [7] ), .B2(\exu.addi.io_imm [7] ), .C1(_08601_ ), .C2(_08612_ ), .ZN(_08613_ ) );
INV_X1 _15124_ ( .A(_08613_ ), .ZN(_08614_ ) );
NOR2_X1 _15125_ ( .A1(_08603_ ), .A2(_08614_ ), .ZN(_08615_ ) );
INV_X1 _15126_ ( .A(_08615_ ), .ZN(_08616_ ) );
XOR2_X1 _15127_ ( .A(\exu.auipc.io_rs1_data [8] ), .B(\exu.addi.io_imm [8] ), .Z(_08617_ ) );
AND2_X1 _15128_ ( .A1(\exu.auipc.io_rs1_data [9] ), .A2(\exu.addi.io_imm [9] ), .ZN(_08618_ ) );
NOR2_X1 _15129_ ( .A1(\exu.auipc.io_rs1_data [9] ), .A2(\exu.addi.io_imm [9] ), .ZN(_08619_ ) );
NOR2_X1 _15130_ ( .A1(_08618_ ), .A2(_08619_ ), .ZN(_08620_ ) );
AND2_X1 _15131_ ( .A1(_08617_ ), .A2(_08620_ ), .ZN(_08621_ ) );
AND2_X1 _15132_ ( .A1(_08616_ ), .A2(_08621_ ), .ZN(_08622_ ) );
XOR2_X1 _15133_ ( .A(\exu.auipc.io_rs1_data [11] ), .B(\exu.addi.io_imm [11] ), .Z(_08623_ ) );
XOR2_X1 _15134_ ( .A(\exu.auipc.io_rs1_data [10] ), .B(\exu.addi.io_imm [10] ), .Z(_08624_ ) );
AND3_X1 _15135_ ( .A1(_08622_ ), .A2(_08623_ ), .A3(_08624_ ), .ZN(_08625_ ) );
XOR2_X1 _15136_ ( .A(\exu.auipc.io_rs1_data [15] ), .B(\exu.addi.io_imm [15] ), .Z(_08626_ ) );
XOR2_X1 _15137_ ( .A(\exu.auipc.io_rs1_data [14] ), .B(\exu.addi.io_imm [14] ), .Z(_08627_ ) );
AND2_X1 _15138_ ( .A1(_08626_ ), .A2(_08627_ ), .ZN(_08628_ ) );
AND2_X1 _15139_ ( .A1(\exu.auipc.io_rs1_data [13] ), .A2(\exu.addi.io_imm [13] ), .ZN(_08629_ ) );
NOR2_X1 _15140_ ( .A1(\exu.auipc.io_rs1_data [13] ), .A2(\exu.addi.io_imm [13] ), .ZN(_08630_ ) );
NOR2_X1 _15141_ ( .A1(_08629_ ), .A2(_08630_ ), .ZN(_08631_ ) );
XOR2_X1 _15142_ ( .A(\exu.auipc.io_rs1_data [12] ), .B(\exu.addi.io_imm [12] ), .Z(_08632_ ) );
AND3_X1 _15143_ ( .A1(_08628_ ), .A2(_08631_ ), .A3(_08632_ ), .ZN(_08633_ ) );
AND2_X1 _15144_ ( .A1(_08625_ ), .A2(_08633_ ), .ZN(_08634_ ) );
AND2_X1 _15145_ ( .A1(\exu.auipc.io_rs1_data [11] ), .A2(\exu.addi.io_imm [11] ), .ZN(_08635_ ) );
AND2_X1 _15146_ ( .A1(\exu.auipc.io_rs1_data [10] ), .A2(\exu.addi.io_imm [10] ), .ZN(_08636_ ) );
AOI21_X1 _15147_ ( .A(_08635_ ), .B1(_08623_ ), .B2(_08636_ ), .ZN(_08637_ ) );
AND2_X1 _15148_ ( .A1(\exu.auipc.io_rs1_data [8] ), .A2(\exu.addi.io_imm [8] ), .ZN(_08638_ ) );
INV_X1 _15149_ ( .A(_08638_ ), .ZN(_08639_ ) );
NOR3_X1 _15150_ ( .A1(_08639_ ), .A2(_08618_ ), .A3(_08619_ ), .ZN(_08640_ ) );
OAI211_X1 _15151_ ( .A(_08623_ ), .B(_08624_ ), .C1(_08640_ ), .C2(_08618_ ), .ZN(_08641_ ) );
NAND2_X1 _15152_ ( .A1(_08637_ ), .A2(_08641_ ), .ZN(_08642_ ) );
NAND2_X1 _15153_ ( .A1(_08642_ ), .A2(_08633_ ), .ZN(_08643_ ) );
AND2_X1 _15154_ ( .A1(\exu.auipc.io_rs1_data [14] ), .A2(\exu.addi.io_imm [14] ), .ZN(_08644_ ) );
AND2_X1 _15155_ ( .A1(_08626_ ), .A2(_08644_ ), .ZN(_08645_ ) );
AND2_X1 _15156_ ( .A1(\exu.auipc.io_rs1_data [12] ), .A2(\exu.addi.io_imm [12] ), .ZN(_08646_ ) );
NAND2_X1 _15157_ ( .A1(_08631_ ), .A2(_08646_ ), .ZN(_08647_ ) );
INV_X1 _15158_ ( .A(\exu.auipc.io_rs1_data [13] ), .ZN(_08648_ ) );
INV_X1 _15159_ ( .A(\exu.addi.io_imm [13] ), .ZN(_08649_ ) );
OAI21_X1 _15160_ ( .A(_08647_ ), .B1(_08648_ ), .B2(_08649_ ), .ZN(_08650_ ) );
AOI221_X4 _15161_ ( .A(_08645_ ), .B1(\exu.auipc.io_rs1_data [15] ), .B2(\exu.addi.io_imm [15] ), .C1(_08628_ ), .C2(_08650_ ), .ZN(_08651_ ) );
AND2_X1 _15162_ ( .A1(_08643_ ), .A2(_08651_ ), .ZN(_08652_ ) );
INV_X1 _15163_ ( .A(_08652_ ), .ZN(_08653_ ) );
OAI21_X1 _15164_ ( .A(_08584_ ), .B1(_08634_ ), .B2(_08653_ ), .ZN(_08654_ ) );
XOR2_X1 _15165_ ( .A(\exu.addi.io_imm [23] ), .B(\exu.auipc.io_rs1_data [23] ), .Z(_08655_ ) );
XOR2_X1 _15166_ ( .A(\exu.addi.io_imm [22] ), .B(\exu.auipc.io_rs1_data [22] ), .Z(_08656_ ) );
AND2_X1 _15167_ ( .A1(_08655_ ), .A2(_08656_ ), .ZN(_08657_ ) );
XOR2_X1 _15168_ ( .A(\exu.addi.io_imm [20] ), .B(\exu.auipc.io_rs1_data [20] ), .Z(_08658_ ) );
AND2_X1 _15169_ ( .A1(\exu.addi.io_imm [21] ), .A2(\exu.auipc.io_rs1_data [21] ), .ZN(_08659_ ) );
NOR2_X1 _15170_ ( .A1(\exu.addi.io_imm [21] ), .A2(\exu.auipc.io_rs1_data [21] ), .ZN(_08660_ ) );
NOR2_X1 _15171_ ( .A1(_08659_ ), .A2(_08660_ ), .ZN(_08661_ ) );
AND2_X1 _15172_ ( .A1(_08658_ ), .A2(_08661_ ), .ZN(_08662_ ) );
NAND2_X1 _15173_ ( .A1(_08657_ ), .A2(_08662_ ), .ZN(_08663_ ) );
OR2_X1 _15174_ ( .A1(_08654_ ), .A2(_08663_ ), .ZN(_08664_ ) );
AND2_X1 _15175_ ( .A1(\exu.addi.io_imm [22] ), .A2(\exu.auipc.io_rs1_data [22] ), .ZN(_08665_ ) );
NAND2_X1 _15176_ ( .A1(_08655_ ), .A2(_08665_ ), .ZN(_08666_ ) );
INV_X1 _15177_ ( .A(\exu.addi.io_imm [23] ), .ZN(_08667_ ) );
INV_X1 _15178_ ( .A(\exu.auipc.io_rs1_data [23] ), .ZN(_08668_ ) );
AND2_X1 _15179_ ( .A1(\exu.addi.io_imm [16] ), .A2(\exu.auipc.io_rs1_data [16] ), .ZN(_08669_ ) );
AND2_X1 _15180_ ( .A1(_08580_ ), .A2(_08669_ ), .ZN(_08670_ ) );
AOI21_X1 _15181_ ( .A(_08670_ ), .B1(\exu.addi.io_imm [17] ), .B2(\exu.auipc.io_rs1_data [17] ), .ZN(_08671_ ) );
INV_X1 _15182_ ( .A(_08583_ ), .ZN(_08672_ ) );
AND2_X1 _15183_ ( .A1(\exu.auipc.io_rs1_data [19] ), .A2(\exu.addi.io_imm [19] ), .ZN(_08673_ ) );
NOR2_X1 _15184_ ( .A1(\exu.auipc.io_rs1_data [19] ), .A2(\exu.addi.io_imm [19] ), .ZN(_08674_ ) );
NOR4_X1 _15185_ ( .A1(_08671_ ), .A2(_08672_ ), .A3(_08673_ ), .A4(_08674_ ), .ZN(_08675_ ) );
NAND2_X1 _15186_ ( .A1(\exu.auipc.io_rs1_data [18] ), .A2(\exu.addi.io_imm [18] ), .ZN(_08676_ ) );
NOR3_X1 _15187_ ( .A1(_08673_ ), .A2(_08674_ ), .A3(_08676_ ), .ZN(_08677_ ) );
NOR3_X1 _15188_ ( .A1(_08675_ ), .A2(_08673_ ), .A3(_08677_ ), .ZN(_08678_ ) );
OAI221_X1 _15189_ ( .A(_08666_ ), .B1(_08667_ ), .B2(_08668_ ), .C1(_08678_ ), .C2(_08663_ ), .ZN(_08679_ ) );
AND2_X1 _15190_ ( .A1(\exu.addi.io_imm [20] ), .A2(\exu.auipc.io_rs1_data [20] ), .ZN(_08680_ ) );
INV_X1 _15191_ ( .A(_08680_ ), .ZN(_08681_ ) );
NOR3_X1 _15192_ ( .A1(_08681_ ), .A2(_08659_ ), .A3(_08660_ ), .ZN(_08682_ ) );
OR2_X1 _15193_ ( .A1(_08682_ ), .A2(_08659_ ), .ZN(_08683_ ) );
AOI21_X1 _15194_ ( .A(_08679_ ), .B1(_08657_ ), .B2(_08683_ ), .ZN(_08684_ ) );
NAND2_X1 _15195_ ( .A1(_08664_ ), .A2(_08684_ ), .ZN(_08685_ ) );
XOR2_X1 _15196_ ( .A(\exu.addi.io_imm [24] ), .B(\exu.auipc.io_rs1_data [24] ), .Z(_08686_ ) );
AND2_X1 _15197_ ( .A1(\exu.addi.io_imm [25] ), .A2(\exu.auipc.io_rs1_data [25] ), .ZN(_08687_ ) );
NOR2_X1 _15198_ ( .A1(\exu.addi.io_imm [25] ), .A2(\exu.auipc.io_rs1_data [25] ), .ZN(_08688_ ) );
NOR2_X1 _15199_ ( .A1(_08687_ ), .A2(_08688_ ), .ZN(_08689_ ) );
AND3_X1 _15200_ ( .A1(_08685_ ), .A2(_08686_ ), .A3(_08689_ ), .ZN(_08690_ ) );
AND2_X1 _15201_ ( .A1(\exu.addi.io_imm [24] ), .A2(\exu.auipc.io_rs1_data [24] ), .ZN(_08691_ ) );
INV_X1 _15202_ ( .A(_08691_ ), .ZN(_08692_ ) );
INV_X1 _15203_ ( .A(_08687_ ), .ZN(_08693_ ) );
AOI21_X1 _15204_ ( .A(_08688_ ), .B1(_08692_ ), .B2(_08693_ ), .ZN(_08694_ ) );
NOR2_X1 _15205_ ( .A1(_08690_ ), .A2(_08694_ ), .ZN(_08695_ ) );
XNOR2_X1 _15206_ ( .A(\exu.addi.io_imm [26] ), .B(\exu.auipc.io_rs1_data [26] ), .ZN(_08696_ ) );
XOR2_X1 _15207_ ( .A(_08695_ ), .B(_08696_ ), .Z(_08697_ ) );
INV_X1 _15208_ ( .A(fanout_net_9 ), .ZN(_08698_ ) );
NOR2_X1 _15209_ ( .A1(_08698_ ), .A2(fanout_net_17 ), .ZN(_08699_ ) );
BUF_X4 _15210_ ( .A(_08699_ ), .Z(_08700_ ) );
NAND2_X1 _15211_ ( .A1(_08697_ ), .A2(_08700_ ), .ZN(_08701_ ) );
BUF_X4 _15212_ ( .A(_08698_ ), .Z(_08702_ ) );
INV_X1 _15213_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_5_A_$_MUX__A_B ), .ZN(_08703_ ) );
AOI21_X1 _15214_ ( .A(_08702_ ), .B1(fanout_net_17 ), .B2(_08703_ ), .ZN(_08704_ ) );
XOR2_X1 _15215_ ( .A(\exu.add.io_rs1_data [10] ), .B(\exu._GEN_0 [10] ), .Z(_08705_ ) );
AND2_X1 _15216_ ( .A1(\exu.add.io_rs1_data [11] ), .A2(\exu._GEN_0 [11] ), .ZN(_08706_ ) );
NOR2_X1 _15217_ ( .A1(\exu.add.io_rs1_data [11] ), .A2(\exu._GEN_0 [11] ), .ZN(_08707_ ) );
NOR2_X1 _15218_ ( .A1(_08706_ ), .A2(_08707_ ), .ZN(_08708_ ) );
NOR2_X1 _15219_ ( .A1(_08705_ ), .A2(_08708_ ), .ZN(_08709_ ) );
AND2_X1 _15220_ ( .A1(\exu.add.io_rs1_data [9] ), .A2(\exu._GEN_0 [9] ), .ZN(_08710_ ) );
NOR2_X1 _15221_ ( .A1(\exu.add.io_rs1_data [9] ), .A2(\exu._GEN_0 [9] ), .ZN(_08711_ ) );
NOR2_X1 _15222_ ( .A1(_08710_ ), .A2(_08711_ ), .ZN(_08712_ ) );
INV_X1 _15223_ ( .A(_08712_ ), .ZN(_08713_ ) );
XOR2_X1 _15224_ ( .A(\exu.add.io_rs1_data [8] ), .B(\exu._GEN_0 [8] ), .Z(_08714_ ) );
INV_X1 _15225_ ( .A(_08714_ ), .ZN(_08715_ ) );
AND3_X1 _15226_ ( .A1(_08709_ ), .A2(_08713_ ), .A3(_08715_ ), .ZN(_08716_ ) );
XOR2_X1 _15227_ ( .A(\exu.add.io_rs1_data [15] ), .B(\exu._GEN_0 [15] ), .Z(_08717_ ) );
XOR2_X1 _15228_ ( .A(\exu.add.io_rs1_data [14] ), .B(\exu._GEN_0 [14] ), .Z(_08718_ ) );
NOR2_X1 _15229_ ( .A1(_08717_ ), .A2(_08718_ ), .ZN(_08719_ ) );
XOR2_X1 _15230_ ( .A(\exu.add.io_rs1_data [12] ), .B(\exu._GEN_0 [12] ), .Z(_08720_ ) );
AND2_X1 _15231_ ( .A1(\exu.add.io_rs1_data [13] ), .A2(\exu._GEN_0 [13] ), .ZN(_08721_ ) );
NOR2_X1 _15232_ ( .A1(\exu.add.io_rs1_data [13] ), .A2(\exu._GEN_0 [13] ), .ZN(_08722_ ) );
NOR2_X1 _15233_ ( .A1(_08721_ ), .A2(_08722_ ), .ZN(_08723_ ) );
NOR2_X1 _15234_ ( .A1(_08720_ ), .A2(_08723_ ), .ZN(_08724_ ) );
AND2_X1 _15235_ ( .A1(_08719_ ), .A2(_08724_ ), .ZN(_08725_ ) );
AND2_X1 _15236_ ( .A1(_08716_ ), .A2(_08725_ ), .ZN(_08726_ ) );
XOR2_X1 _15237_ ( .A(\exu.add.io_rs1_data [6] ), .B(\exu._GEN_0 [6] ), .Z(_08727_ ) );
AND2_X2 _15238_ ( .A1(\exu.add.io_rs1_data [7] ), .A2(\exu._GEN_0 [7] ), .ZN(_08728_ ) );
NOR2_X1 _15239_ ( .A1(\exu.add.io_rs1_data [7] ), .A2(\exu._GEN_0 [7] ), .ZN(_08729_ ) );
NOR2_X1 _15240_ ( .A1(_08728_ ), .A2(_08729_ ), .ZN(_08730_ ) );
NOR2_X1 _15241_ ( .A1(_08727_ ), .A2(_08730_ ), .ZN(_08731_ ) );
XOR2_X1 _15242_ ( .A(\exu.add.io_rs1_data [4] ), .B(\exu._GEN_0 [4] ), .Z(_08732_ ) );
AND2_X1 _15243_ ( .A1(\exu.add.io_rs1_data [5] ), .A2(\exu._GEN_0 [5] ), .ZN(_08733_ ) );
NOR2_X1 _15244_ ( .A1(\exu.add.io_rs1_data [5] ), .A2(\exu._GEN_0 [5] ), .ZN(_08734_ ) );
NOR2_X1 _15245_ ( .A1(_08733_ ), .A2(_08734_ ), .ZN(_08735_ ) );
NOR2_X1 _15246_ ( .A1(_08732_ ), .A2(_08735_ ), .ZN(_08736_ ) );
AND2_X1 _15247_ ( .A1(_08731_ ), .A2(_08736_ ), .ZN(_08737_ ) );
XOR2_X1 _15248_ ( .A(\exu.add.io_rs1_data [3] ), .B(\exu._GEN_0 [3] ), .Z(_08738_ ) );
INV_X1 _15249_ ( .A(_08738_ ), .ZN(_08739_ ) );
XOR2_X1 _15250_ ( .A(\exu.add.io_rs1_data [0] ), .B(\exu._GEN_0 [0] ), .Z(_08740_ ) );
INV_X1 _15251_ ( .A(_08740_ ), .ZN(_08741_ ) );
AND4_X1 _15252_ ( .A1(_08726_ ), .A2(_08737_ ), .A3(_08739_ ), .A4(_08741_ ), .ZN(_08742_ ) );
XOR2_X1 _15253_ ( .A(\exu.add.io_rs1_data [19] ), .B(\exu._GEN_0 [19] ), .Z(_08743_ ) );
XOR2_X1 _15254_ ( .A(\exu.add.io_rs1_data [18] ), .B(\exu._GEN_0 [18] ), .Z(_08744_ ) );
NOR2_X1 _15255_ ( .A1(_08743_ ), .A2(_08744_ ), .ZN(_08745_ ) );
XOR2_X1 _15256_ ( .A(\exu.add.io_rs1_data [17] ), .B(\exu._GEN_0 [17] ), .Z(_08746_ ) );
INV_X1 _15257_ ( .A(_08746_ ), .ZN(_08747_ ) );
XOR2_X1 _15258_ ( .A(\exu.add.io_rs1_data [16] ), .B(\exu._GEN_0 [16] ), .Z(_08748_ ) );
INV_X1 _15259_ ( .A(_08748_ ), .ZN(_08749_ ) );
AND3_X1 _15260_ ( .A1(_08745_ ), .A2(_08747_ ), .A3(_08749_ ), .ZN(_08750_ ) );
XOR2_X1 _15261_ ( .A(\exu.add.io_rs1_data [23] ), .B(\exu._GEN_0 [23] ), .Z(_08751_ ) );
XOR2_X1 _15262_ ( .A(\exu.add.io_rs1_data [22] ), .B(\exu._GEN_0 [22] ), .Z(_08752_ ) );
NOR2_X1 _15263_ ( .A1(_08751_ ), .A2(_08752_ ), .ZN(_08753_ ) );
XOR2_X1 _15264_ ( .A(\exu.add.io_rs1_data [20] ), .B(\exu._GEN_0 [20] ), .Z(_08754_ ) );
AND2_X1 _15265_ ( .A1(\exu.add.io_rs1_data [21] ), .A2(\exu._GEN_0 [21] ), .ZN(_08755_ ) );
NOR2_X1 _15266_ ( .A1(\exu.add.io_rs1_data [21] ), .A2(\exu._GEN_0 [21] ), .ZN(_08756_ ) );
NOR2_X1 _15267_ ( .A1(_08755_ ), .A2(_08756_ ), .ZN(_08757_ ) );
NOR2_X1 _15268_ ( .A1(_08754_ ), .A2(_08757_ ), .ZN(_08758_ ) );
AND2_X1 _15269_ ( .A1(_08753_ ), .A2(_08758_ ), .ZN(_08759_ ) );
AND2_X1 _15270_ ( .A1(_08750_ ), .A2(_08759_ ), .ZN(_08760_ ) );
XOR2_X1 _15271_ ( .A(\exu._GEN_0 [31] ), .B(\exu.add.io_rs1_data [31] ), .Z(_08761_ ) );
XOR2_X1 _15272_ ( .A(\exu.add.io_rs1_data [30] ), .B(\exu._GEN_0 [30] ), .Z(_08762_ ) );
NOR2_X1 _15273_ ( .A1(_08761_ ), .A2(_08762_ ), .ZN(_08763_ ) );
XOR2_X1 _15274_ ( .A(\exu.add.io_rs1_data [29] ), .B(\exu._GEN_0 [29] ), .Z(_08764_ ) );
XOR2_X1 _15275_ ( .A(\exu.add.io_rs1_data [28] ), .B(\exu._GEN_0 [28] ), .Z(_08765_ ) );
NOR2_X1 _15276_ ( .A1(_08764_ ), .A2(_08765_ ), .ZN(_08766_ ) );
AND2_X1 _15277_ ( .A1(_08763_ ), .A2(_08766_ ), .ZN(_08767_ ) );
XOR2_X1 _15278_ ( .A(\exu.add.io_rs1_data [25] ), .B(\exu._GEN_0 [25] ), .Z(_08768_ ) );
XOR2_X1 _15279_ ( .A(\exu.add.io_rs1_data [24] ), .B(\exu._GEN_0 [24] ), .Z(_08769_ ) );
NOR2_X1 _15280_ ( .A1(_08768_ ), .A2(_08769_ ), .ZN(_08770_ ) );
XOR2_X1 _15281_ ( .A(\exu.add.io_rs1_data [27] ), .B(\exu._GEN_0 [27] ), .Z(_08771_ ) );
XOR2_X1 _15282_ ( .A(\exu.add.io_rs1_data [26] ), .B(\exu._GEN_0 [26] ), .Z(_08772_ ) );
NOR2_X1 _15283_ ( .A1(_08771_ ), .A2(_08772_ ), .ZN(_08773_ ) );
AND2_X1 _15284_ ( .A1(_08770_ ), .A2(_08773_ ), .ZN(_08774_ ) );
AND2_X1 _15285_ ( .A1(_08767_ ), .A2(_08774_ ), .ZN(_08775_ ) );
AND2_X1 _15286_ ( .A1(_08760_ ), .A2(_08775_ ), .ZN(_08776_ ) );
NAND2_X1 _15287_ ( .A1(_08742_ ), .A2(_08776_ ), .ZN(_08777_ ) );
XOR2_X2 _15288_ ( .A(\exu.add.io_rs1_data [1] ), .B(\exu._GEN_0 [1] ), .Z(_08778_ ) );
XOR2_X1 _15289_ ( .A(\exu.add.io_rs1_data [2] ), .B(\exu._GEN_0 [2] ), .Z(_08779_ ) );
OR2_X1 _15290_ ( .A1(_08778_ ), .A2(_08779_ ), .ZN(_08780_ ) );
NOR2_X2 _15291_ ( .A1(_08777_ ), .A2(_08780_ ), .ZN(_08781_ ) );
INV_X1 _15292_ ( .A(\exu.beq.io_is ), .ZN(_08782_ ) );
NOR2_X1 _15293_ ( .A1(_08782_ ), .A2(fanout_net_17 ), .ZN(_08783_ ) );
AND2_X2 _15294_ ( .A1(_08781_ ), .A2(_08783_ ), .ZN(_08784_ ) );
INV_X1 _15295_ ( .A(_08784_ ), .ZN(_08785_ ) );
CLKBUF_X2 _15296_ ( .A(_08785_ ), .Z(_08786_ ) );
OR2_X1 _15297_ ( .A1(_08697_ ), .A2(_08786_ ), .ZN(_08787_ ) );
BUF_X4 _15298_ ( .A(_08782_ ), .Z(_08788_ ) );
NOR2_X1 _15299_ ( .A1(_08784_ ), .A2(_08788_ ), .ZN(_08789_ ) );
INV_X1 _15300_ ( .A(_08789_ ), .ZN(_08790_ ) );
AND2_X1 _15301_ ( .A1(\exu.auipc.io_rs1_data [3] ), .A2(\exu.auipc.io_rs1_data [2] ), .ZN(_08791_ ) );
AND2_X1 _15302_ ( .A1(\exu.auipc.io_rs1_data [5] ), .A2(\exu.auipc.io_rs1_data [4] ), .ZN(_08792_ ) );
AND2_X1 _15303_ ( .A1(_08791_ ), .A2(_08792_ ), .ZN(_08793_ ) );
AND2_X1 _15304_ ( .A1(\exu.auipc.io_rs1_data [7] ), .A2(\exu.auipc.io_rs1_data [6] ), .ZN(_08794_ ) );
AND2_X1 _15305_ ( .A1(_08793_ ), .A2(_08794_ ), .ZN(_08795_ ) );
INV_X1 _15306_ ( .A(_08795_ ), .ZN(_08796_ ) );
NAND2_X1 _15307_ ( .A1(\exu.auipc.io_rs1_data [9] ), .A2(\exu.auipc.io_rs1_data [8] ), .ZN(_08797_ ) );
NOR2_X1 _15308_ ( .A1(_08796_ ), .A2(_08797_ ), .ZN(_08798_ ) );
NAND2_X1 _15309_ ( .A1(\exu.auipc.io_rs1_data [11] ), .A2(\exu.auipc.io_rs1_data [10] ), .ZN(_08799_ ) );
INV_X1 _15310_ ( .A(\exu.auipc.io_rs1_data [12] ), .ZN(_08800_ ) );
NOR3_X1 _15311_ ( .A1(_08799_ ), .A2(_08648_ ), .A3(_08800_ ), .ZN(_08801_ ) );
AND2_X1 _15312_ ( .A1(\exu.auipc.io_rs1_data [15] ), .A2(\exu.auipc.io_rs1_data [14] ), .ZN(_08802_ ) );
AND4_X1 _15313_ ( .A1(\exu.auipc.io_rs1_data [17] ), .A2(_08801_ ), .A3(\exu.auipc.io_rs1_data [16] ), .A4(_08802_ ), .ZN(_08803_ ) );
AND2_X1 _15314_ ( .A1(_08798_ ), .A2(_08803_ ), .ZN(_08804_ ) );
AND4_X1 _15315_ ( .A1(\exu.auipc.io_rs1_data [22] ), .A2(\exu.auipc.io_rs1_data [23] ), .A3(\exu.auipc.io_rs1_data [24] ), .A4(\exu.auipc.io_rs1_data [25] ), .ZN(_08805_ ) );
AND2_X1 _15316_ ( .A1(\exu.auipc.io_rs1_data [19] ), .A2(\exu.auipc.io_rs1_data [18] ), .ZN(_08806_ ) );
AND4_X1 _15317_ ( .A1(\exu.auipc.io_rs1_data [21] ), .A2(_08805_ ), .A3(\exu.auipc.io_rs1_data [20] ), .A4(_08806_ ), .ZN(_08807_ ) );
AND2_X1 _15318_ ( .A1(_08804_ ), .A2(_08807_ ), .ZN(_08808_ ) );
OR2_X1 _15319_ ( .A1(_08808_ ), .A2(_08703_ ), .ZN(_08809_ ) );
NAND3_X1 _15320_ ( .A1(_08804_ ), .A2(_08703_ ), .A3(_08807_ ), .ZN(_08810_ ) );
AND2_X1 _15321_ ( .A1(_08809_ ), .A2(_08810_ ), .ZN(_08811_ ) );
INV_X1 _15322_ ( .A(\exu.bne.io_is ), .ZN(_08812_ ) );
NOR2_X1 _15323_ ( .A1(_08812_ ), .A2(fanout_net_17 ), .ZN(_08813_ ) );
INV_X1 _15324_ ( .A(_08813_ ), .ZN(_08814_ ) );
NOR2_X2 _15325_ ( .A1(_08781_ ), .A2(_08814_ ), .ZN(_08815_ ) );
NOR3_X1 _15326_ ( .A1(_08815_ ), .A2(_08811_ ), .A3(_08812_ ), .ZN(_08816_ ) );
INV_X1 _15327_ ( .A(_08697_ ), .ZN(_08817_ ) );
INV_X1 _15328_ ( .A(_08726_ ), .ZN(_08818_ ) );
INV_X1 _15329_ ( .A(\exu.add.io_rs1_data [2] ), .ZN(_08819_ ) );
NOR2_X1 _15330_ ( .A1(_08819_ ), .A2(\exu._GEN_0 [2] ), .ZN(_08820_ ) );
INV_X1 _15331_ ( .A(\exu.add.io_rs1_data [0] ), .ZN(_08821_ ) );
AOI21_X1 _15332_ ( .A(_08778_ ), .B1(_08821_ ), .B2(\exu._GEN_0 [0] ), .ZN(_08822_ ) );
INV_X1 _15333_ ( .A(\exu._GEN_0 [1] ), .ZN(_08823_ ) );
AOI21_X1 _15334_ ( .A(_08822_ ), .B1(\exu.add.io_rs1_data [1] ), .B2(_08823_ ), .ZN(_08824_ ) );
NOR2_X1 _15335_ ( .A1(_08824_ ), .A2(_08779_ ), .ZN(_08825_ ) );
INV_X1 _15336_ ( .A(\exu._GEN_0 [3] ), .ZN(_08826_ ) );
AOI211_X1 _15337_ ( .A(_08820_ ), .B(_08825_ ), .C1(\exu.add.io_rs1_data [3] ), .C2(_08826_ ), .ZN(_08827_ ) );
NOR2_X1 _15338_ ( .A1(_08826_ ), .A2(\exu.add.io_rs1_data [3] ), .ZN(_08828_ ) );
NOR2_X2 _15339_ ( .A1(_08827_ ), .A2(_08828_ ), .ZN(_08829_ ) );
NAND2_X1 _15340_ ( .A1(_08829_ ), .A2(_08737_ ), .ZN(_08830_ ) );
INV_X1 _15341_ ( .A(\exu.add.io_rs1_data [6] ), .ZN(_08831_ ) );
NOR3_X1 _15342_ ( .A1(_08730_ ), .A2(_08831_ ), .A3(\exu._GEN_0 [6] ), .ZN(_08832_ ) );
INV_X1 _15343_ ( .A(\exu._GEN_0 [7] ), .ZN(_08833_ ) );
INV_X1 _15344_ ( .A(\exu.add.io_rs1_data [4] ), .ZN(_08834_ ) );
NOR3_X1 _15345_ ( .A1(_08735_ ), .A2(_08834_ ), .A3(\exu._GEN_0 [4] ), .ZN(_08835_ ) );
INV_X1 _15346_ ( .A(\exu._GEN_0 [5] ), .ZN(_08836_ ) );
AOI21_X1 _15347_ ( .A(_08835_ ), .B1(\exu.add.io_rs1_data [5] ), .B2(_08836_ ), .ZN(_08837_ ) );
INV_X1 _15348_ ( .A(_08837_ ), .ZN(_08838_ ) );
AOI221_X4 _15349_ ( .A(_08832_ ), .B1(\exu.add.io_rs1_data [7] ), .B2(_08833_ ), .C1(_08838_ ), .C2(_08731_ ), .ZN(_08839_ ) );
AOI21_X4 _15350_ ( .A(_08818_ ), .B1(_08830_ ), .B2(_08839_ ), .ZN(_08840_ ) );
INV_X1 _15351_ ( .A(\exu.add.io_rs1_data [8] ), .ZN(_08841_ ) );
NOR2_X1 _15352_ ( .A1(_08841_ ), .A2(\exu._GEN_0 [8] ), .ZN(_08842_ ) );
INV_X1 _15353_ ( .A(_08842_ ), .ZN(_08843_ ) );
NOR2_X1 _15354_ ( .A1(_08712_ ), .A2(_08843_ ), .ZN(_08844_ ) );
INV_X1 _15355_ ( .A(\exu._GEN_0 [9] ), .ZN(_08845_ ) );
AOI21_X1 _15356_ ( .A(_08844_ ), .B1(\exu.add.io_rs1_data [9] ), .B2(_08845_ ), .ZN(_08846_ ) );
INV_X1 _15357_ ( .A(_08709_ ), .ZN(_08847_ ) );
INV_X1 _15358_ ( .A(\exu.add.io_rs1_data [11] ), .ZN(_08848_ ) );
OAI22_X1 _15359_ ( .A1(_08846_ ), .A2(_08847_ ), .B1(_08848_ ), .B2(\exu._GEN_0 [11] ), .ZN(_08849_ ) );
INV_X1 _15360_ ( .A(\exu.add.io_rs1_data [10] ), .ZN(_08850_ ) );
NOR3_X1 _15361_ ( .A1(_08708_ ), .A2(_08850_ ), .A3(\exu._GEN_0 [10] ), .ZN(_08851_ ) );
NOR2_X1 _15362_ ( .A1(_08849_ ), .A2(_08851_ ), .ZN(_08852_ ) );
INV_X1 _15363_ ( .A(_08725_ ), .ZN(_08853_ ) );
NOR2_X1 _15364_ ( .A1(_08852_ ), .A2(_08853_ ), .ZN(_08854_ ) );
INV_X1 _15365_ ( .A(\exu.add.io_rs1_data [12] ), .ZN(_08855_ ) );
NOR3_X1 _15366_ ( .A1(_08723_ ), .A2(_08855_ ), .A3(\exu._GEN_0 [12] ), .ZN(_08856_ ) );
INV_X1 _15367_ ( .A(\exu._GEN_0 [13] ), .ZN(_08857_ ) );
AOI21_X1 _15368_ ( .A(_08856_ ), .B1(\exu.add.io_rs1_data [13] ), .B2(_08857_ ), .ZN(_08858_ ) );
NOR3_X1 _15369_ ( .A1(_08858_ ), .A2(_08717_ ), .A3(_08718_ ), .ZN(_08859_ ) );
INV_X1 _15370_ ( .A(\exu.add.io_rs1_data [14] ), .ZN(_08860_ ) );
NOR3_X1 _15371_ ( .A1(_08717_ ), .A2(_08860_ ), .A3(\exu._GEN_0 [14] ), .ZN(_08861_ ) );
INV_X1 _15372_ ( .A(\exu.add.io_rs1_data [15] ), .ZN(_08862_ ) );
NOR2_X1 _15373_ ( .A1(_08862_ ), .A2(\exu._GEN_0 [15] ), .ZN(_08863_ ) );
NOR4_X1 _15374_ ( .A1(_08854_ ), .A2(_08859_ ), .A3(_08861_ ), .A4(_08863_ ), .ZN(_08864_ ) );
INV_X1 _15375_ ( .A(_08864_ ), .ZN(_08865_ ) );
OAI21_X1 _15376_ ( .A(_08776_ ), .B1(_08840_ ), .B2(_08865_ ), .ZN(_08866_ ) );
INV_X1 _15377_ ( .A(\exu.add.io_rs1_data [28] ), .ZN(_08867_ ) );
NOR3_X1 _15378_ ( .A1(_08764_ ), .A2(_08867_ ), .A3(\exu._GEN_0 [28] ), .ZN(_08868_ ) );
INV_X1 _15379_ ( .A(\exu.add.io_rs1_data [29] ), .ZN(_08869_ ) );
NOR2_X1 _15380_ ( .A1(_08869_ ), .A2(\exu._GEN_0 [29] ), .ZN(_08870_ ) );
OAI21_X1 _15381_ ( .A(_08763_ ), .B1(_08868_ ), .B2(_08870_ ), .ZN(_08871_ ) );
INV_X1 _15382_ ( .A(\exu._GEN_0 [30] ), .ZN(_08872_ ) );
NAND2_X1 _15383_ ( .A1(_08872_ ), .A2(\exu.add.io_rs1_data [30] ), .ZN(_08873_ ) );
OR2_X1 _15384_ ( .A1(_08761_ ), .A2(_08873_ ), .ZN(_08874_ ) );
INV_X1 _15385_ ( .A(\exu.add.io_rs1_data [31] ), .ZN(_08875_ ) );
OAI211_X1 _15386_ ( .A(_08871_ ), .B(_08874_ ), .C1(\exu._GEN_0 [31] ), .C2(_08875_ ), .ZN(_08876_ ) );
INV_X1 _15387_ ( .A(\exu.add.io_rs1_data [16] ), .ZN(_08877_ ) );
NOR3_X1 _15388_ ( .A1(_08746_ ), .A2(_08877_ ), .A3(\exu._GEN_0 [16] ), .ZN(_08878_ ) );
INV_X1 _15389_ ( .A(\exu._GEN_0 [17] ), .ZN(_08879_ ) );
AOI21_X1 _15390_ ( .A(_08878_ ), .B1(\exu.add.io_rs1_data [17] ), .B2(_08879_ ), .ZN(_08880_ ) );
INV_X1 _15391_ ( .A(_08745_ ), .ZN(_08881_ ) );
INV_X1 _15392_ ( .A(\exu.add.io_rs1_data [19] ), .ZN(_08882_ ) );
OAI22_X1 _15393_ ( .A1(_08880_ ), .A2(_08881_ ), .B1(_08882_ ), .B2(\exu._GEN_0 [19] ), .ZN(_08883_ ) );
INV_X1 _15394_ ( .A(\exu.add.io_rs1_data [18] ), .ZN(_08884_ ) );
NOR3_X1 _15395_ ( .A1(_08743_ ), .A2(_08884_ ), .A3(\exu._GEN_0 [18] ), .ZN(_08885_ ) );
OAI21_X1 _15396_ ( .A(_08759_ ), .B1(_08883_ ), .B2(_08885_ ), .ZN(_08886_ ) );
INV_X1 _15397_ ( .A(\exu.add.io_rs1_data [22] ), .ZN(_08887_ ) );
NOR2_X1 _15398_ ( .A1(_08887_ ), .A2(\exu._GEN_0 [22] ), .ZN(_08888_ ) );
INV_X1 _15399_ ( .A(_08888_ ), .ZN(_08889_ ) );
OR2_X1 _15400_ ( .A1(_08751_ ), .A2(_08889_ ), .ZN(_08890_ ) );
INV_X1 _15401_ ( .A(\exu.add.io_rs1_data [20] ), .ZN(_08891_ ) );
NOR2_X1 _15402_ ( .A1(_08891_ ), .A2(\exu._GEN_0 [20] ), .ZN(_08892_ ) );
INV_X1 _15403_ ( .A(_08892_ ), .ZN(_08893_ ) );
NOR2_X1 _15404_ ( .A1(_08757_ ), .A2(_08893_ ), .ZN(_08894_ ) );
INV_X1 _15405_ ( .A(\exu._GEN_0 [21] ), .ZN(_08895_ ) );
AOI21_X1 _15406_ ( .A(_08894_ ), .B1(\exu.add.io_rs1_data [21] ), .B2(_08895_ ), .ZN(_08896_ ) );
INV_X1 _15407_ ( .A(_08896_ ), .ZN(_08897_ ) );
INV_X1 _15408_ ( .A(\exu._GEN_0 [23] ), .ZN(_08898_ ) );
AOI22_X1 _15409_ ( .A1(_08897_ ), .A2(_08753_ ), .B1(\exu.add.io_rs1_data [23] ), .B2(_08898_ ), .ZN(_08899_ ) );
AND3_X1 _15410_ ( .A1(_08886_ ), .A2(_08890_ ), .A3(_08899_ ), .ZN(_08900_ ) );
INV_X1 _15411_ ( .A(_08775_ ), .ZN(_08901_ ) );
NOR2_X1 _15412_ ( .A1(_08900_ ), .A2(_08901_ ), .ZN(_08902_ ) );
INV_X1 _15413_ ( .A(\exu.add.io_rs1_data [24] ), .ZN(_08903_ ) );
NOR2_X1 _15414_ ( .A1(_08903_ ), .A2(\exu._GEN_0 [24] ), .ZN(_08904_ ) );
INV_X1 _15415_ ( .A(_08904_ ), .ZN(_08905_ ) );
NOR2_X1 _15416_ ( .A1(_08768_ ), .A2(_08905_ ), .ZN(_08906_ ) );
INV_X1 _15417_ ( .A(_08906_ ), .ZN(_08907_ ) );
INV_X1 _15418_ ( .A(\exu.add.io_rs1_data [25] ), .ZN(_08908_ ) );
OAI21_X1 _15419_ ( .A(_08907_ ), .B1(_08908_ ), .B2(\exu._GEN_0 [25] ), .ZN(_08909_ ) );
AND2_X1 _15420_ ( .A1(_08909_ ), .A2(_08773_ ), .ZN(_08910_ ) );
INV_X1 _15421_ ( .A(\exu.add.io_rs1_data [26] ), .ZN(_08911_ ) );
NOR3_X1 _15422_ ( .A1(_08771_ ), .A2(_08911_ ), .A3(\exu._GEN_0 [26] ), .ZN(_08912_ ) );
INV_X1 _15423_ ( .A(\exu.add.io_rs1_data [27] ), .ZN(_08913_ ) );
NOR2_X1 _15424_ ( .A1(_08913_ ), .A2(\exu._GEN_0 [27] ), .ZN(_08914_ ) );
NOR3_X1 _15425_ ( .A1(_08910_ ), .A2(_08912_ ), .A3(_08914_ ), .ZN(_08915_ ) );
INV_X1 _15426_ ( .A(_08915_ ), .ZN(_08916_ ) );
AOI211_X1 _15427_ ( .A(_08876_ ), .B(_08902_ ), .C1(_08767_ ), .C2(_08916_ ), .ZN(_08917_ ) );
AND2_X2 _15428_ ( .A1(_08866_ ), .A2(_08917_ ), .ZN(_08918_ ) );
INV_X1 _15429_ ( .A(_08761_ ), .ZN(_08919_ ) );
XNOR2_X2 _15430_ ( .A(_08918_ ), .B(_08919_ ), .ZN(_08920_ ) );
INV_X1 _15431_ ( .A(_08920_ ), .ZN(_08921_ ) );
INV_X1 _15432_ ( .A(\exu.bge.io_is ), .ZN(_08922_ ) );
NOR2_X1 _15433_ ( .A1(_08922_ ), .A2(fanout_net_17 ), .ZN(_08923_ ) );
AND2_X2 _15434_ ( .A1(_08921_ ), .A2(_08923_ ), .ZN(_08924_ ) );
BUF_X4 _15435_ ( .A(_08924_ ), .Z(_08925_ ) );
INV_X1 _15436_ ( .A(_08925_ ), .ZN(_08926_ ) );
OR2_X1 _15437_ ( .A1(_08697_ ), .A2(_08926_ ), .ZN(_08927_ ) );
NOR2_X4 _15438_ ( .A1(_08925_ ), .A2(_08922_ ), .ZN(_08928_ ) );
INV_X1 _15439_ ( .A(_08928_ ), .ZN(_08929_ ) );
BUF_X4 _15440_ ( .A(_08929_ ), .Z(_08930_ ) );
INV_X2 _15441_ ( .A(\exu.bgeu.io_is ), .ZN(_08931_ ) );
NOR2_X1 _15442_ ( .A1(_08931_ ), .A2(fanout_net_17 ), .ZN(_08932_ ) );
INV_X1 _15443_ ( .A(_08932_ ), .ZN(_08933_ ) );
NOR2_X1 _15444_ ( .A1(_08918_ ), .A2(_08933_ ), .ZN(_08934_ ) );
BUF_X4 _15445_ ( .A(_08934_ ), .Z(_08935_ ) );
INV_X1 _15446_ ( .A(_08935_ ), .ZN(_08936_ ) );
NOR2_X1 _15447_ ( .A1(_08697_ ), .A2(_08936_ ), .ZN(_08937_ ) );
NOR2_X1 _15448_ ( .A1(_08934_ ), .A2(_08931_ ), .ZN(_08938_ ) );
INV_X1 _15449_ ( .A(_08811_ ), .ZN(_08939_ ) );
INV_X1 _15450_ ( .A(fanout_net_7 ), .ZN(_08940_ ) );
NOR2_X1 _15451_ ( .A1(_08940_ ), .A2(fanout_net_17 ), .ZN(_08941_ ) );
AND2_X1 _15452_ ( .A1(_08918_ ), .A2(_08941_ ), .ZN(_08942_ ) );
BUF_X2 _15453_ ( .A(_08942_ ), .Z(_08943_ ) );
NAND2_X1 _15454_ ( .A1(_08697_ ), .A2(_08943_ ), .ZN(_08944_ ) );
BUF_X4 _15455_ ( .A(_08943_ ), .Z(_08945_ ) );
OAI211_X1 _15456_ ( .A(_08944_ ), .B(fanout_net_7 ), .C1(_08945_ ), .C2(_08939_ ), .ZN(_08946_ ) );
INV_X1 _15457_ ( .A(fanout_net_6 ), .ZN(_08947_ ) );
AND3_X1 _15458_ ( .A1(fanout_net_17 ), .A2(fanout_net_11 ), .A3(\exu.addi._io_rd_T_4_$_NOT__Y_5_A_$_MUX__A_B ), .ZN(_08948_ ) );
INV_X1 _15459_ ( .A(fanout_net_11 ), .ZN(_08949_ ) );
NAND3_X1 _15460_ ( .A1(_08809_ ), .A2(exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ), .A3(_08810_ ), .ZN(_08950_ ) );
AND3_X1 _15461_ ( .A1(\exu.csrrs.io_csr_rdata [3] ), .A2(\exu.csrrs.io_csr_rdata [2] ), .A3(\exu.csrrs.io_csr_rdata [4] ), .ZN(_08951_ ) );
NAND3_X1 _15462_ ( .A1(_08951_ ), .A2(\exu.csrrs.io_csr_rdata [6] ), .A3(\exu.csrrs.io_csr_rdata [5] ), .ZN(_08952_ ) );
INV_X1 _15463_ ( .A(\exu.csrrs.io_csr_rdata [7] ), .ZN(_08953_ ) );
NOR2_X1 _15464_ ( .A1(_08952_ ), .A2(_08953_ ), .ZN(_08954_ ) );
NAND2_X1 _15465_ ( .A1(_08954_ ), .A2(\exu.csrrs.io_csr_rdata [8] ), .ZN(_08955_ ) );
INV_X1 _15466_ ( .A(\exu.csrrs.io_csr_rdata [9] ), .ZN(_08956_ ) );
NOR2_X1 _15467_ ( .A1(_08955_ ), .A2(_08956_ ), .ZN(_08957_ ) );
NAND4_X1 _15468_ ( .A1(\exu.csrrs.io_csr_rdata [16] ), .A2(\exu.csrrs.io_csr_rdata [14] ), .A3(\exu.csrrs.io_csr_rdata [15] ), .A4(\exu.csrrs.io_csr_rdata [17] ), .ZN(_08958_ ) );
NAND2_X1 _15469_ ( .A1(\exu.csrrs.io_csr_rdata [12] ), .A2(\exu.csrrs.io_csr_rdata [13] ), .ZN(_08959_ ) );
INV_X1 _15470_ ( .A(\exu.csrrs.io_csr_rdata [11] ), .ZN(_08960_ ) );
INV_X1 _15471_ ( .A(\exu.csrrs.io_csr_rdata [10] ), .ZN(_08961_ ) );
NOR4_X1 _15472_ ( .A1(_08958_ ), .A2(_08959_ ), .A3(_08960_ ), .A4(_08961_ ), .ZN(_08962_ ) );
AND2_X1 _15473_ ( .A1(_08957_ ), .A2(_08962_ ), .ZN(_08963_ ) );
AND2_X1 _15474_ ( .A1(\exu.csrrs.io_csr_rdata [18] ), .A2(\exu.csrrs.io_csr_rdata [19] ), .ZN(_08964_ ) );
AND3_X1 _15475_ ( .A1(_08964_ ), .A2(\exu.csrrs.io_csr_rdata [20] ), .A3(\exu.csrrs.io_csr_rdata [21] ), .ZN(_08965_ ) );
AND2_X1 _15476_ ( .A1(\exu.csrrs.io_csr_rdata [25] ), .A2(\exu.csrrs.io_csr_rdata [24] ), .ZN(_08966_ ) );
AND2_X1 _15477_ ( .A1(\exu.csrrs.io_csr_rdata [22] ), .A2(\exu.csrrs.io_csr_rdata [23] ), .ZN(_08967_ ) );
AND3_X1 _15478_ ( .A1(_08965_ ), .A2(_08966_ ), .A3(_08967_ ), .ZN(_08968_ ) );
AND2_X1 _15479_ ( .A1(_08963_ ), .A2(_08968_ ), .ZN(_08969_ ) );
XOR2_X1 _15480_ ( .A(_08969_ ), .B(\ifu.io_out_bits_pc_$_NOT__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ), .Z(_08970_ ) );
NOR2_X1 _15481_ ( .A1(_08949_ ), .A2(fanout_net_17 ), .ZN(_08971_ ) );
BUF_X4 _15482_ ( .A(_08971_ ), .Z(_08972_ ) );
AOI221_X4 _15483_ ( .A(_08948_ ), .B1(_08949_ ), .B2(_08950_ ), .C1(_08970_ ), .C2(_08972_ ), .ZN(_08973_ ) );
OAI211_X1 _15484_ ( .A(_08946_ ), .B(_08947_ ), .C1(fanout_net_7 ), .C2(_08973_ ), .ZN(_08974_ ) );
NOR2_X1 _15485_ ( .A1(_08947_ ), .A2(fanout_net_17 ), .ZN(_08975_ ) );
AND2_X2 _15486_ ( .A1(_08920_ ), .A2(_08975_ ), .ZN(_08976_ ) );
INV_X1 _15487_ ( .A(_08976_ ), .ZN(_08977_ ) );
INV_X1 _15488_ ( .A(fanout_net_17 ), .ZN(_08978_ ) );
AND2_X1 _15489_ ( .A1(_08920_ ), .A2(_08978_ ), .ZN(_08979_ ) );
OAI22_X1 _15490_ ( .A1(_08817_ ), .A2(_08977_ ), .B1(_08979_ ), .B2(_08939_ ), .ZN(_08980_ ) );
AOI21_X1 _15491_ ( .A(\exu.bgeu.io_is ), .B1(_08980_ ), .B2(fanout_net_6 ), .ZN(_08981_ ) );
AOI221_X4 _15492_ ( .A(_08937_ ), .B1(_08938_ ), .B2(_08939_ ), .C1(_08974_ ), .C2(_08981_ ), .ZN(_08982_ ) );
OAI221_X1 _15493_ ( .A(_08927_ ), .B1(_08930_ ), .B2(_08811_ ), .C1(_08982_ ), .C2(\exu.bge.io_is ), .ZN(_08983_ ) );
BUF_X4 _15494_ ( .A(_08812_ ), .Z(_08984_ ) );
AOI221_X4 _15495_ ( .A(_08816_ ), .B1(_08815_ ), .B2(_08817_ ), .C1(_08983_ ), .C2(_08984_ ), .ZN(_08985_ ) );
OAI221_X1 _15496_ ( .A(_08787_ ), .B1(_08790_ ), .B2(_08811_ ), .C1(_08985_ ), .C2(\exu.beq.io_is ), .ZN(_08986_ ) );
AOI221_X4 _15497_ ( .A(fanout_net_8 ), .B1(_08701_ ), .B2(_08704_ ), .C1(_08986_ ), .C2(_08702_ ), .ZN(_08987_ ) );
INV_X1 _15498_ ( .A(fanout_net_8 ), .ZN(_08988_ ) );
BUF_X4 _15499_ ( .A(_08988_ ), .Z(_08989_ ) );
NOR2_X1 _15500_ ( .A1(_08989_ ), .A2(fanout_net_17 ), .ZN(_08990_ ) );
BUF_X4 _15501_ ( .A(_08990_ ), .Z(_08991_ ) );
AOI211_X1 _15502_ ( .A(fanout_net_10 ), .B(_08987_ ), .C1(\exu.csrrs.io_csr_rdata [26] ), .C2(_08991_ ), .ZN(_08992_ ) );
XNOR2_X1 _15503_ ( .A(\exu.auipc.io_rs1_data [22] ), .B(\idu.io_in_bits_pc [22] ), .ZN(_08993_ ) );
XNOR2_X1 _15504_ ( .A(\exu.auipc.io_rs1_data [23] ), .B(\idu.io_in_bits_pc [23] ), .ZN(_08994_ ) );
XNOR2_X1 _15505_ ( .A(\exu.auipc.io_rs1_data [19] ), .B(\idu.io_in_bits_pc [19] ), .ZN(_08995_ ) );
XNOR2_X1 _15506_ ( .A(\exu.auipc.io_rs1_data [18] ), .B(\idu.io_in_bits_pc [18] ), .ZN(_08996_ ) );
AND4_X1 _15507_ ( .A1(_08993_ ), .A2(_08994_ ), .A3(_08995_ ), .A4(_08996_ ), .ZN(_08997_ ) );
XNOR2_X1 _15508_ ( .A(\exu.auipc.io_rs1_data [29] ), .B(\idu.io_in_bits_pc [29] ), .ZN(_08998_ ) );
XNOR2_X1 _15509_ ( .A(\exu.auipc.io_rs1_data [25] ), .B(\idu.io_in_bits_pc [25] ), .ZN(_08999_ ) );
XNOR2_X1 _15510_ ( .A(\exu.auipc.io_rs1_data [28] ), .B(\idu.io_in_bits_pc [28] ), .ZN(_09000_ ) );
XNOR2_X1 _15511_ ( .A(\exu.auipc.io_rs1_data [24] ), .B(\idu.io_in_bits_pc [24] ), .ZN(_09001_ ) );
AND4_X1 _15512_ ( .A1(_08998_ ), .A2(_08999_ ), .A3(_09000_ ), .A4(_09001_ ), .ZN(_09002_ ) );
XNOR2_X1 _15513_ ( .A(\exu.auipc.io_rs1_data [4] ), .B(\idu.io_in_bits_pc [4] ), .ZN(_09003_ ) );
XNOR2_X1 _15514_ ( .A(\exu.auipc.io_rs1_data [5] ), .B(\idu.io_in_bits_pc [5] ), .ZN(_09004_ ) );
XNOR2_X1 _15515_ ( .A(\exu.auipc.io_rs1_data [1] ), .B(\idu.io_in_bits_pc [1] ), .ZN(_09005_ ) );
XNOR2_X1 _15516_ ( .A(\exu.auipc.io_rs1_data [0] ), .B(\idu.io_in_bits_pc [0] ), .ZN(_09006_ ) );
AND4_X1 _15517_ ( .A1(_09003_ ), .A2(_09004_ ), .A3(_09005_ ), .A4(_09006_ ), .ZN(_09007_ ) );
XNOR2_X1 _15518_ ( .A(\exu.auipc.io_rs1_data [11] ), .B(\idu.io_in_bits_pc [11] ), .ZN(_09008_ ) );
XNOR2_X1 _15519_ ( .A(\exu.auipc.io_rs1_data [15] ), .B(\idu.io_in_bits_pc [15] ), .ZN(_09009_ ) );
XNOR2_X1 _15520_ ( .A(\exu.auipc.io_rs1_data [14] ), .B(\idu.io_in_bits_pc [14] ), .ZN(_09010_ ) );
XNOR2_X1 _15521_ ( .A(\exu.auipc.io_rs1_data [10] ), .B(\idu.io_in_bits_pc [10] ), .ZN(_09011_ ) );
AND4_X1 _15522_ ( .A1(_09008_ ), .A2(_09009_ ), .A3(_09010_ ), .A4(_09011_ ), .ZN(_09012_ ) );
AND4_X1 _15523_ ( .A1(_08997_ ), .A2(_09002_ ), .A3(_09007_ ), .A4(_09012_ ), .ZN(_09013_ ) );
XNOR2_X1 _15524_ ( .A(\exu.auipc.io_rs1_data [21] ), .B(\idu.io_in_bits_pc [21] ), .ZN(_09014_ ) );
XNOR2_X1 _15525_ ( .A(\exu.auipc.io_rs1_data [17] ), .B(\idu.io_in_bits_pc [17] ), .ZN(_09015_ ) );
XNOR2_X1 _15526_ ( .A(\exu.auipc.io_rs1_data [20] ), .B(\idu.io_in_bits_pc [20] ), .ZN(_09016_ ) );
XNOR2_X1 _15527_ ( .A(\exu.auipc.io_rs1_data [16] ), .B(\idu.io_in_bits_pc [16] ), .ZN(_09017_ ) );
AND4_X1 _15528_ ( .A1(_09014_ ), .A2(_09015_ ), .A3(_09016_ ), .A4(_09017_ ), .ZN(_09018_ ) );
XNOR2_X1 _15529_ ( .A(\exu.auipc.io_rs1_data [26] ), .B(\idu.io_in_bits_pc [26] ), .ZN(_09019_ ) );
XNOR2_X1 _15530_ ( .A(\exu.auipc.io_rs1_data [27] ), .B(\idu.io_in_bits_pc [27] ), .ZN(_09020_ ) );
XNOR2_X1 _15531_ ( .A(\idu.io_in_bits_pc [31] ), .B(\exu.auipc.io_rs1_data [31] ), .ZN(_09021_ ) );
XNOR2_X1 _15532_ ( .A(\idu.io_in_bits_pc [30] ), .B(\exu.auipc.io_rs1_data [30] ), .ZN(_09022_ ) );
AND4_X1 _15533_ ( .A1(_09019_ ), .A2(_09020_ ), .A3(_09021_ ), .A4(_09022_ ), .ZN(_09023_ ) );
XNOR2_X1 _15534_ ( .A(\exu.auipc.io_rs1_data [6] ), .B(\idu.io_in_bits_pc [6] ), .ZN(_09024_ ) );
XNOR2_X1 _15535_ ( .A(\exu.auipc.io_rs1_data [2] ), .B(\idu.io_in_bits_pc [2] ), .ZN(_09025_ ) );
XNOR2_X1 _15536_ ( .A(\exu.auipc.io_rs1_data [3] ), .B(\idu.io_in_bits_pc [3] ), .ZN(_09026_ ) );
XNOR2_X1 _15537_ ( .A(\exu.auipc.io_rs1_data [7] ), .B(\idu.io_in_bits_pc [7] ), .ZN(_09027_ ) );
AND4_X1 _15538_ ( .A1(_09024_ ), .A2(_09025_ ), .A3(_09026_ ), .A4(_09027_ ), .ZN(_09028_ ) );
XNOR2_X1 _15539_ ( .A(\exu.auipc.io_rs1_data [12] ), .B(\idu.io_in_bits_pc [12] ), .ZN(_09029_ ) );
XNOR2_X1 _15540_ ( .A(\exu.auipc.io_rs1_data [13] ), .B(\idu.io_in_bits_pc [13] ), .ZN(_09030_ ) );
XNOR2_X1 _15541_ ( .A(\exu.auipc.io_rs1_data [9] ), .B(\idu.io_in_bits_pc [9] ), .ZN(_09031_ ) );
XNOR2_X1 _15542_ ( .A(\exu.auipc.io_rs1_data [8] ), .B(\idu.io_in_bits_pc [8] ), .ZN(_09032_ ) );
AND4_X1 _15543_ ( .A1(_09029_ ), .A2(_09030_ ), .A3(_09031_ ), .A4(_09032_ ), .ZN(_09033_ ) );
AND4_X1 _15544_ ( .A1(_09018_ ), .A2(_09023_ ), .A3(_09028_ ), .A4(_09033_ ), .ZN(_09034_ ) );
INV_X1 _15545_ ( .A(exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ), .ZN(_09035_ ) );
BUF_X2 _15546_ ( .A(_09035_ ), .Z(_09036_ ) );
NAND3_X1 _15547_ ( .A1(_09013_ ), .A2(_09034_ ), .A3(_09036_ ), .ZN(_09037_ ) );
NOR2_X1 _15548_ ( .A1(_09037_ ), .A2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_09038_ ) );
INV_X1 _15549_ ( .A(_09038_ ), .ZN(_09039_ ) );
CLKBUF_X2 _15550_ ( .A(_09039_ ), .Z(_09040_ ) );
INV_X1 _15551_ ( .A(fanout_net_10 ), .ZN(_09041_ ) );
BUF_X4 _15552_ ( .A(_09041_ ), .Z(_09042_ ) );
AND2_X1 _15553_ ( .A1(\exu.add.io_rs1_data [19] ), .A2(\exu.addi.io_imm [19] ), .ZN(_09043_ ) );
NOR2_X1 _15554_ ( .A1(\exu.add.io_rs1_data [19] ), .A2(\exu.addi.io_imm [19] ), .ZN(_09044_ ) );
NOR2_X1 _15555_ ( .A1(_09043_ ), .A2(_09044_ ), .ZN(_09045_ ) );
AND2_X1 _15556_ ( .A1(\exu.add.io_rs1_data [18] ), .A2(\exu.addi.io_imm [18] ), .ZN(_09046_ ) );
NOR2_X1 _15557_ ( .A1(\exu.add.io_rs1_data [18] ), .A2(\exu.addi.io_imm [18] ), .ZN(_09047_ ) );
NOR2_X1 _15558_ ( .A1(_09046_ ), .A2(_09047_ ), .ZN(_09048_ ) );
AND2_X1 _15559_ ( .A1(_09045_ ), .A2(_09048_ ), .ZN(_09049_ ) );
XOR2_X1 _15560_ ( .A(\exu.add.io_rs1_data [4] ), .B(\exu.addi.io_imm [4] ), .Z(_09050_ ) );
AND2_X1 _15561_ ( .A1(\exu.add.io_rs1_data [1] ), .A2(\exu.addi.io_imm [1] ), .ZN(_09051_ ) );
INV_X1 _15562_ ( .A(_09051_ ), .ZN(_09052_ ) );
AND2_X1 _15563_ ( .A1(\exu.addi.io_imm [0] ), .A2(\exu.add.io_rs1_data [0] ), .ZN(_09053_ ) );
INV_X1 _15564_ ( .A(_09053_ ), .ZN(_09054_ ) );
NOR2_X1 _15565_ ( .A1(\exu.add.io_rs1_data [1] ), .A2(\exu.addi.io_imm [1] ), .ZN(_09055_ ) );
OAI21_X1 _15566_ ( .A(_09052_ ), .B1(_09054_ ), .B2(_09055_ ), .ZN(_09056_ ) );
AND2_X1 _15567_ ( .A1(\exu.add.io_rs1_data [2] ), .A2(\exu.addi.io_imm [2] ), .ZN(_09057_ ) );
NOR2_X1 _15568_ ( .A1(\exu.add.io_rs1_data [2] ), .A2(\exu.addi.io_imm [2] ), .ZN(_09058_ ) );
NOR2_X1 _15569_ ( .A1(_09057_ ), .A2(_09058_ ), .ZN(_09059_ ) );
NAND2_X1 _15570_ ( .A1(_09056_ ), .A2(_09059_ ), .ZN(_09060_ ) );
AND2_X1 _15571_ ( .A1(\exu.add.io_rs1_data [3] ), .A2(\exu.addi.io_imm [3] ), .ZN(_09061_ ) );
INV_X1 _15572_ ( .A(_09061_ ), .ZN(_09062_ ) );
INV_X1 _15573_ ( .A(_09057_ ), .ZN(_09063_ ) );
NAND3_X1 _15574_ ( .A1(_09060_ ), .A2(_09062_ ), .A3(_09063_ ), .ZN(_09064_ ) );
NOR2_X1 _15575_ ( .A1(\exu.add.io_rs1_data [3] ), .A2(\exu.addi.io_imm [3] ), .ZN(_09065_ ) );
INV_X1 _15576_ ( .A(_09065_ ), .ZN(_09066_ ) );
AND2_X1 _15577_ ( .A1(\exu.add.io_rs1_data [5] ), .A2(\exu.addi.io_imm [5] ), .ZN(_09067_ ) );
NOR2_X1 _15578_ ( .A1(\exu.add.io_rs1_data [5] ), .A2(\exu.addi.io_imm [5] ), .ZN(_09068_ ) );
NOR2_X1 _15579_ ( .A1(_09067_ ), .A2(_09068_ ), .ZN(_09069_ ) );
AND4_X1 _15580_ ( .A1(_09050_ ), .A2(_09064_ ), .A3(_09066_ ), .A4(_09069_ ), .ZN(_09070_ ) );
AND2_X1 _15581_ ( .A1(\exu.add.io_rs1_data [4] ), .A2(\exu.addi.io_imm [4] ), .ZN(_09071_ ) );
AND2_X1 _15582_ ( .A1(_09069_ ), .A2(_09071_ ), .ZN(_09072_ ) );
NOR3_X1 _15583_ ( .A1(_09070_ ), .A2(_09067_ ), .A3(_09072_ ), .ZN(_09073_ ) );
AND2_X1 _15584_ ( .A1(\exu.add.io_rs1_data [6] ), .A2(\exu.addi.io_imm [6] ), .ZN(_09074_ ) );
NOR2_X1 _15585_ ( .A1(\exu.add.io_rs1_data [6] ), .A2(\exu.addi.io_imm [6] ), .ZN(_09075_ ) );
NOR3_X1 _15586_ ( .A1(_09073_ ), .A2(_09074_ ), .A3(_09075_ ), .ZN(_09076_ ) );
AND2_X1 _15587_ ( .A1(\exu.add.io_rs1_data [7] ), .A2(\exu.addi.io_imm [7] ), .ZN(_09077_ ) );
NOR3_X1 _15588_ ( .A1(_09076_ ), .A2(_09077_ ), .A3(_09074_ ), .ZN(_09078_ ) );
NOR2_X1 _15589_ ( .A1(\exu.add.io_rs1_data [7] ), .A2(\exu.addi.io_imm [7] ), .ZN(_09079_ ) );
AND2_X1 _15590_ ( .A1(\exu.add.io_rs1_data [8] ), .A2(\exu.addi.io_imm [8] ), .ZN(_09080_ ) );
NOR2_X1 _15591_ ( .A1(\exu.add.io_rs1_data [8] ), .A2(\exu.addi.io_imm [8] ), .ZN(_09081_ ) );
NOR2_X1 _15592_ ( .A1(_09080_ ), .A2(_09081_ ), .ZN(_09082_ ) );
AND2_X1 _15593_ ( .A1(\exu.addi.io_imm [9] ), .A2(\exu.add.io_rs1_data [9] ), .ZN(_09083_ ) );
NOR2_X1 _15594_ ( .A1(\exu.addi.io_imm [9] ), .A2(\exu.add.io_rs1_data [9] ), .ZN(_09084_ ) );
NOR2_X1 _15595_ ( .A1(_09083_ ), .A2(_09084_ ), .ZN(_09085_ ) );
NAND2_X1 _15596_ ( .A1(_09082_ ), .A2(_09085_ ), .ZN(_09086_ ) );
AND2_X1 _15597_ ( .A1(\exu.add.io_rs1_data [10] ), .A2(\exu.addi.io_imm [10] ), .ZN(_09087_ ) );
NOR2_X1 _15598_ ( .A1(\exu.add.io_rs1_data [10] ), .A2(\exu.addi.io_imm [10] ), .ZN(_09088_ ) );
NOR2_X1 _15599_ ( .A1(_09087_ ), .A2(_09088_ ), .ZN(_09089_ ) );
AND2_X1 _15600_ ( .A1(\exu.add.io_rs1_data [11] ), .A2(\exu.addi.io_imm [11] ), .ZN(_09090_ ) );
NOR2_X1 _15601_ ( .A1(\exu.add.io_rs1_data [11] ), .A2(\exu.addi.io_imm [11] ), .ZN(_09091_ ) );
NOR2_X1 _15602_ ( .A1(_09090_ ), .A2(_09091_ ), .ZN(_09092_ ) );
NAND2_X1 _15603_ ( .A1(_09089_ ), .A2(_09092_ ), .ZN(_09093_ ) );
NOR4_X1 _15604_ ( .A1(_09078_ ), .A2(_09079_ ), .A3(_09086_ ), .A4(_09093_ ), .ZN(_09094_ ) );
INV_X1 _15605_ ( .A(_09084_ ), .ZN(_09095_ ) );
AOI21_X1 _15606_ ( .A(_09083_ ), .B1(_09095_ ), .B2(_09080_ ), .ZN(_09096_ ) );
OR2_X1 _15607_ ( .A1(_09093_ ), .A2(_09096_ ), .ZN(_09097_ ) );
INV_X1 _15608_ ( .A(_09090_ ), .ZN(_09098_ ) );
INV_X1 _15609_ ( .A(_09091_ ), .ZN(_09099_ ) );
NAND3_X1 _15610_ ( .A1(_09098_ ), .A2(_09099_ ), .A3(_09087_ ), .ZN(_09100_ ) );
NAND3_X1 _15611_ ( .A1(_09097_ ), .A2(_09098_ ), .A3(_09100_ ), .ZN(_09101_ ) );
OR2_X1 _15612_ ( .A1(_09094_ ), .A2(_09101_ ), .ZN(_09102_ ) );
AND2_X1 _15613_ ( .A1(\exu.add.io_rs1_data [15] ), .A2(\exu.addi.io_imm [15] ), .ZN(_09103_ ) );
NOR2_X1 _15614_ ( .A1(\exu.add.io_rs1_data [15] ), .A2(\exu.addi.io_imm [15] ), .ZN(_09104_ ) );
NOR2_X1 _15615_ ( .A1(_09103_ ), .A2(_09104_ ), .ZN(_09105_ ) );
AND2_X1 _15616_ ( .A1(\exu.add.io_rs1_data [14] ), .A2(\exu.addi.io_imm [14] ), .ZN(_09106_ ) );
NOR2_X1 _15617_ ( .A1(\exu.add.io_rs1_data [14] ), .A2(\exu.addi.io_imm [14] ), .ZN(_09107_ ) );
NOR2_X1 _15618_ ( .A1(_09106_ ), .A2(_09107_ ), .ZN(_09108_ ) );
AND2_X1 _15619_ ( .A1(\exu.addi.io_imm [13] ), .A2(\exu.add.io_rs1_data [13] ), .ZN(_09109_ ) );
NOR2_X1 _15620_ ( .A1(\exu.addi.io_imm [13] ), .A2(\exu.add.io_rs1_data [13] ), .ZN(_09110_ ) );
NOR2_X1 _15621_ ( .A1(_09109_ ), .A2(_09110_ ), .ZN(_09111_ ) );
AND2_X1 _15622_ ( .A1(\exu.add.io_rs1_data [12] ), .A2(\exu.addi.io_imm [12] ), .ZN(_09112_ ) );
NOR2_X1 _15623_ ( .A1(\exu.add.io_rs1_data [12] ), .A2(\exu.addi.io_imm [12] ), .ZN(_09113_ ) );
NOR2_X1 _15624_ ( .A1(_09112_ ), .A2(_09113_ ), .ZN(_09114_ ) );
AND2_X1 _15625_ ( .A1(_09111_ ), .A2(_09114_ ), .ZN(_09115_ ) );
NAND4_X1 _15626_ ( .A1(_09102_ ), .A2(_09105_ ), .A3(_09108_ ), .A4(_09115_ ), .ZN(_09116_ ) );
AOI21_X1 _15627_ ( .A(_09109_ ), .B1(_09111_ ), .B2(_09112_ ), .ZN(_09117_ ) );
INV_X1 _15628_ ( .A(_09108_ ), .ZN(_09118_ ) );
NOR4_X1 _15629_ ( .A1(_09117_ ), .A2(_09118_ ), .A3(_09103_ ), .A4(_09104_ ), .ZN(_09119_ ) );
INV_X1 _15630_ ( .A(\exu.addi.io_imm [14] ), .ZN(_09120_ ) );
NOR4_X1 _15631_ ( .A1(_09103_ ), .A2(_09104_ ), .A3(_08860_ ), .A4(_09120_ ), .ZN(_09121_ ) );
NOR3_X1 _15632_ ( .A1(_09119_ ), .A2(_09103_ ), .A3(_09121_ ), .ZN(_09122_ ) );
NAND2_X1 _15633_ ( .A1(_09116_ ), .A2(_09122_ ), .ZN(_09123_ ) );
AND2_X1 _15634_ ( .A1(\exu.add.io_rs1_data [16] ), .A2(\exu.addi.io_imm [16] ), .ZN(_09124_ ) );
NOR2_X1 _15635_ ( .A1(\exu.add.io_rs1_data [16] ), .A2(\exu.addi.io_imm [16] ), .ZN(_09125_ ) );
NOR2_X1 _15636_ ( .A1(_09124_ ), .A2(_09125_ ), .ZN(_09126_ ) );
AND2_X1 _15637_ ( .A1(\exu.add.io_rs1_data [17] ), .A2(\exu.addi.io_imm [17] ), .ZN(_09127_ ) );
NOR2_X1 _15638_ ( .A1(\exu.add.io_rs1_data [17] ), .A2(\exu.addi.io_imm [17] ), .ZN(_09128_ ) );
NOR2_X1 _15639_ ( .A1(_09127_ ), .A2(_09128_ ), .ZN(_09129_ ) );
AND4_X1 _15640_ ( .A1(_09049_ ), .A2(_09123_ ), .A3(_09126_ ), .A4(_09129_ ), .ZN(_09130_ ) );
INV_X1 _15641_ ( .A(_09128_ ), .ZN(_09131_ ) );
AOI21_X1 _15642_ ( .A(_09127_ ), .B1(_09131_ ), .B2(_09124_ ), .ZN(_09132_ ) );
INV_X1 _15643_ ( .A(_09048_ ), .ZN(_09133_ ) );
NOR4_X1 _15644_ ( .A1(_09132_ ), .A2(_09133_ ), .A3(_09043_ ), .A4(_09044_ ), .ZN(_09134_ ) );
INV_X1 _15645_ ( .A(\exu.addi.io_imm [18] ), .ZN(_09135_ ) );
NOR3_X1 _15646_ ( .A1(_09044_ ), .A2(_08884_ ), .A3(_09135_ ), .ZN(_09136_ ) );
OR3_X1 _15647_ ( .A1(_09134_ ), .A2(_09043_ ), .A3(_09136_ ), .ZN(_09137_ ) );
OR2_X1 _15648_ ( .A1(_09130_ ), .A2(_09137_ ), .ZN(_09138_ ) );
AND2_X1 _15649_ ( .A1(\exu.add.io_rs1_data [23] ), .A2(\exu.addi.io_imm [23] ), .ZN(_09139_ ) );
NOR2_X1 _15650_ ( .A1(\exu.add.io_rs1_data [23] ), .A2(\exu.addi.io_imm [23] ), .ZN(_09140_ ) );
NOR2_X1 _15651_ ( .A1(_09139_ ), .A2(_09140_ ), .ZN(_09141_ ) );
AND2_X1 _15652_ ( .A1(\exu.add.io_rs1_data [22] ), .A2(\exu.addi.io_imm [22] ), .ZN(_09142_ ) );
NOR2_X1 _15653_ ( .A1(\exu.add.io_rs1_data [22] ), .A2(\exu.addi.io_imm [22] ), .ZN(_09143_ ) );
NOR2_X1 _15654_ ( .A1(_09142_ ), .A2(_09143_ ), .ZN(_09144_ ) );
AND2_X1 _15655_ ( .A1(\exu.add.io_rs1_data [21] ), .A2(\exu.addi.io_imm [21] ), .ZN(_09145_ ) );
NOR2_X1 _15656_ ( .A1(\exu.add.io_rs1_data [21] ), .A2(\exu.addi.io_imm [21] ), .ZN(_09146_ ) );
NOR2_X1 _15657_ ( .A1(_09145_ ), .A2(_09146_ ), .ZN(_09147_ ) );
AND2_X1 _15658_ ( .A1(\exu.add.io_rs1_data [20] ), .A2(\exu.addi.io_imm [20] ), .ZN(_09148_ ) );
NOR2_X1 _15659_ ( .A1(\exu.add.io_rs1_data [20] ), .A2(\exu.addi.io_imm [20] ), .ZN(_09149_ ) );
NOR2_X1 _15660_ ( .A1(_09148_ ), .A2(_09149_ ), .ZN(_09150_ ) );
AND2_X1 _15661_ ( .A1(_09147_ ), .A2(_09150_ ), .ZN(_09151_ ) );
NAND4_X1 _15662_ ( .A1(_09138_ ), .A2(_09141_ ), .A3(_09144_ ), .A4(_09151_ ), .ZN(_09152_ ) );
AOI21_X1 _15663_ ( .A(_09145_ ), .B1(_09147_ ), .B2(_09148_ ), .ZN(_09153_ ) );
INV_X1 _15664_ ( .A(_09141_ ), .ZN(_09154_ ) );
INV_X1 _15665_ ( .A(_09144_ ), .ZN(_09155_ ) );
NOR3_X1 _15666_ ( .A1(_09153_ ), .A2(_09154_ ), .A3(_09155_ ), .ZN(_09156_ ) );
INV_X1 _15667_ ( .A(\exu.addi.io_imm [22] ), .ZN(_09157_ ) );
NOR4_X1 _15668_ ( .A1(_09139_ ), .A2(_09140_ ), .A3(_08887_ ), .A4(_09157_ ), .ZN(_09158_ ) );
NOR3_X1 _15669_ ( .A1(_09156_ ), .A2(_09139_ ), .A3(_09158_ ), .ZN(_09159_ ) );
NAND2_X1 _15670_ ( .A1(_09152_ ), .A2(_09159_ ), .ZN(_09160_ ) );
AND2_X1 _15671_ ( .A1(\exu.add.io_rs1_data [24] ), .A2(\exu.addi.io_imm [24] ), .ZN(_09161_ ) );
NOR2_X1 _15672_ ( .A1(\exu.add.io_rs1_data [24] ), .A2(\exu.addi.io_imm [24] ), .ZN(_09162_ ) );
NOR2_X1 _15673_ ( .A1(_09161_ ), .A2(_09162_ ), .ZN(_09163_ ) );
AND2_X1 _15674_ ( .A1(\exu.add.io_rs1_data [25] ), .A2(\exu.addi.io_imm [25] ), .ZN(_09164_ ) );
NOR2_X1 _15675_ ( .A1(\exu.add.io_rs1_data [25] ), .A2(\exu.addi.io_imm [25] ), .ZN(_09165_ ) );
NOR2_X1 _15676_ ( .A1(_09164_ ), .A2(_09165_ ), .ZN(_09166_ ) );
AND3_X1 _15677_ ( .A1(_09160_ ), .A2(_09163_ ), .A3(_09166_ ), .ZN(_09167_ ) );
AND2_X1 _15678_ ( .A1(_09166_ ), .A2(_09161_ ), .ZN(_09168_ ) );
NOR3_X1 _15679_ ( .A1(_09167_ ), .A2(_09164_ ), .A3(_09168_ ), .ZN(_09169_ ) );
AND2_X1 _15680_ ( .A1(\exu.add.io_rs1_data [26] ), .A2(\exu.addi.io_imm [26] ), .ZN(_09170_ ) );
NOR2_X1 _15681_ ( .A1(\exu.add.io_rs1_data [26] ), .A2(\exu.addi.io_imm [26] ), .ZN(_09171_ ) );
NOR2_X1 _15682_ ( .A1(_09170_ ), .A2(_09171_ ), .ZN(_09172_ ) );
XNOR2_X1 _15683_ ( .A(_09169_ ), .B(_09172_ ), .ZN(\exu.addi._io_rd_T_4 [26] ) );
NOR2_X1 _15684_ ( .A1(_09041_ ), .A2(fanout_net_17 ), .ZN(_09173_ ) );
BUF_X2 _15685_ ( .A(_09173_ ), .Z(_09174_ ) );
AND2_X1 _15686_ ( .A1(\exu.addi._io_rd_T_4 [26] ), .A2(_09174_ ), .ZN(_09175_ ) );
INV_X1 _15687_ ( .A(_09173_ ), .ZN(_09176_ ) );
BUF_X2 _15688_ ( .A(_09176_ ), .Z(_09177_ ) );
AOI211_X1 _15689_ ( .A(_09042_ ), .B(_09175_ ), .C1(_08703_ ), .C2(_09177_ ), .ZN(_09178_ ) );
OR3_X1 _15690_ ( .A1(_08992_ ), .A2(_09040_ ), .A3(_09178_ ), .ZN(_09179_ ) );
NOR2_X1 _15691_ ( .A1(fanout_net_14 ), .A2(fanout_net_15 ), .ZN(_09180_ ) );
BUF_X4 _15692_ ( .A(_09180_ ), .Z(_09181_ ) );
BUF_X4 _15693_ ( .A(_09181_ ), .Z(_09182_ ) );
BUF_X4 _15694_ ( .A(_09182_ ), .Z(_09183_ ) );
BUF_X2 _15695_ ( .A(_09038_ ), .Z(_09184_ ) );
BUF_X2 _15696_ ( .A(_09184_ ), .Z(_09185_ ) );
OR2_X1 _15697_ ( .A1(_09185_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_1_A_$_MUX__Y_B ), .ZN(_09186_ ) );
NAND3_X1 _15698_ ( .A1(_09179_ ), .A2(_09183_ ), .A3(_09186_ ), .ZN(_09187_ ) );
OAI21_X1 _15699_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_1_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09188_ ) );
AND2_X2 _15700_ ( .A1(_09187_ ), .A2(_09188_ ), .ZN(_09189_ ) );
BUF_X4 _15701_ ( .A(_08978_ ), .Z(_09190_ ) );
BUF_X4 _15702_ ( .A(_09190_ ), .Z(_09191_ ) );
BUF_X4 _15703_ ( .A(_09191_ ), .Z(_09192_ ) );
NAND3_X1 _15704_ ( .A1(_09192_ ), .A2(fanout_net_8 ), .A3(\exu.csrrs.io_csr_rdata [4] ), .ZN(_09193_ ) );
INV_X1 _15705_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_27_A_$_MUX__A_B ), .ZN(_09194_ ) );
NAND2_X1 _15706_ ( .A1(_08791_ ), .A2(_09194_ ), .ZN(_09195_ ) );
INV_X1 _15707_ ( .A(\exu.auipc.io_rs1_data [3] ), .ZN(_09196_ ) );
INV_X1 _15708_ ( .A(\exu.auipc.io_rs1_data [2] ), .ZN(_09197_ ) );
OAI21_X1 _15709_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_27_A_$_MUX__A_B ), .B1(_09196_ ), .B2(_09197_ ), .ZN(_09198_ ) );
AND2_X1 _15710_ ( .A1(_09195_ ), .A2(_09198_ ), .ZN(_09199_ ) );
INV_X1 _15711_ ( .A(_09199_ ), .ZN(_09200_ ) );
OAI211_X1 _15712_ ( .A(\exu.bne.io_is ), .B(_09200_ ), .C1(_08781_ ), .C2(fanout_net_17 ), .ZN(_09201_ ) );
INV_X2 _15713_ ( .A(_08815_ ), .ZN(_09202_ ) );
XOR2_X1 _15714_ ( .A(_08598_ ), .B(_08585_ ), .Z(_09203_ ) );
AND3_X1 _15715_ ( .A1(_08921_ ), .A2(_08923_ ), .A3(_09203_ ), .ZN(_09204_ ) );
AOI211_X1 _15716_ ( .A(_08922_ ), .B(_09204_ ), .C1(_08926_ ), .C2(_09199_ ), .ZN(_09205_ ) );
AND4_X1 _15717_ ( .A1(_08866_ ), .A2(_08917_ ), .A3(_08941_ ), .A4(_09203_ ), .ZN(_09206_ ) );
INV_X1 _15718_ ( .A(_08943_ ), .ZN(_09207_ ) );
AOI211_X1 _15719_ ( .A(_08940_ ), .B(_09206_ ), .C1(_09207_ ), .C2(_09199_ ), .ZN(_09208_ ) );
NOR2_X1 _15720_ ( .A1(_09035_ ), .A2(fanout_net_11 ), .ZN(_09209_ ) );
INV_X1 _15721_ ( .A(_09209_ ), .ZN(_09210_ ) );
BUF_X4 _15722_ ( .A(_08949_ ), .Z(_09211_ ) );
AND2_X1 _15723_ ( .A1(fanout_net_17 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_27_A_$_MUX__A_B ), .ZN(_09212_ ) );
OAI22_X1 _15724_ ( .A1(_09200_ ), .A2(_09210_ ), .B1(_09211_ ), .B2(_09212_ ), .ZN(_09213_ ) );
INV_X1 _15725_ ( .A(_08971_ ), .ZN(_09214_ ) );
AND3_X1 _15726_ ( .A1(\exu.csrrs.io_csr_rdata [3] ), .A2(\exu.csrrs.io_csr_rdata [2] ), .A3(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ), .ZN(_09215_ ) );
AOI21_X1 _15727_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ), .B1(\exu.csrrs.io_csr_rdata [3] ), .B2(\exu.csrrs.io_csr_rdata [2] ), .ZN(_09216_ ) );
OR3_X1 _15728_ ( .A1(_09214_ ), .A2(_09215_ ), .A3(_09216_ ), .ZN(_09217_ ) );
AOI21_X1 _15729_ ( .A(fanout_net_7 ), .B1(_09213_ ), .B2(_09217_ ), .ZN(_09218_ ) );
OAI21_X1 _15730_ ( .A(_08947_ ), .B1(_09208_ ), .B2(_09218_ ), .ZN(_09219_ ) );
BUF_X4 _15731_ ( .A(_08976_ ), .Z(_09220_ ) );
MUX2_X1 _15732_ ( .A(_09199_ ), .B(_09203_ ), .S(_09220_ ), .Z(_09221_ ) );
BUF_X4 _15733_ ( .A(_08947_ ), .Z(_09222_ ) );
OAI211_X1 _15734_ ( .A(_08931_ ), .B(_09219_ ), .C1(_09221_ ), .C2(_09222_ ), .ZN(_09223_ ) );
MUX2_X1 _15735_ ( .A(_09199_ ), .B(_09203_ ), .S(_08935_ ), .Z(_09224_ ) );
AOI21_X1 _15736_ ( .A(\exu.bge.io_is ), .B1(_09224_ ), .B2(\exu.bgeu.io_is ), .ZN(_09225_ ) );
AOI21_X1 _15737_ ( .A(_09205_ ), .B1(_09223_ ), .B2(_09225_ ), .ZN(_09226_ ) );
OAI221_X1 _15738_ ( .A(_09201_ ), .B1(_09202_ ), .B2(_09203_ ), .C1(_09226_ ), .C2(\exu.bne.io_is ), .ZN(_09227_ ) );
NAND2_X1 _15739_ ( .A1(_09227_ ), .A2(_08788_ ), .ZN(_09228_ ) );
NOR3_X1 _15740_ ( .A1(_08777_ ), .A2(_08782_ ), .A3(_08780_ ), .ZN(_09229_ ) );
NAND3_X1 _15741_ ( .A1(_09203_ ), .A2(_09191_ ), .A3(_09229_ ), .ZN(_09230_ ) );
AND2_X2 _15742_ ( .A1(_09229_ ), .A2(_09190_ ), .ZN(_09231_ ) );
OAI211_X1 _15743_ ( .A(_09230_ ), .B(\exu.beq.io_is ), .C1(_09231_ ), .C2(_09200_ ), .ZN(_09232_ ) );
AOI21_X1 _15744_ ( .A(fanout_net_9 ), .B1(_09228_ ), .B2(_09232_ ), .ZN(_09233_ ) );
MUX2_X1 _15745_ ( .A(_09194_ ), .B(_09203_ ), .S(_08699_ ), .Z(_09234_ ) );
OAI21_X1 _15746_ ( .A(_08989_ ), .B1(_09234_ ), .B2(_08698_ ), .ZN(_09235_ ) );
OAI211_X1 _15747_ ( .A(_09042_ ), .B(_09193_ ), .C1(_09233_ ), .C2(_09235_ ), .ZN(_09236_ ) );
NAND2_X1 _15748_ ( .A1(_09064_ ), .A2(_09066_ ), .ZN(_09237_ ) );
XNOR2_X1 _15749_ ( .A(_09237_ ), .B(_09050_ ), .ZN(\exu.addi._io_rd_T_4 [4] ) );
NAND2_X1 _15750_ ( .A1(\exu.addi._io_rd_T_4 [4] ), .A2(_09174_ ), .ZN(_09238_ ) );
OAI211_X1 _15751_ ( .A(_09238_ ), .B(fanout_net_10 ), .C1(_09192_ ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_27_A_$_MUX__A_B ), .ZN(_09239_ ) );
NAND3_X1 _15752_ ( .A1(_09236_ ), .A2(_09038_ ), .A3(_09239_ ), .ZN(_09240_ ) );
INV_X1 _15753_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__Y_B ), .ZN(_09241_ ) );
OAI21_X1 _15754_ ( .A(_09241_ ), .B1(_09037_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_09242_ ) );
NAND2_X1 _15755_ ( .A1(_09240_ ), .A2(_09242_ ), .ZN(\ifu.io_out_bits_pc [4] ) );
NAND2_X1 _15756_ ( .A1(\ifu.io_out_bits_pc [4] ), .A2(_09180_ ), .ZN(_09243_ ) );
OAI21_X1 _15757_ ( .A(_09241_ ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09244_ ) );
NAND2_X2 _15758_ ( .A1(_09243_ ), .A2(_09244_ ), .ZN(_09245_ ) );
BUF_X4 _15759_ ( .A(_09245_ ), .Z(_09246_ ) );
MUX2_X1 _15760_ ( .A(\icache.tag_reg_0 [21] ), .B(\icache.tag_reg_1 [21] ), .S(_09246_ ), .Z(_09247_ ) );
XOR2_X1 _15761_ ( .A(_09189_ ), .B(_09247_ ), .Z(_09248_ ) );
BUF_X4 _15762_ ( .A(_08788_ ), .Z(_09249_ ) );
BUF_X4 _15763_ ( .A(_08922_ ), .Z(_09250_ ) );
BUF_X4 _15764_ ( .A(_09250_ ), .Z(_09251_ ) );
BUF_X4 _15765_ ( .A(_09222_ ), .Z(_09252_ ) );
BUF_X4 _15766_ ( .A(_09252_ ), .Z(_09253_ ) );
BUF_X4 _15767_ ( .A(_08940_ ), .Z(_09254_ ) );
BUF_X4 _15768_ ( .A(_09254_ ), .Z(_09255_ ) );
BUF_X4 _15769_ ( .A(_09255_ ), .Z(_09256_ ) );
BUF_X2 _15770_ ( .A(_09207_ ), .Z(_09257_ ) );
AND2_X1 _15771_ ( .A1(_08685_ ), .A2(_08686_ ), .ZN(_09258_ ) );
INV_X1 _15772_ ( .A(_08689_ ), .ZN(_09259_ ) );
OR3_X1 _15773_ ( .A1(_09258_ ), .A2(_08691_ ), .A3(_09259_ ), .ZN(_09260_ ) );
OAI21_X1 _15774_ ( .A(_09259_ ), .B1(_09258_ ), .B2(_08691_ ), .ZN(_09261_ ) );
AOI21_X1 _15775_ ( .A(_09257_ ), .B1(_09260_ ), .B2(_09261_ ), .ZN(_09262_ ) );
AND3_X1 _15776_ ( .A1(_08806_ ), .A2(\exu.auipc.io_rs1_data [21] ), .A3(\exu.auipc.io_rs1_data [20] ), .ZN(_09263_ ) );
AND3_X1 _15777_ ( .A1(_08798_ ), .A2(_09263_ ), .A3(_08803_ ), .ZN(_09264_ ) );
NAND3_X1 _15778_ ( .A1(_09264_ ), .A2(\exu.auipc.io_rs1_data [22] ), .A3(\exu.auipc.io_rs1_data [23] ), .ZN(_09265_ ) );
NOR2_X1 _15779_ ( .A1(_09265_ ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_7_A_$_MUX__A_B ), .ZN(_09266_ ) );
INV_X1 _15780_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_6_A_$_MUX__A_B ), .ZN(_09267_ ) );
XNOR2_X1 _15781_ ( .A(_09266_ ), .B(_09267_ ), .ZN(_09268_ ) );
INV_X1 _15782_ ( .A(_09268_ ), .ZN(_09269_ ) );
AOI211_X1 _15783_ ( .A(_09256_ ), .B(_09262_ ), .C1(_09257_ ), .C2(_09269_ ), .ZN(_09270_ ) );
BUF_X4 _15784_ ( .A(_09214_ ), .Z(_09271_ ) );
NOR3_X1 _15785_ ( .A1(_08955_ ), .A2(_08961_ ), .A3(_08956_ ), .ZN(_09272_ ) );
AND3_X1 _15786_ ( .A1(_09272_ ), .A2(\exu.csrrs.io_csr_rdata [11] ), .A3(\exu.csrrs.io_csr_rdata [12] ), .ZN(_09273_ ) );
AND2_X1 _15787_ ( .A1(_09273_ ), .A2(\exu.csrrs.io_csr_rdata [13] ), .ZN(_09274_ ) );
AND2_X1 _15788_ ( .A1(_09274_ ), .A2(\exu.csrrs.io_csr_rdata [14] ), .ZN(_09275_ ) );
AND2_X1 _15789_ ( .A1(_09275_ ), .A2(\exu.csrrs.io_csr_rdata [15] ), .ZN(_09276_ ) );
AND2_X1 _15790_ ( .A1(_09276_ ), .A2(\exu.csrrs.io_csr_rdata [16] ), .ZN(_09277_ ) );
AND2_X1 _15791_ ( .A1(_09277_ ), .A2(\exu.csrrs.io_csr_rdata [17] ), .ZN(_09278_ ) );
AND2_X1 _15792_ ( .A1(_09278_ ), .A2(\exu.csrrs.io_csr_rdata [18] ), .ZN(_09279_ ) );
AND3_X1 _15793_ ( .A1(_09279_ ), .A2(\exu.csrrs.io_csr_rdata [20] ), .A3(\exu.csrrs.io_csr_rdata [19] ), .ZN(_09280_ ) );
AND2_X1 _15794_ ( .A1(_09280_ ), .A2(\exu.csrrs.io_csr_rdata [21] ), .ZN(_09281_ ) );
AND2_X1 _15795_ ( .A1(_09281_ ), .A2(\exu.csrrs.io_csr_rdata [22] ), .ZN(_09282_ ) );
AND2_X1 _15796_ ( .A1(_09282_ ), .A2(\exu.csrrs.io_csr_rdata [23] ), .ZN(_09283_ ) );
AOI21_X1 _15797_ ( .A(_09271_ ), .B1(_09283_ ), .B2(_08966_ ), .ZN(_09284_ ) );
AND4_X1 _15798_ ( .A1(\exu.csrrs.io_csr_rdata [24] ), .A2(_08963_ ), .A3(_08967_ ), .A4(_08965_ ), .ZN(_09285_ ) );
OAI21_X1 _15799_ ( .A(_09284_ ), .B1(\exu.csrrs.io_csr_rdata [25] ), .B2(_09285_ ), .ZN(_09286_ ) );
OAI211_X1 _15800_ ( .A(_09286_ ), .B(fanout_net_11 ), .C1(_09191_ ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_6_A_$_MUX__A_B ), .ZN(_09287_ ) );
BUF_X2 _15801_ ( .A(_09211_ ), .Z(_09288_ ) );
OAI21_X1 _15802_ ( .A(_09288_ ), .B1(_09268_ ), .B2(_09036_ ), .ZN(_09289_ ) );
AOI21_X1 _15803_ ( .A(fanout_net_7 ), .B1(_09287_ ), .B2(_09289_ ), .ZN(_09290_ ) );
OAI21_X1 _15804_ ( .A(_09253_ ), .B1(_09270_ ), .B2(_09290_ ), .ZN(_09291_ ) );
NAND2_X1 _15805_ ( .A1(_09260_ ), .A2(_09261_ ), .ZN(_09292_ ) );
BUF_X4 _15806_ ( .A(_09220_ ), .Z(_09293_ ) );
NAND2_X1 _15807_ ( .A1(_09292_ ), .A2(_09293_ ), .ZN(_09294_ ) );
OAI211_X1 _15808_ ( .A(_09294_ ), .B(fanout_net_6 ), .C1(_09293_ ), .C2(_09268_ ), .ZN(_09295_ ) );
AOI21_X1 _15809_ ( .A(\exu.bgeu.io_is ), .B1(_09291_ ), .B2(_09295_ ), .ZN(_09296_ ) );
BUF_X2 _15810_ ( .A(_08936_ ), .Z(_09297_ ) );
BUF_X2 _15811_ ( .A(_08938_ ), .Z(_09298_ ) );
INV_X1 _15812_ ( .A(_09298_ ), .ZN(_09299_ ) );
OAI22_X1 _15813_ ( .A1(_09292_ ), .A2(_09297_ ), .B1(_09299_ ), .B2(_09269_ ), .ZN(_09300_ ) );
OAI21_X1 _15814_ ( .A(_09251_ ), .B1(_09296_ ), .B2(_09300_ ), .ZN(_09301_ ) );
INV_X1 _15815_ ( .A(_09292_ ), .ZN(_09302_ ) );
BUF_X4 _15816_ ( .A(_08925_ ), .Z(_09303_ ) );
AOI22_X1 _15817_ ( .A1(_09302_ ), .A2(_09303_ ), .B1(_08928_ ), .B2(_09268_ ), .ZN(_09304_ ) );
AOI21_X1 _15818_ ( .A(\exu.bne.io_is ), .B1(_09301_ ), .B2(_09304_ ), .ZN(_09305_ ) );
BUF_X4 _15819_ ( .A(_09202_ ), .Z(_09306_ ) );
NOR2_X1 _15820_ ( .A1(_08815_ ), .A2(_08812_ ), .ZN(_09307_ ) );
INV_X1 _15821_ ( .A(_09307_ ), .ZN(_09308_ ) );
BUF_X4 _15822_ ( .A(_09308_ ), .Z(_09309_ ) );
OAI22_X1 _15823_ ( .A1(_09292_ ), .A2(_09306_ ), .B1(_09309_ ), .B2(_09269_ ), .ZN(_09310_ ) );
OAI21_X1 _15824_ ( .A(_09249_ ), .B1(_09305_ ), .B2(_09310_ ), .ZN(_09311_ ) );
BUF_X4 _15825_ ( .A(_08784_ ), .Z(_09312_ ) );
BUF_X4 _15826_ ( .A(_08789_ ), .Z(_09313_ ) );
AOI22_X1 _15827_ ( .A1(_09302_ ), .A2(_09312_ ), .B1(_09313_ ), .B2(_09268_ ), .ZN(_09314_ ) );
AOI21_X1 _15828_ ( .A(fanout_net_9 ), .B1(_09311_ ), .B2(_09314_ ), .ZN(_09315_ ) );
AND2_X1 _15829_ ( .A1(fanout_net_9 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_6_A_$_MUX__A_B ), .ZN(_09316_ ) );
BUF_X4 _15830_ ( .A(_08700_ ), .Z(_09317_ ) );
MUX2_X1 _15831_ ( .A(_09316_ ), .B(_09302_ ), .S(_09317_ ), .Z(_09318_ ) );
NOR3_X1 _15832_ ( .A1(_09315_ ), .A2(fanout_net_8 ), .A3(_09318_ ), .ZN(_09319_ ) );
AOI211_X1 _15833_ ( .A(fanout_net_10 ), .B(_09319_ ), .C1(\exu.csrrs.io_csr_rdata [25] ), .C2(_08991_ ), .ZN(_09320_ ) );
BUF_X4 _15834_ ( .A(_09042_ ), .Z(_09321_ ) );
INV_X1 _15835_ ( .A(_09163_ ), .ZN(_09322_ ) );
AOI21_X1 _15836_ ( .A(_09322_ ), .B1(_09152_ ), .B2(_09159_ ), .ZN(_09323_ ) );
NOR2_X1 _15837_ ( .A1(_09323_ ), .A2(_09161_ ), .ZN(_09324_ ) );
XNOR2_X1 _15838_ ( .A(_09324_ ), .B(_09166_ ), .ZN(\exu.addi._io_rd_T_4 [25] ) );
AND2_X1 _15839_ ( .A1(\exu.addi._io_rd_T_4 [25] ), .A2(_09174_ ), .ZN(_09325_ ) );
AOI211_X1 _15840_ ( .A(_09321_ ), .B(_09325_ ), .C1(fanout_net_17 ), .C2(_09267_ ), .ZN(_09326_ ) );
OR3_X1 _15841_ ( .A1(_09320_ ), .A2(_09040_ ), .A3(_09326_ ), .ZN(_09327_ ) );
BUF_X4 _15842_ ( .A(_09185_ ), .Z(_09328_ ) );
OR2_X1 _15843_ ( .A1(_09328_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_2_A_$_MUX__Y_B ), .ZN(_09329_ ) );
NAND3_X1 _15844_ ( .A1(_09327_ ), .A2(_09183_ ), .A3(_09329_ ), .ZN(_09330_ ) );
OAI21_X1 _15845_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_2_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09331_ ) );
BUF_X4 _15846_ ( .A(_09246_ ), .Z(_09332_ ) );
NAND2_X1 _15847_ ( .A1(_09332_ ), .A2(\icache.tag_reg_1 [20] ), .ZN(_09333_ ) );
BUF_X4 _15848_ ( .A(_09243_ ), .Z(_09334_ ) );
BUF_X2 _15849_ ( .A(_09334_ ), .Z(_09335_ ) );
BUF_X4 _15850_ ( .A(_09244_ ), .Z(_09336_ ) );
BUF_X2 _15851_ ( .A(_09336_ ), .Z(_09337_ ) );
NAND3_X1 _15852_ ( .A1(_09335_ ), .A2(\icache.tag_reg_0 [20] ), .A3(_09337_ ), .ZN(_09338_ ) );
AND4_X1 _15853_ ( .A1(_09330_ ), .A2(_09331_ ), .A3(_09333_ ), .A4(_09338_ ), .ZN(_09339_ ) );
AOI22_X1 _15854_ ( .A1(_09330_ ), .A2(_09331_ ), .B1(_09333_ ), .B2(_09338_ ), .ZN(_09340_ ) );
OR3_X1 _15855_ ( .A1(_09248_ ), .A2(_09339_ ), .A3(_09340_ ), .ZN(_09341_ ) );
INV_X1 _15856_ ( .A(\ifu.io_out_bits_pc_$_MUX__Y_9_A_$_MUX__Y_A_$_OR__Y_B_$_ANDNOT__Y_A ), .ZN(_09342_ ) );
AND2_X2 _15857_ ( .A1(_08990_ ), .A2(_09342_ ), .ZN(_09343_ ) );
XOR2_X1 _15858_ ( .A(\exu.addi.io_imm [27] ), .B(\exu.auipc.io_rs1_data [27] ), .Z(_09344_ ) );
INV_X1 _15859_ ( .A(_09344_ ), .ZN(_09345_ ) );
NOR2_X1 _15860_ ( .A1(_09345_ ), .A2(_08696_ ), .ZN(_09346_ ) );
NAND4_X1 _15861_ ( .A1(_08685_ ), .A2(_09346_ ), .A3(_08686_ ), .A4(_08689_ ), .ZN(_09347_ ) );
AND2_X1 _15862_ ( .A1(\exu.addi.io_imm [26] ), .A2(\exu.auipc.io_rs1_data [26] ), .ZN(_09348_ ) );
AND2_X1 _15863_ ( .A1(_09344_ ), .A2(_09348_ ), .ZN(_09349_ ) );
AOI221_X4 _15864_ ( .A(_09349_ ), .B1(\exu.addi.io_imm [27] ), .B2(\exu.auipc.io_rs1_data [27] ), .C1(_09346_ ), .C2(_08694_ ), .ZN(_09350_ ) );
AND2_X1 _15865_ ( .A1(_09347_ ), .A2(_09350_ ), .ZN(_09351_ ) );
XNOR2_X1 _15866_ ( .A(\exu.addi.io_imm [28] ), .B(\exu.auipc.io_rs1_data [28] ), .ZN(_09352_ ) );
XOR2_X1 _15867_ ( .A(_09351_ ), .B(_09352_ ), .Z(_09353_ ) );
BUF_X2 _15868_ ( .A(_08945_ ), .Z(_09354_ ) );
AND2_X1 _15869_ ( .A1(_09353_ ), .A2(_09354_ ), .ZN(_09355_ ) );
AND3_X1 _15870_ ( .A1(_08808_ ), .A2(\exu.auipc.io_rs1_data [27] ), .A3(\exu.auipc.io_rs1_data [26] ), .ZN(_09356_ ) );
XNOR2_X1 _15871_ ( .A(_09356_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_3_A_$_MUX__A_B ), .ZN(_09357_ ) );
AOI211_X1 _15872_ ( .A(_09256_ ), .B(_09355_ ), .C1(_09257_ ), .C2(_09357_ ), .ZN(_09358_ ) );
NAND3_X1 _15873_ ( .A1(fanout_net_17 ), .A2(fanout_net_11 ), .A3(\exu.addi._io_rd_T_4_$_NOT__Y_3_A_$_MUX__A_B ), .ZN(_09359_ ) );
AND3_X1 _15874_ ( .A1(_08969_ ), .A2(\exu.csrrs.io_csr_rdata [27] ), .A3(\exu.csrrs.io_csr_rdata [26] ), .ZN(_09360_ ) );
XOR2_X1 _15875_ ( .A(_09360_ ), .B(\exu.csrrs.io_csr_rdata [28] ), .Z(_09361_ ) );
AND2_X1 _15876_ ( .A1(_09357_ ), .A2(exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ), .ZN(_09362_ ) );
OAI221_X1 _15877_ ( .A(_09359_ ), .B1(_09271_ ), .B2(_09361_ ), .C1(_09362_ ), .C2(fanout_net_11 ), .ZN(_09363_ ) );
AND2_X1 _15878_ ( .A1(_09363_ ), .A2(_09256_ ), .ZN(_09364_ ) );
OAI21_X1 _15879_ ( .A(_09253_ ), .B1(_09358_ ), .B2(_09364_ ), .ZN(_09365_ ) );
NAND2_X1 _15880_ ( .A1(_09353_ ), .A2(_09293_ ), .ZN(_09366_ ) );
INV_X1 _15881_ ( .A(_09357_ ), .ZN(_09367_ ) );
OAI211_X1 _15882_ ( .A(_09366_ ), .B(fanout_net_6 ), .C1(_09293_ ), .C2(_09367_ ), .ZN(_09368_ ) );
AOI21_X1 _15883_ ( .A(\exu.bgeu.io_is ), .B1(_09365_ ), .B2(_09368_ ), .ZN(_09369_ ) );
OAI22_X1 _15884_ ( .A1(_09353_ ), .A2(_09297_ ), .B1(_09299_ ), .B2(_09357_ ), .ZN(_09370_ ) );
OAI21_X1 _15885_ ( .A(_09251_ ), .B1(_09369_ ), .B2(_09370_ ), .ZN(_09371_ ) );
INV_X1 _15886_ ( .A(_09353_ ), .ZN(_09372_ ) );
AOI22_X1 _15887_ ( .A1(_09372_ ), .A2(_09303_ ), .B1(_08928_ ), .B2(_09367_ ), .ZN(_09373_ ) );
AOI21_X1 _15888_ ( .A(\exu.bne.io_is ), .B1(_09371_ ), .B2(_09373_ ), .ZN(_09374_ ) );
OAI22_X1 _15889_ ( .A1(_09353_ ), .A2(_09306_ ), .B1(_09309_ ), .B2(_09357_ ), .ZN(_09375_ ) );
OAI21_X1 _15890_ ( .A(_09249_ ), .B1(_09374_ ), .B2(_09375_ ), .ZN(_09376_ ) );
AOI22_X1 _15891_ ( .A1(_09372_ ), .A2(_09312_ ), .B1(_09313_ ), .B2(_09367_ ), .ZN(_09377_ ) );
AOI21_X1 _15892_ ( .A(fanout_net_9 ), .B1(_09376_ ), .B2(_09377_ ), .ZN(_09378_ ) );
MUX2_X1 _15893_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_3_A_$_MUX__A_B ), .B(_09372_ ), .S(_09317_ ), .Z(_09379_ ) );
AOI21_X1 _15894_ ( .A(_09378_ ), .B1(fanout_net_9 ), .B2(_09379_ ), .ZN(_09380_ ) );
AOI221_X4 _15895_ ( .A(fanout_net_10 ), .B1(\exu.csrrs.io_csr_rdata [28] ), .B2(_09343_ ), .C1(_09380_ ), .C2(\ifu.io_out_bits_pc_$_MUX__Y_9_A_$_MUX__Y_A_$_OR__Y_B_$_ANDNOT__Y_A ), .ZN(_09381_ ) );
INV_X1 _15896_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_3_A_$_MUX__A_B ), .ZN(_09382_ ) );
AND2_X1 _15897_ ( .A1(\exu.add.io_rs1_data [27] ), .A2(\exu.addi.io_imm [27] ), .ZN(_09383_ ) );
NOR2_X1 _15898_ ( .A1(\exu.add.io_rs1_data [27] ), .A2(\exu.addi.io_imm [27] ), .ZN(_09384_ ) );
INV_X1 _15899_ ( .A(_09172_ ), .ZN(_09385_ ) );
OR4_X1 _15900_ ( .A1(_09383_ ), .A2(_09169_ ), .A3(_09384_ ), .A4(_09385_ ), .ZN(_09386_ ) );
NOR2_X1 _15901_ ( .A1(_09383_ ), .A2(_09384_ ), .ZN(_09387_ ) );
AOI21_X1 _15902_ ( .A(_09383_ ), .B1(_09387_ ), .B2(_09170_ ), .ZN(_09388_ ) );
AND2_X1 _15903_ ( .A1(\exu.add.io_rs1_data [28] ), .A2(\exu.addi.io_imm [28] ), .ZN(_09389_ ) );
NOR2_X1 _15904_ ( .A1(\exu.add.io_rs1_data [28] ), .A2(\exu.addi.io_imm [28] ), .ZN(_09390_ ) );
NOR2_X1 _15905_ ( .A1(_09389_ ), .A2(_09390_ ), .ZN(_09391_ ) );
INV_X1 _15906_ ( .A(_09391_ ), .ZN(_09392_ ) );
AND3_X1 _15907_ ( .A1(_09386_ ), .A2(_09388_ ), .A3(_09392_ ), .ZN(_09393_ ) );
AOI21_X1 _15908_ ( .A(_09392_ ), .B1(_09386_ ), .B2(_09388_ ), .ZN(_09394_ ) );
NOR2_X1 _15909_ ( .A1(_09393_ ), .A2(_09394_ ), .ZN(\exu.addi._io_rd_T_4 [28] ) );
BUF_X4 _15910_ ( .A(_09192_ ), .Z(_09395_ ) );
BUF_X4 _15911_ ( .A(_09395_ ), .Z(_09396_ ) );
MUX2_X1 _15912_ ( .A(_09382_ ), .B(\exu.addi._io_rd_T_4 [28] ), .S(_09396_ ), .Z(_09397_ ) );
NOR2_X1 _15913_ ( .A1(_09397_ ), .A2(_09321_ ), .ZN(_09398_ ) );
OAI21_X1 _15914_ ( .A(_09328_ ), .B1(_09381_ ), .B2(_09398_ ), .ZN(_09399_ ) );
INV_X1 _15915_ ( .A(\ifu.pc [28] ), .ZN(_09400_ ) );
BUF_X4 _15916_ ( .A(_09037_ ), .Z(_09401_ ) );
BUF_X4 _15917_ ( .A(_09401_ ), .Z(_09402_ ) );
OAI21_X1 _15918_ ( .A(_09400_ ), .B1(_09402_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_09403_ ) );
NAND3_X1 _15919_ ( .A1(_09399_ ), .A2(_09183_ ), .A3(_09403_ ), .ZN(_09404_ ) );
OAI21_X1 _15920_ ( .A(\ifu.pc [28] ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09405_ ) );
AND2_X1 _15921_ ( .A1(_09404_ ), .A2(_09405_ ), .ZN(_09406_ ) );
MUX2_X1 _15922_ ( .A(\icache.tag_reg_0 [23] ), .B(\icache.tag_reg_1 [23] ), .S(_09332_ ), .Z(_09407_ ) );
XNOR2_X1 _15923_ ( .A(_09406_ ), .B(_09407_ ), .ZN(_09408_ ) );
BUF_X4 _15924_ ( .A(_08702_ ), .Z(_09409_ ) );
BUF_X4 _15925_ ( .A(_09409_ ), .Z(_09410_ ) );
BUF_X4 _15926_ ( .A(_08984_ ), .Z(_09411_ ) );
BUF_X4 _15927_ ( .A(_08931_ ), .Z(_09412_ ) );
BUF_X4 _15928_ ( .A(_09412_ ), .Z(_09413_ ) );
BUF_X4 _15929_ ( .A(_08972_ ), .Z(_09414_ ) );
AND2_X1 _15930_ ( .A1(fanout_net_11 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_4_A_$_MUX__A_B ), .ZN(_09415_ ) );
OR2_X1 _15931_ ( .A1(_09414_ ), .A2(_09415_ ), .ZN(_09416_ ) );
INV_X1 _15932_ ( .A(_09360_ ), .ZN(_09417_ ) );
AND4_X1 _15933_ ( .A1(\exu.csrrs.io_csr_rdata [26] ), .A2(_08957_ ), .A3(_08968_ ), .A4(_08962_ ), .ZN(_09418_ ) );
OAI211_X1 _15934_ ( .A(_09417_ ), .B(_09414_ ), .C1(\exu.csrrs.io_csr_rdata [27] ), .C2(_09418_ ), .ZN(_09419_ ) );
XNOR2_X1 _15935_ ( .A(_08810_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_4_A_$_MUX__A_B ), .ZN(_09420_ ) );
OR2_X1 _15936_ ( .A1(_09420_ ), .A2(_09036_ ), .ZN(_09421_ ) );
AOI221_X4 _15937_ ( .A(fanout_net_7 ), .B1(_09416_ ), .B2(_09419_ ), .C1(_09421_ ), .C2(_09288_ ), .ZN(_09422_ ) );
NOR2_X1 _15938_ ( .A1(_08695_ ), .A2(_08696_ ), .ZN(_09423_ ) );
OR3_X1 _15939_ ( .A1(_09423_ ), .A2(_09345_ ), .A3(_09348_ ), .ZN(_09424_ ) );
OAI21_X1 _15940_ ( .A(_09345_ ), .B1(_09423_ ), .B2(_09348_ ), .ZN(_09425_ ) );
NAND2_X1 _15941_ ( .A1(_09424_ ), .A2(_09425_ ), .ZN(_09426_ ) );
INV_X1 _15942_ ( .A(_09426_ ), .ZN(_09427_ ) );
BUF_X2 _15943_ ( .A(_08918_ ), .Z(_09428_ ) );
AND2_X1 _15944_ ( .A1(_09428_ ), .A2(_09190_ ), .ZN(_09429_ ) );
OAI22_X1 _15945_ ( .A1(_09427_ ), .A2(_09257_ ), .B1(_09429_ ), .B2(_09420_ ), .ZN(_09430_ ) );
AOI211_X1 _15946_ ( .A(fanout_net_6 ), .B(_09422_ ), .C1(_09430_ ), .C2(fanout_net_7 ), .ZN(_09431_ ) );
BUF_X4 _15947_ ( .A(_08977_ ), .Z(_09432_ ) );
AOI21_X1 _15948_ ( .A(_09432_ ), .B1(_09424_ ), .B2(_09425_ ), .ZN(_09433_ ) );
INV_X1 _15949_ ( .A(_09420_ ), .ZN(_09434_ ) );
AOI211_X1 _15950_ ( .A(_09253_ ), .B(_09433_ ), .C1(_09432_ ), .C2(_09434_ ), .ZN(_09435_ ) );
OAI21_X1 _15951_ ( .A(_09413_ ), .B1(_09431_ ), .B2(_09435_ ), .ZN(_09436_ ) );
BUF_X4 _15952_ ( .A(_08935_ ), .Z(_09437_ ) );
AOI22_X1 _15953_ ( .A1(_09427_ ), .A2(_09437_ ), .B1(_09298_ ), .B2(_09420_ ), .ZN(_09438_ ) );
AOI21_X1 _15954_ ( .A(\exu.bge.io_is ), .B1(_09436_ ), .B2(_09438_ ), .ZN(_09439_ ) );
BUF_X2 _15955_ ( .A(_08926_ ), .Z(_09440_ ) );
OAI22_X1 _15956_ ( .A1(_09426_ ), .A2(_09440_ ), .B1(_08930_ ), .B2(_09434_ ), .ZN(_09441_ ) );
OAI21_X1 _15957_ ( .A(_09411_ ), .B1(_09439_ ), .B2(_09441_ ), .ZN(_09442_ ) );
BUF_X4 _15958_ ( .A(_08815_ ), .Z(_09443_ ) );
BUF_X4 _15959_ ( .A(_09307_ ), .Z(_09444_ ) );
AOI22_X1 _15960_ ( .A1(_09427_ ), .A2(_09443_ ), .B1(_09444_ ), .B2(_09420_ ), .ZN(_09445_ ) );
AOI21_X1 _15961_ ( .A(\exu.beq.io_is ), .B1(_09442_ ), .B2(_09445_ ), .ZN(_09446_ ) );
NAND3_X1 _15962_ ( .A1(_09424_ ), .A2(_09312_ ), .A3(_09425_ ), .ZN(_09447_ ) );
BUF_X4 _15963_ ( .A(_08790_ ), .Z(_09448_ ) );
OAI21_X1 _15964_ ( .A(_09447_ ), .B1(_09448_ ), .B2(_09434_ ), .ZN(_09449_ ) );
OAI21_X1 _15965_ ( .A(_09410_ ), .B1(_09446_ ), .B2(_09449_ ), .ZN(_09450_ ) );
NAND2_X1 _15966_ ( .A1(fanout_net_9 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_4_A_$_MUX__A_B ), .ZN(_09451_ ) );
BUF_X4 _15967_ ( .A(_09317_ ), .Z(_09452_ ) );
MUX2_X1 _15968_ ( .A(_09451_ ), .B(_09426_ ), .S(_09452_ ), .Z(_09453_ ) );
NAND3_X1 _15969_ ( .A1(_09450_ ), .A2(_08989_ ), .A3(_09453_ ), .ZN(_09454_ ) );
INV_X1 _15970_ ( .A(\exu.csrrs.io_csr_rdata [27] ), .ZN(_09455_ ) );
INV_X1 _15971_ ( .A(_08990_ ), .ZN(_09456_ ) );
OAI211_X1 _15972_ ( .A(_09454_ ), .B(_09321_ ), .C1(_09455_ ), .C2(_09456_ ), .ZN(_09457_ ) );
NOR2_X1 _15973_ ( .A1(_09169_ ), .A2(_09385_ ), .ZN(_09458_ ) );
NOR2_X1 _15974_ ( .A1(_09458_ ), .A2(_09170_ ), .ZN(_09459_ ) );
XNOR2_X1 _15975_ ( .A(_09459_ ), .B(_09387_ ), .ZN(\exu.addi._io_rd_T_4 [27] ) );
BUF_X2 _15976_ ( .A(_09174_ ), .Z(_09460_ ) );
NAND2_X1 _15977_ ( .A1(\exu.addi._io_rd_T_4 [27] ), .A2(_09460_ ), .ZN(_09461_ ) );
BUF_X4 _15978_ ( .A(_09396_ ), .Z(_09462_ ) );
BUF_X4 _15979_ ( .A(_09462_ ), .Z(_09463_ ) );
OAI211_X1 _15980_ ( .A(_09461_ ), .B(fanout_net_10 ), .C1(_09463_ ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_4_A_$_MUX__A_B ), .ZN(_09464_ ) );
NAND3_X1 _15981_ ( .A1(_09457_ ), .A2(_09328_ ), .A3(_09464_ ), .ZN(_09465_ ) );
BUF_X2 _15982_ ( .A(_09183_ ), .Z(_09466_ ) );
OR2_X1 _15983_ ( .A1(_09328_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_09467_ ) );
NAND3_X1 _15984_ ( .A1(_09465_ ), .A2(_09466_ ), .A3(_09467_ ), .ZN(_09468_ ) );
OAI21_X1 _15985_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09469_ ) );
NAND2_X1 _15986_ ( .A1(_09332_ ), .A2(\icache.tag_reg_1 [22] ), .ZN(_09470_ ) );
NAND3_X1 _15987_ ( .A1(_09335_ ), .A2(\icache.tag_reg_0 [22] ), .A3(_09337_ ), .ZN(_09471_ ) );
AOI22_X1 _15988_ ( .A1(_09468_ ), .A2(_09469_ ), .B1(_09470_ ), .B2(_09471_ ), .ZN(_09472_ ) );
AND4_X1 _15989_ ( .A1(_09468_ ), .A2(_09469_ ), .A3(_09470_ ), .A4(_09471_ ), .ZN(_09473_ ) );
NOR4_X1 _15990_ ( .A1(_09341_ ), .A2(_09408_ ), .A3(_09472_ ), .A4(_09473_ ), .ZN(_09474_ ) );
AND2_X1 _15991_ ( .A1(_08654_ ), .A2(_08678_ ), .ZN(_09475_ ) );
INV_X1 _15992_ ( .A(_08658_ ), .ZN(_09476_ ) );
NOR4_X1 _15993_ ( .A1(_09475_ ), .A2(_08659_ ), .A3(_08660_ ), .A4(_09476_ ), .ZN(_09477_ ) );
NOR2_X1 _15994_ ( .A1(_09477_ ), .A2(_08683_ ), .ZN(_09478_ ) );
XNOR2_X1 _15995_ ( .A(\exu.addi.io_imm [22] ), .B(\exu.auipc.io_rs1_data [22] ), .ZN(_09479_ ) );
NOR2_X1 _15996_ ( .A1(_09478_ ), .A2(_09479_ ), .ZN(_09480_ ) );
NOR2_X1 _15997_ ( .A1(_09480_ ), .A2(_08665_ ), .ZN(_09481_ ) );
XNOR2_X1 _15998_ ( .A(_09481_ ), .B(_08655_ ), .ZN(_09482_ ) );
AND2_X1 _15999_ ( .A1(_09482_ ), .A2(_09354_ ), .ZN(_09483_ ) );
NAND2_X1 _16000_ ( .A1(_09264_ ), .A2(\exu.auipc.io_rs1_data [22] ), .ZN(_09484_ ) );
XNOR2_X1 _16001_ ( .A(_09484_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_8_A_$_MUX__A_B ), .ZN(_09485_ ) );
INV_X1 _16002_ ( .A(_09485_ ), .ZN(_09486_ ) );
AOI211_X1 _16003_ ( .A(_09256_ ), .B(_09483_ ), .C1(_09257_ ), .C2(_09486_ ), .ZN(_09487_ ) );
AND2_X1 _16004_ ( .A1(_08963_ ), .A2(_08965_ ), .ZN(_09488_ ) );
NAND2_X1 _16005_ ( .A1(_09488_ ), .A2(_08967_ ), .ZN(_09489_ ) );
AND3_X1 _16006_ ( .A1(_08963_ ), .A2(\exu.csrrs.io_csr_rdata [22] ), .A3(_08965_ ), .ZN(_09490_ ) );
OAI211_X1 _16007_ ( .A(_09489_ ), .B(_09414_ ), .C1(\exu.csrrs.io_csr_rdata [23] ), .C2(_09490_ ), .ZN(_09491_ ) );
OAI211_X1 _16008_ ( .A(_09491_ ), .B(fanout_net_11 ), .C1(_09191_ ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_8_A_$_MUX__A_B ), .ZN(_09492_ ) );
OAI21_X1 _16009_ ( .A(_09288_ ), .B1(_09485_ ), .B2(_09036_ ), .ZN(_09493_ ) );
AOI21_X1 _16010_ ( .A(fanout_net_7 ), .B1(_09492_ ), .B2(_09493_ ), .ZN(_09494_ ) );
OAI21_X1 _16011_ ( .A(_09253_ ), .B1(_09487_ ), .B2(_09494_ ), .ZN(_09495_ ) );
NAND2_X1 _16012_ ( .A1(_09482_ ), .A2(_09293_ ), .ZN(_09496_ ) );
OAI211_X1 _16013_ ( .A(_09496_ ), .B(fanout_net_6 ), .C1(_09293_ ), .C2(_09485_ ), .ZN(_09497_ ) );
AOI21_X1 _16014_ ( .A(\exu.bgeu.io_is ), .B1(_09495_ ), .B2(_09497_ ), .ZN(_09498_ ) );
OAI22_X1 _16015_ ( .A1(_09482_ ), .A2(_09297_ ), .B1(_09299_ ), .B2(_09486_ ), .ZN(_09499_ ) );
OAI21_X1 _16016_ ( .A(_09251_ ), .B1(_09498_ ), .B2(_09499_ ), .ZN(_09500_ ) );
NAND2_X1 _16017_ ( .A1(_09482_ ), .A2(_09303_ ), .ZN(_09501_ ) );
OAI211_X1 _16018_ ( .A(_09501_ ), .B(\exu.bge.io_is ), .C1(_09303_ ), .C2(_09485_ ), .ZN(_09502_ ) );
AOI21_X1 _16019_ ( .A(\exu.bne.io_is ), .B1(_09500_ ), .B2(_09502_ ), .ZN(_09503_ ) );
OAI22_X1 _16020_ ( .A1(_09482_ ), .A2(_09306_ ), .B1(_09309_ ), .B2(_09486_ ), .ZN(_09504_ ) );
OAI21_X1 _16021_ ( .A(_09249_ ), .B1(_09503_ ), .B2(_09504_ ), .ZN(_09505_ ) );
INV_X1 _16022_ ( .A(_09482_ ), .ZN(_09506_ ) );
AOI22_X1 _16023_ ( .A1(_09506_ ), .A2(_09312_ ), .B1(_09313_ ), .B2(_09485_ ), .ZN(_09507_ ) );
AOI21_X1 _16024_ ( .A(fanout_net_9 ), .B1(_09505_ ), .B2(_09507_ ), .ZN(_09508_ ) );
AND2_X1 _16025_ ( .A1(fanout_net_9 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_8_A_$_MUX__A_B ), .ZN(_09509_ ) );
MUX2_X1 _16026_ ( .A(_09509_ ), .B(_09506_ ), .S(_09317_ ), .Z(_09510_ ) );
NOR3_X1 _16027_ ( .A1(_09508_ ), .A2(fanout_net_8 ), .A3(_09510_ ), .ZN(_09511_ ) );
AOI211_X1 _16028_ ( .A(fanout_net_10 ), .B(_09511_ ), .C1(\exu.csrrs.io_csr_rdata [23] ), .C2(_08991_ ), .ZN(_09512_ ) );
OAI21_X1 _16029_ ( .A(_09151_ ), .B1(_09130_ ), .B2(_09137_ ), .ZN(_09513_ ) );
AOI21_X1 _16030_ ( .A(_09155_ ), .B1(_09513_ ), .B2(_09153_ ), .ZN(_09514_ ) );
NOR2_X1 _16031_ ( .A1(_09514_ ), .A2(_09142_ ), .ZN(_09515_ ) );
XNOR2_X1 _16032_ ( .A(_09515_ ), .B(_09141_ ), .ZN(\exu.addi._io_rd_T_4 [23] ) );
NAND2_X1 _16033_ ( .A1(\exu.addi._io_rd_T_4 [23] ), .A2(_09174_ ), .ZN(_09516_ ) );
OAI211_X1 _16034_ ( .A(_09516_ ), .B(fanout_net_10 ), .C1(_09462_ ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_8_A_$_MUX__A_B ), .ZN(_09517_ ) );
INV_X1 _16035_ ( .A(_09517_ ), .ZN(_09518_ ) );
OR3_X1 _16036_ ( .A1(_09512_ ), .A2(_09040_ ), .A3(_09518_ ), .ZN(_09519_ ) );
OR2_X1 _16037_ ( .A1(_09328_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_4_A_$_MUX__Y_B ), .ZN(_09520_ ) );
NAND3_X1 _16038_ ( .A1(_09519_ ), .A2(_09466_ ), .A3(_09520_ ), .ZN(_09521_ ) );
OAI21_X1 _16039_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_4_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09522_ ) );
AND2_X1 _16040_ ( .A1(_09521_ ), .A2(_09522_ ), .ZN(_09523_ ) );
MUX2_X1 _16041_ ( .A(\icache.tag_reg_0 [18] ), .B(\icache.tag_reg_1 [18] ), .S(_09332_ ), .Z(_09524_ ) );
XNOR2_X1 _16042_ ( .A(_09523_ ), .B(_09524_ ), .ZN(_09525_ ) );
XNOR2_X1 _16043_ ( .A(_09478_ ), .B(_08656_ ), .ZN(_09526_ ) );
OR2_X1 _16044_ ( .A1(_09526_ ), .A2(_08786_ ), .ZN(_09527_ ) );
INV_X1 _16045_ ( .A(\exu.auipc.io_rs1_data [22] ), .ZN(_09528_ ) );
XNOR2_X1 _16046_ ( .A(_09264_ ), .B(_09528_ ), .ZN(_09529_ ) );
NOR2_X1 _16047_ ( .A1(_09526_ ), .A2(_09306_ ), .ZN(_09530_ ) );
INV_X1 _16048_ ( .A(_09529_ ), .ZN(_09531_ ) );
OAI211_X1 _16049_ ( .A(\exu.bge.io_is ), .B(_09531_ ), .C1(_08920_ ), .C2(fanout_net_17 ), .ZN(_09532_ ) );
NOR2_X1 _16050_ ( .A1(_09526_ ), .A2(_08936_ ), .ZN(_09533_ ) );
OAI211_X1 _16051_ ( .A(fanout_net_6 ), .B(_09531_ ), .C1(_08921_ ), .C2(fanout_net_17 ), .ZN(_09534_ ) );
INV_X1 _16052_ ( .A(_09429_ ), .ZN(_09535_ ) );
AOI22_X1 _16053_ ( .A1(_09526_ ), .A2(_08945_ ), .B1(_09535_ ), .B2(_09529_ ), .ZN(_09536_ ) );
OAI21_X1 _16054_ ( .A(_09222_ ), .B1(_09536_ ), .B2(_09254_ ), .ZN(_09537_ ) );
NAND2_X1 _16055_ ( .A1(fanout_net_11 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_9_A_$_MUX__A_B ), .ZN(_09538_ ) );
XOR2_X1 _16056_ ( .A(_09488_ ), .B(\exu.csrrs.io_csr_rdata [22] ), .Z(_09539_ ) );
MUX2_X1 _16057_ ( .A(_09538_ ), .B(_09539_ ), .S(_08972_ ), .Z(_09540_ ) );
OAI21_X1 _16058_ ( .A(_09211_ ), .B1(_09531_ ), .B2(_09036_ ), .ZN(_09541_ ) );
AND3_X1 _16059_ ( .A1(_09540_ ), .A2(_09254_ ), .A3(_09541_ ), .ZN(_09542_ ) );
OAI221_X1 _16060_ ( .A(_09534_ ), .B1(_08977_ ), .B2(_09526_ ), .C1(_09537_ ), .C2(_09542_ ), .ZN(_09543_ ) );
AOI221_X4 _16061_ ( .A(_09533_ ), .B1(_09298_ ), .B2(_09531_ ), .C1(_09543_ ), .C2(_09412_ ), .ZN(_09544_ ) );
OAI221_X1 _16062_ ( .A(_09532_ ), .B1(_09440_ ), .B2(_09526_ ), .C1(_09544_ ), .C2(\exu.bge.io_is ), .ZN(_09545_ ) );
AOI221_X4 _16063_ ( .A(_09530_ ), .B1(_09444_ ), .B2(_09531_ ), .C1(_09545_ ), .C2(_09411_ ), .ZN(_09546_ ) );
OAI221_X1 _16064_ ( .A(_09527_ ), .B1(_09448_ ), .B2(_09529_ ), .C1(_09546_ ), .C2(\exu.beq.io_is ), .ZN(_09547_ ) );
NAND2_X1 _16065_ ( .A1(_09547_ ), .A2(_09409_ ), .ZN(_09548_ ) );
NAND2_X1 _16066_ ( .A1(fanout_net_9 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_9_A_$_MUX__A_B ), .ZN(_09549_ ) );
MUX2_X1 _16067_ ( .A(_09549_ ), .B(_09526_ ), .S(_09317_ ), .Z(_09550_ ) );
AND3_X1 _16068_ ( .A1(_09548_ ), .A2(\ifu.io_out_bits_pc_$_MUX__Y_9_A_$_MUX__Y_A_$_OR__Y_B_$_ANDNOT__Y_A ), .A3(_09550_ ), .ZN(_09551_ ) );
AOI211_X1 _16069_ ( .A(fanout_net_10 ), .B(_09551_ ), .C1(\exu.csrrs.io_csr_rdata [22] ), .C2(_09343_ ), .ZN(_09552_ ) );
AND3_X1 _16070_ ( .A1(_09513_ ), .A2(_09155_ ), .A3(_09153_ ), .ZN(_09553_ ) );
OAI21_X1 _16071_ ( .A(_09462_ ), .B1(_09553_ ), .B2(_09514_ ), .ZN(_09554_ ) );
NAND2_X1 _16072_ ( .A1(fanout_net_17 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_9_A_$_MUX__A_B ), .ZN(_09555_ ) );
AOI21_X1 _16073_ ( .A(_09321_ ), .B1(_09554_ ), .B2(_09555_ ), .ZN(_09556_ ) );
OAI21_X1 _16074_ ( .A(_09328_ ), .B1(_09552_ ), .B2(_09556_ ), .ZN(_09557_ ) );
INV_X1 _16075_ ( .A(\ifu.pc [22] ), .ZN(_09558_ ) );
OAI21_X1 _16076_ ( .A(_09558_ ), .B1(_09402_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_09559_ ) );
NAND2_X1 _16077_ ( .A1(_09557_ ), .A2(_09559_ ), .ZN(_09560_ ) );
NAND2_X1 _16078_ ( .A1(_09560_ ), .A2(_09466_ ), .ZN(_09561_ ) );
OAI21_X1 _16079_ ( .A(_09558_ ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09562_ ) );
NAND2_X1 _16080_ ( .A1(_09561_ ), .A2(_09562_ ), .ZN(_09563_ ) );
MUX2_X1 _16081_ ( .A(\icache.tag_reg_0 [17] ), .B(\icache.tag_reg_1 [17] ), .S(_09332_ ), .Z(_09564_ ) );
XOR2_X1 _16082_ ( .A(_09563_ ), .B(_09564_ ), .Z(_09565_ ) );
OAI21_X1 _16083_ ( .A(fanout_net_9 ), .B1(_09395_ ), .B2(\exu.addi._io_rd_T_4_$_NOT__Y_10_A_$_MUX__A_B ), .ZN(_09566_ ) );
AOI21_X1 _16084_ ( .A(_09476_ ), .B1(_08654_ ), .B2(_08678_ ), .ZN(_09567_ ) );
OR3_X1 _16085_ ( .A1(_09567_ ), .A2(_08661_ ), .A3(_08680_ ), .ZN(_09568_ ) );
OAI21_X1 _16086_ ( .A(_08661_ ), .B1(_09567_ ), .B2(_08680_ ), .ZN(_09569_ ) );
AND2_X1 _16087_ ( .A1(_09568_ ), .A2(_09569_ ), .ZN(_09570_ ) );
AOI21_X1 _16088_ ( .A(_09566_ ), .B1(_09570_ ), .B2(_09317_ ), .ZN(_09571_ ) );
OR2_X1 _16089_ ( .A1(_09570_ ), .A2(_08786_ ), .ZN(_09572_ ) );
AND3_X1 _16090_ ( .A1(_08798_ ), .A2(_08806_ ), .A3(_08803_ ), .ZN(_09573_ ) );
INV_X1 _16091_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_11_A_$_MUX__A_B ), .ZN(_09574_ ) );
NAND2_X1 _16092_ ( .A1(_09573_ ), .A2(_09574_ ), .ZN(_09575_ ) );
XNOR2_X1 _16093_ ( .A(_09575_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_10_A_$_MUX__A_B ), .ZN(_09576_ ) );
INV_X1 _16094_ ( .A(_09576_ ), .ZN(_09577_ ) );
AOI21_X1 _16095_ ( .A(_09202_ ), .B1(_09568_ ), .B2(_09569_ ), .ZN(_09578_ ) );
OR2_X1 _16096_ ( .A1(_09570_ ), .A2(_09440_ ), .ZN(_09579_ ) );
AOI21_X1 _16097_ ( .A(_08936_ ), .B1(_09568_ ), .B2(_09569_ ), .ZN(_09580_ ) );
INV_X1 _16098_ ( .A(_09488_ ), .ZN(_09581_ ) );
NAND3_X1 _16099_ ( .A1(_08957_ ), .A2(_08964_ ), .A3(_08962_ ), .ZN(_09582_ ) );
INV_X1 _16100_ ( .A(\exu.csrrs.io_csr_rdata [20] ), .ZN(_09583_ ) );
NOR2_X1 _16101_ ( .A1(_09582_ ), .A2(_09583_ ), .ZN(_09584_ ) );
OAI211_X1 _16102_ ( .A(_09581_ ), .B(_08972_ ), .C1(_09584_ ), .C2(\exu.csrrs.io_csr_rdata [21] ), .ZN(_09585_ ) );
AND2_X1 _16103_ ( .A1(\exu.addi._io_rd_T_4_$_NOT__Y_10_A_$_MUX__A_B ), .A2(fanout_net_11 ), .ZN(_09586_ ) );
OAI21_X1 _16104_ ( .A(_09585_ ), .B1(_08972_ ), .B2(_09586_ ), .ZN(_09587_ ) );
NOR2_X1 _16105_ ( .A1(_09576_ ), .A2(_09035_ ), .ZN(_09588_ ) );
OAI211_X1 _16106_ ( .A(_09587_ ), .B(_09254_ ), .C1(_09588_ ), .C2(fanout_net_11 ), .ZN(_09589_ ) );
AOI22_X1 _16107_ ( .A1(_09570_ ), .A2(_08945_ ), .B1(_09535_ ), .B2(_09577_ ), .ZN(_09590_ ) );
OAI211_X1 _16108_ ( .A(_09222_ ), .B(_09589_ ), .C1(_09590_ ), .C2(_09254_ ), .ZN(_09591_ ) );
MUX2_X1 _16109_ ( .A(_09577_ ), .B(_09570_ ), .S(_09220_ ), .Z(_09592_ ) );
OAI21_X1 _16110_ ( .A(_09591_ ), .B1(_09252_ ), .B2(_09592_ ), .ZN(_09593_ ) );
AOI221_X4 _16111_ ( .A(_09580_ ), .B1(_09298_ ), .B2(_09576_ ), .C1(_09593_ ), .C2(_09412_ ), .ZN(_09594_ ) );
OAI221_X1 _16112_ ( .A(_09579_ ), .B1(_08930_ ), .B2(_09577_ ), .C1(_09594_ ), .C2(\exu.bge.io_is ), .ZN(_09595_ ) );
AOI221_X4 _16113_ ( .A(_09578_ ), .B1(_09444_ ), .B2(_09576_ ), .C1(_09595_ ), .C2(_09411_ ), .ZN(_09596_ ) );
OAI221_X1 _16114_ ( .A(_09572_ ), .B1(_09448_ ), .B2(_09577_ ), .C1(_09596_ ), .C2(\exu.beq.io_is ), .ZN(_09597_ ) );
AOI21_X1 _16115_ ( .A(_09571_ ), .B1(_09597_ ), .B2(_09409_ ), .ZN(_09598_ ) );
AOI221_X4 _16116_ ( .A(fanout_net_10 ), .B1(\exu.csrrs.io_csr_rdata [21] ), .B2(_09343_ ), .C1(_09598_ ), .C2(\ifu.io_out_bits_pc_$_MUX__Y_9_A_$_MUX__Y_A_$_OR__Y_B_$_ANDNOT__Y_A ), .ZN(_09599_ ) );
AND2_X1 _16117_ ( .A1(_09138_ ), .A2(_09150_ ), .ZN(_09600_ ) );
NOR2_X1 _16118_ ( .A1(_09600_ ), .A2(_09148_ ), .ZN(_09601_ ) );
XNOR2_X1 _16119_ ( .A(_09601_ ), .B(_09147_ ), .ZN(\exu.addi._io_rd_T_4 [21] ) );
OR2_X1 _16120_ ( .A1(\exu.addi._io_rd_T_4 [21] ), .A2(fanout_net_17 ), .ZN(_09602_ ) );
NAND2_X1 _16121_ ( .A1(fanout_net_17 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_10_A_$_MUX__A_B ), .ZN(_09603_ ) );
AOI21_X1 _16122_ ( .A(_09321_ ), .B1(_09602_ ), .B2(_09603_ ), .ZN(_09604_ ) );
OAI21_X1 _16123_ ( .A(_09185_ ), .B1(_09599_ ), .B2(_09604_ ), .ZN(_09605_ ) );
INV_X1 _16124_ ( .A(\ifu.pc [21] ), .ZN(_09606_ ) );
OAI21_X1 _16125_ ( .A(_09606_ ), .B1(_09402_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_09607_ ) );
NAND2_X1 _16126_ ( .A1(_09605_ ), .A2(_09607_ ), .ZN(_09608_ ) );
NAND2_X1 _16127_ ( .A1(_09608_ ), .A2(_09183_ ), .ZN(_09609_ ) );
OAI21_X1 _16128_ ( .A(_09606_ ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09610_ ) );
AND2_X1 _16129_ ( .A1(_09609_ ), .A2(_09610_ ), .ZN(_09611_ ) );
MUX2_X1 _16130_ ( .A(\icache.tag_reg_0 [16] ), .B(\icache.tag_reg_1 [16] ), .S(_09332_ ), .Z(_09612_ ) );
XNOR2_X1 _16131_ ( .A(_09611_ ), .B(_09612_ ), .ZN(_09613_ ) );
XOR2_X1 _16132_ ( .A(_08685_ ), .B(_08686_ ), .Z(_09614_ ) );
AND2_X1 _16133_ ( .A1(_09614_ ), .A2(_09354_ ), .ZN(_09615_ ) );
INV_X1 _16134_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_7_A_$_MUX__A_B ), .ZN(_09616_ ) );
XNOR2_X1 _16135_ ( .A(_09265_ ), .B(_09616_ ), .ZN(_09617_ ) );
AOI211_X1 _16136_ ( .A(_09256_ ), .B(_09615_ ), .C1(_09257_ ), .C2(_09617_ ), .ZN(_09618_ ) );
INV_X1 _16137_ ( .A(_09617_ ), .ZN(_09619_ ) );
AND2_X1 _16138_ ( .A1(fanout_net_17 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_7_A_$_MUX__A_B ), .ZN(_09620_ ) );
OAI22_X1 _16139_ ( .A1(_09619_ ), .A2(_09210_ ), .B1(_09288_ ), .B2(_09620_ ), .ZN(_09621_ ) );
AND2_X1 _16140_ ( .A1(_09489_ ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_9_A_$_MUX__A_B_$_MUX__B_1_A_$_XOR__Y_A_$_NOR__A_Y_$_XOR__A_B ), .ZN(_09622_ ) );
NOR2_X1 _16141_ ( .A1(_09489_ ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_9_A_$_MUX__A_B_$_MUX__B_1_A_$_XOR__Y_A_$_NOR__A_Y_$_XOR__A_B ), .ZN(_09623_ ) );
OAI21_X1 _16142_ ( .A(_09414_ ), .B1(_09622_ ), .B2(_09623_ ), .ZN(_09624_ ) );
AOI21_X1 _16143_ ( .A(fanout_net_7 ), .B1(_09621_ ), .B2(_09624_ ), .ZN(_09625_ ) );
OAI21_X1 _16144_ ( .A(_09253_ ), .B1(_09618_ ), .B2(_09625_ ), .ZN(_09626_ ) );
NAND2_X1 _16145_ ( .A1(_09614_ ), .A2(_09293_ ), .ZN(_09627_ ) );
OAI211_X1 _16146_ ( .A(_09627_ ), .B(fanout_net_6 ), .C1(_09293_ ), .C2(_09619_ ), .ZN(_09628_ ) );
AOI21_X1 _16147_ ( .A(\exu.bgeu.io_is ), .B1(_09626_ ), .B2(_09628_ ), .ZN(_09629_ ) );
OAI22_X1 _16148_ ( .A1(_09614_ ), .A2(_09297_ ), .B1(_09299_ ), .B2(_09617_ ), .ZN(_09630_ ) );
OAI21_X1 _16149_ ( .A(_09251_ ), .B1(_09629_ ), .B2(_09630_ ), .ZN(_09631_ ) );
INV_X1 _16150_ ( .A(_09614_ ), .ZN(_09632_ ) );
AOI22_X1 _16151_ ( .A1(_09632_ ), .A2(_09303_ ), .B1(_08928_ ), .B2(_09619_ ), .ZN(_09633_ ) );
AOI21_X1 _16152_ ( .A(\exu.bne.io_is ), .B1(_09631_ ), .B2(_09633_ ), .ZN(_09634_ ) );
OAI22_X1 _16153_ ( .A1(_09614_ ), .A2(_09306_ ), .B1(_09309_ ), .B2(_09617_ ), .ZN(_09635_ ) );
OAI21_X1 _16154_ ( .A(_09249_ ), .B1(_09634_ ), .B2(_09635_ ), .ZN(_09636_ ) );
AOI22_X1 _16155_ ( .A1(_09632_ ), .A2(_09312_ ), .B1(_09313_ ), .B2(_09619_ ), .ZN(_09637_ ) );
AOI21_X1 _16156_ ( .A(fanout_net_9 ), .B1(_09636_ ), .B2(_09637_ ), .ZN(_09638_ ) );
OAI21_X1 _16157_ ( .A(fanout_net_9 ), .B1(_09396_ ), .B2(\exu.addi._io_rd_T_4_$_NOT__Y_7_A_$_MUX__A_B ), .ZN(_09639_ ) );
AOI21_X1 _16158_ ( .A(_09639_ ), .B1(_09614_ ), .B2(_09452_ ), .ZN(_09640_ ) );
NOR3_X1 _16159_ ( .A1(_09638_ ), .A2(fanout_net_8 ), .A3(_09640_ ), .ZN(_09641_ ) );
AOI211_X1 _16160_ ( .A(fanout_net_10 ), .B(_09641_ ), .C1(\exu.csrrs.io_csr_rdata [24] ), .C2(_08991_ ), .ZN(_09642_ ) );
NAND3_X1 _16161_ ( .A1(fanout_net_17 ), .A2(fanout_net_10 ), .A3(\exu.addi._io_rd_T_4_$_NOT__Y_7_A_$_MUX__A_B ), .ZN(_09643_ ) );
XNOR2_X1 _16162_ ( .A(_09160_ ), .B(_09322_ ), .ZN(\exu.addi._io_rd_T_4 [24] ) );
OAI21_X1 _16163_ ( .A(_09643_ ), .B1(\exu.addi._io_rd_T_4 [24] ), .B2(_09177_ ), .ZN(_09644_ ) );
OAI21_X1 _16164_ ( .A(_09328_ ), .B1(_09642_ ), .B2(_09644_ ), .ZN(_09645_ ) );
OAI21_X1 _16165_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_3_A_$_MUX__Y_B ), .B1(_09402_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_09646_ ) );
NAND3_X1 _16166_ ( .A1(_09645_ ), .A2(_09183_ ), .A3(_09646_ ), .ZN(_09647_ ) );
INV_X1 _16167_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_3_A_$_MUX__Y_B ), .ZN(_09648_ ) );
OAI21_X1 _16168_ ( .A(_09648_ ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09649_ ) );
NAND2_X1 _16169_ ( .A1(_09647_ ), .A2(_09649_ ), .ZN(_09650_ ) );
NOR2_X1 _16170_ ( .A1(_09332_ ), .A2(\icache.tag_reg_0 [19] ), .ZN(_09651_ ) );
AOI21_X1 _16171_ ( .A(\icache.tag_reg_1 [19] ), .B1(_09335_ ), .B2(_09337_ ), .ZN(_09652_ ) );
NOR2_X1 _16172_ ( .A1(_09651_ ), .A2(_09652_ ), .ZN(_09653_ ) );
XNOR2_X1 _16173_ ( .A(_09650_ ), .B(_09653_ ), .ZN(_09654_ ) );
AND4_X1 _16174_ ( .A1(_09525_ ), .A2(_09565_ ), .A3(_09613_ ), .A4(_09654_ ), .ZN(_09655_ ) );
NAND2_X1 _16175_ ( .A1(_09474_ ), .A2(_09655_ ), .ZN(_09656_ ) );
BUF_X4 _16176_ ( .A(_09321_ ), .Z(_09657_ ) );
XNOR2_X1 _16177_ ( .A(\exu.addi.io_imm [29] ), .B(\exu.auipc.io_rs1_data [29] ), .ZN(_09658_ ) );
AOI211_X1 _16178_ ( .A(_09658_ ), .B(_09352_ ), .C1(_09347_ ), .C2(_09350_ ), .ZN(_09659_ ) );
AND2_X1 _16179_ ( .A1(\exu.addi.io_imm [29] ), .A2(\exu.auipc.io_rs1_data [29] ), .ZN(_09660_ ) );
NAND2_X1 _16180_ ( .A1(\exu.addi.io_imm [28] ), .A2(\exu.auipc.io_rs1_data [28] ), .ZN(_09661_ ) );
NOR2_X1 _16181_ ( .A1(_09658_ ), .A2(_09661_ ), .ZN(_09662_ ) );
NOR3_X1 _16182_ ( .A1(_09659_ ), .A2(_09660_ ), .A3(_09662_ ), .ZN(_09663_ ) );
XNOR2_X1 _16183_ ( .A(\exu.addi.io_imm [30] ), .B(\exu.auipc.io_rs1_data [30] ), .ZN(_09664_ ) );
XOR2_X1 _16184_ ( .A(_09663_ ), .B(_09664_ ), .Z(_09665_ ) );
NAND2_X1 _16185_ ( .A1(_09665_ ), .A2(_09452_ ), .ZN(_09666_ ) );
INV_X1 _16186_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_1_A_$_MUX__A_B ), .ZN(_09667_ ) );
AOI21_X1 _16187_ ( .A(_09409_ ), .B1(fanout_net_17 ), .B2(_09667_ ), .ZN(_09668_ ) );
OR2_X1 _16188_ ( .A1(_09665_ ), .A2(_08786_ ), .ZN(_09669_ ) );
AND4_X1 _16189_ ( .A1(\exu.auipc.io_rs1_data [28] ), .A2(\exu.auipc.io_rs1_data [27] ), .A3(\exu.auipc.io_rs1_data [29] ), .A4(\exu.auipc.io_rs1_data [26] ), .ZN(_09670_ ) );
NAND3_X1 _16190_ ( .A1(_08804_ ), .A2(_08807_ ), .A3(_09670_ ), .ZN(_09671_ ) );
XNOR2_X1 _16191_ ( .A(_09671_ ), .B(_09667_ ), .ZN(_09672_ ) );
NOR2_X1 _16192_ ( .A1(_09665_ ), .A2(_09306_ ), .ZN(_09673_ ) );
INV_X1 _16193_ ( .A(_09672_ ), .ZN(_09674_ ) );
OR2_X1 _16194_ ( .A1(_09665_ ), .A2(_09440_ ), .ZN(_09675_ ) );
NOR2_X1 _16195_ ( .A1(_09665_ ), .A2(_09297_ ), .ZN(_09676_ ) );
NAND2_X1 _16196_ ( .A1(_09665_ ), .A2(_09220_ ), .ZN(_09677_ ) );
OAI211_X1 _16197_ ( .A(_09677_ ), .B(fanout_net_6 ), .C1(_09220_ ), .C2(_09674_ ), .ZN(_09678_ ) );
MUX2_X1 _16198_ ( .A(_09672_ ), .B(_09665_ ), .S(_08945_ ), .Z(_09679_ ) );
AND3_X1 _16199_ ( .A1(_09282_ ), .A2(\exu.csrrs.io_csr_rdata [24] ), .A3(\exu.csrrs.io_csr_rdata [23] ), .ZN(_09680_ ) );
AND3_X1 _16200_ ( .A1(_09680_ ), .A2(\exu.csrrs.io_csr_rdata [25] ), .A3(\exu.csrrs.io_csr_rdata [26] ), .ZN(_09681_ ) );
NAND3_X1 _16201_ ( .A1(_09681_ ), .A2(\exu.csrrs.io_csr_rdata [28] ), .A3(\exu.csrrs.io_csr_rdata [27] ), .ZN(_09682_ ) );
INV_X1 _16202_ ( .A(\exu.csrrs.io_csr_rdata [29] ), .ZN(_09683_ ) );
NOR2_X1 _16203_ ( .A1(_09682_ ), .A2(_09683_ ), .ZN(_09684_ ) );
AOI21_X1 _16204_ ( .A(_09214_ ), .B1(_09684_ ), .B2(\ifu.io_out_bits_pc_$_MUX__Y_13_A_$_MUX__Y_A_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ), .ZN(_09685_ ) );
OAI21_X1 _16205_ ( .A(_09685_ ), .B1(\ifu.io_out_bits_pc_$_MUX__Y_13_A_$_MUX__Y_A_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ), .B2(_09684_ ), .ZN(_09686_ ) );
AND2_X1 _16206_ ( .A1(fanout_net_17 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_1_A_$_MUX__A_B ), .ZN(_09687_ ) );
OAI22_X1 _16207_ ( .A1(_09674_ ), .A2(_09210_ ), .B1(_09211_ ), .B2(_09687_ ), .ZN(_09688_ ) );
AND2_X1 _16208_ ( .A1(_09686_ ), .A2(_09688_ ), .ZN(_09689_ ) );
MUX2_X1 _16209_ ( .A(_09679_ ), .B(_09689_ ), .S(_09255_ ), .Z(_09690_ ) );
OAI21_X1 _16210_ ( .A(_09678_ ), .B1(_09690_ ), .B2(fanout_net_6 ), .ZN(_09691_ ) );
AOI221_X4 _16211_ ( .A(_09676_ ), .B1(_09298_ ), .B2(_09674_ ), .C1(_09691_ ), .C2(_09413_ ), .ZN(_09692_ ) );
OAI221_X1 _16212_ ( .A(_09675_ ), .B1(_08930_ ), .B2(_09672_ ), .C1(_09692_ ), .C2(\exu.bge.io_is ), .ZN(_09693_ ) );
AOI221_X4 _16213_ ( .A(_09673_ ), .B1(_09444_ ), .B2(_09674_ ), .C1(_09693_ ), .C2(_09411_ ), .ZN(_09694_ ) );
OAI221_X1 _16214_ ( .A(_09669_ ), .B1(_09448_ ), .B2(_09672_ ), .C1(_09694_ ), .C2(\exu.beq.io_is ), .ZN(_09695_ ) );
AOI221_X4 _16215_ ( .A(_09342_ ), .B1(_09666_ ), .B2(_09668_ ), .C1(_09695_ ), .C2(_09409_ ), .ZN(_09696_ ) );
AND4_X1 _16216_ ( .A1(_09462_ ), .A2(_09342_ ), .A3(fanout_net_8 ), .A4(\exu.csrrs.io_csr_rdata [30] ), .ZN(_09697_ ) );
OAI21_X1 _16217_ ( .A(_09657_ ), .B1(_09696_ ), .B2(_09697_ ), .ZN(_09698_ ) );
AND2_X1 _16218_ ( .A1(\exu.add.io_rs1_data [29] ), .A2(\exu.addi.io_imm [29] ), .ZN(_09699_ ) );
NOR2_X1 _16219_ ( .A1(\exu.add.io_rs1_data [29] ), .A2(\exu.addi.io_imm [29] ), .ZN(_09700_ ) );
NOR2_X1 _16220_ ( .A1(_09699_ ), .A2(_09700_ ), .ZN(_09701_ ) );
INV_X1 _16221_ ( .A(_09701_ ), .ZN(_09702_ ) );
AOI211_X1 _16222_ ( .A(_09392_ ), .B(_09702_ ), .C1(_09386_ ), .C2(_09388_ ), .ZN(_09703_ ) );
INV_X1 _16223_ ( .A(\exu.addi.io_imm [28] ), .ZN(_09704_ ) );
NOR4_X1 _16224_ ( .A1(_09699_ ), .A2(_09700_ ), .A3(_08867_ ), .A4(_09704_ ), .ZN(_09705_ ) );
NOR3_X1 _16225_ ( .A1(_09703_ ), .A2(_09699_ ), .A3(_09705_ ), .ZN(_09706_ ) );
AND2_X1 _16226_ ( .A1(\exu.add.io_rs1_data [30] ), .A2(\exu.addi.io_imm [30] ), .ZN(_09707_ ) );
NOR2_X1 _16227_ ( .A1(\exu.add.io_rs1_data [30] ), .A2(\exu.addi.io_imm [30] ), .ZN(_09708_ ) );
NOR2_X1 _16228_ ( .A1(_09707_ ), .A2(_09708_ ), .ZN(_09709_ ) );
XNOR2_X1 _16229_ ( .A(_09706_ ), .B(_09709_ ), .ZN(\exu.addi._io_rd_T_4 [30] ) );
OR2_X1 _16230_ ( .A1(\exu.addi._io_rd_T_4 [30] ), .A2(_09177_ ), .ZN(_09710_ ) );
OAI211_X1 _16231_ ( .A(_09710_ ), .B(fanout_net_10 ), .C1(_09463_ ), .C2(_09667_ ), .ZN(_09711_ ) );
NAND3_X1 _16232_ ( .A1(_09698_ ), .A2(_09328_ ), .A3(_09711_ ), .ZN(_09712_ ) );
INV_X1 _16233_ ( .A(\ifu.pc [30] ), .ZN(_09713_ ) );
OAI21_X1 _16234_ ( .A(_09713_ ), .B1(_09402_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_09714_ ) );
NAND3_X1 _16235_ ( .A1(_09712_ ), .A2(_09466_ ), .A3(_09714_ ), .ZN(_09715_ ) );
OAI21_X1 _16236_ ( .A(\ifu.pc [30] ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09716_ ) );
AND2_X1 _16237_ ( .A1(_09715_ ), .A2(_09716_ ), .ZN(_09717_ ) );
NOR2_X1 _16238_ ( .A1(_09332_ ), .A2(\icache.tag_reg_0 [25] ), .ZN(_09718_ ) );
AOI21_X1 _16239_ ( .A(\icache.tag_reg_1 [25] ), .B1(_09335_ ), .B2(_09337_ ), .ZN(_09719_ ) );
OR2_X1 _16240_ ( .A1(_09718_ ), .A2(_09719_ ), .ZN(_09720_ ) );
XNOR2_X1 _16241_ ( .A(_09717_ ), .B(_09720_ ), .ZN(_09721_ ) );
NOR2_X1 _16242_ ( .A1(_09663_ ), .A2(_09664_ ), .ZN(_09722_ ) );
AND2_X1 _16243_ ( .A1(\exu.addi.io_imm [30] ), .A2(\exu.auipc.io_rs1_data [30] ), .ZN(_09723_ ) );
XNOR2_X1 _16244_ ( .A(\exu.addi.io_imm [31] ), .B(\exu.auipc.io_rs1_data [31] ), .ZN(_09724_ ) );
OR3_X1 _16245_ ( .A1(_09722_ ), .A2(_09723_ ), .A3(_09724_ ), .ZN(_09725_ ) );
OAI21_X1 _16246_ ( .A(_09724_ ), .B1(_09722_ ), .B2(_09723_ ), .ZN(_09726_ ) );
NAND2_X1 _16247_ ( .A1(_09725_ ), .A2(_09726_ ), .ZN(_09727_ ) );
NAND2_X1 _16248_ ( .A1(_09727_ ), .A2(_09354_ ), .ZN(_09728_ ) );
INV_X1 _16249_ ( .A(_08808_ ), .ZN(_09729_ ) );
NAND4_X1 _16250_ ( .A1(\exu.auipc.io_rs1_data [28] ), .A2(\exu.auipc.io_rs1_data [27] ), .A3(\exu.auipc.io_rs1_data [29] ), .A4(\exu.auipc.io_rs1_data [26] ), .ZN(_09730_ ) );
OR4_X1 _16251_ ( .A1(\exu.addi._io_rd_T_4_$_NOT__Y_1_A_$_MUX__A_B ), .A2(_09729_ ), .A3(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_MUX__A_B ), .A4(_09730_ ), .ZN(_09731_ ) );
OAI21_X1 _16252_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_MUX__A_B ), .B1(_09671_ ), .B2(\exu.addi._io_rd_T_4_$_NOT__Y_1_A_$_MUX__A_B ), .ZN(_09732_ ) );
NAND2_X1 _16253_ ( .A1(_09731_ ), .A2(_09732_ ), .ZN(_09733_ ) );
OAI211_X1 _16254_ ( .A(_09728_ ), .B(fanout_net_7 ), .C1(_09733_ ), .C2(_09354_ ), .ZN(_09734_ ) );
INV_X1 _16255_ ( .A(_09733_ ), .ZN(_09735_ ) );
AND2_X1 _16256_ ( .A1(fanout_net_17 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_MUX__A_B ), .ZN(_09736_ ) );
INV_X1 _16257_ ( .A(_09736_ ), .ZN(_09737_ ) );
AOI22_X1 _16258_ ( .A1(_09735_ ), .A2(_09209_ ), .B1(fanout_net_11 ), .B2(_09737_ ), .ZN(_09738_ ) );
AND4_X1 _16259_ ( .A1(\exu.csrrs.io_csr_rdata [28] ), .A2(\exu.csrrs.io_csr_rdata [29] ), .A3(\exu.csrrs.io_csr_rdata [27] ), .A4(\exu.csrrs.io_csr_rdata [26] ), .ZN(_09739_ ) );
NAND3_X1 _16260_ ( .A1(_08969_ ), .A2(\exu.csrrs.io_csr_rdata [30] ), .A3(_09739_ ), .ZN(_09740_ ) );
INV_X1 _16261_ ( .A(\exu.csrrs.io_csr_rdata [31] ), .ZN(_09741_ ) );
NAND2_X1 _16262_ ( .A1(_09740_ ), .A2(_09741_ ), .ZN(_09742_ ) );
NAND4_X1 _16263_ ( .A1(_08969_ ), .A2(\exu.csrrs.io_csr_rdata [30] ), .A3(\exu.csrrs.io_csr_rdata [31] ), .A4(_09739_ ), .ZN(_09743_ ) );
AOI21_X1 _16264_ ( .A(_09271_ ), .B1(_09742_ ), .B2(_09743_ ), .ZN(_09744_ ) );
OAI21_X1 _16265_ ( .A(_09256_ ), .B1(_09738_ ), .B2(_09744_ ), .ZN(_09745_ ) );
AOI21_X1 _16266_ ( .A(fanout_net_6 ), .B1(_09734_ ), .B2(_09745_ ), .ZN(_09746_ ) );
AOI21_X1 _16267_ ( .A(_09432_ ), .B1(_09725_ ), .B2(_09726_ ), .ZN(_09747_ ) );
AOI211_X1 _16268_ ( .A(_09253_ ), .B(_09747_ ), .C1(_09735_ ), .C2(_09432_ ), .ZN(_09748_ ) );
OAI21_X1 _16269_ ( .A(_09413_ ), .B1(_09746_ ), .B2(_09748_ ), .ZN(_09749_ ) );
INV_X1 _16270_ ( .A(_09727_ ), .ZN(_09750_ ) );
AOI22_X1 _16271_ ( .A1(_09750_ ), .A2(_09437_ ), .B1(_09733_ ), .B2(_09298_ ), .ZN(_09751_ ) );
AOI21_X1 _16272_ ( .A(\exu.bge.io_is ), .B1(_09749_ ), .B2(_09751_ ), .ZN(_09752_ ) );
OAI22_X1 _16273_ ( .A1(_09727_ ), .A2(_09440_ ), .B1(_09735_ ), .B2(_08930_ ), .ZN(_09753_ ) );
OAI21_X1 _16274_ ( .A(_09411_ ), .B1(_09752_ ), .B2(_09753_ ), .ZN(_09754_ ) );
AOI22_X1 _16275_ ( .A1(_09750_ ), .A2(_09443_ ), .B1(_09733_ ), .B2(_09444_ ), .ZN(_09755_ ) );
AOI21_X1 _16276_ ( .A(\exu.beq.io_is ), .B1(_09754_ ), .B2(_09755_ ), .ZN(_09756_ ) );
NAND3_X1 _16277_ ( .A1(_09725_ ), .A2(_09726_ ), .A3(_09312_ ), .ZN(_09757_ ) );
OAI21_X1 _16278_ ( .A(_09757_ ), .B1(_09735_ ), .B2(_09448_ ), .ZN(_09758_ ) );
OAI21_X1 _16279_ ( .A(_09409_ ), .B1(_09756_ ), .B2(_09758_ ), .ZN(_09759_ ) );
OAI21_X1 _16280_ ( .A(_09737_ ), .B1(_09727_ ), .B2(fanout_net_17 ), .ZN(_09760_ ) );
AOI21_X1 _16281_ ( .A(_09342_ ), .B1(_09760_ ), .B2(fanout_net_9 ), .ZN(_09761_ ) );
AOI22_X1 _16282_ ( .A1(_09759_ ), .A2(_09761_ ), .B1(\exu.csrrs.io_csr_rdata [31] ), .B2(_09343_ ), .ZN(_09762_ ) );
NOR2_X1 _16283_ ( .A1(_09762_ ), .A2(fanout_net_10 ), .ZN(_09763_ ) );
NOR3_X1 _16284_ ( .A1(_09706_ ), .A2(_09707_ ), .A3(_09708_ ), .ZN(_09764_ ) );
NOR2_X1 _16285_ ( .A1(_09764_ ), .A2(_09707_ ), .ZN(_09765_ ) );
XOR2_X1 _16286_ ( .A(\exu.add.io_rs1_data [31] ), .B(\exu.addi.io_imm [31] ), .Z(_09766_ ) );
XNOR2_X1 _16287_ ( .A(_09765_ ), .B(_09766_ ), .ZN(\exu.addi._io_rd_T_4 [31] ) );
NOR2_X1 _16288_ ( .A1(\exu.addi._io_rd_T_4 [31] ), .A2(_09177_ ), .ZN(_09767_ ) );
AOI211_X1 _16289_ ( .A(_09321_ ), .B(_09767_ ), .C1(fanout_net_17 ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_MUX__A_B ), .ZN(_09768_ ) );
OR3_X1 _16290_ ( .A1(_09763_ ), .A2(_09040_ ), .A3(_09768_ ), .ZN(_09769_ ) );
OAI211_X1 _16291_ ( .A(_09769_ ), .B(_09466_ ), .C1(\ifu.pc [31] ), .C2(_09328_ ), .ZN(_09770_ ) );
OAI21_X1 _16292_ ( .A(\ifu.pc [31] ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09771_ ) );
AND2_X1 _16293_ ( .A1(_09770_ ), .A2(_09771_ ), .ZN(_09772_ ) );
MUX2_X1 _16294_ ( .A(\icache.tag_reg_0 [26] ), .B(\icache.tag_reg_1 [26] ), .S(_09332_ ), .Z(_09773_ ) );
XOR2_X1 _16295_ ( .A(_09772_ ), .B(_09773_ ), .Z(_09774_ ) );
BUF_X4 _16296_ ( .A(_09328_ ), .Z(_09775_ ) );
NAND2_X1 _16297_ ( .A1(fanout_net_17 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_2_A_$_MUX__A_B ), .ZN(_09776_ ) );
NOR2_X1 _16298_ ( .A1(_09394_ ), .A2(_09389_ ), .ZN(_09777_ ) );
XNOR2_X1 _16299_ ( .A(_09777_ ), .B(_09702_ ), .ZN(_09778_ ) );
INV_X1 _16300_ ( .A(_09778_ ), .ZN(\exu.addi._io_rd_T_4 [29] ) );
OAI211_X1 _16301_ ( .A(fanout_net_10 ), .B(_09776_ ), .C1(\exu.addi._io_rd_T_4 [29] ), .C2(fanout_net_18 ), .ZN(_09779_ ) );
OR2_X1 _16302_ ( .A1(_09351_ ), .A2(_09352_ ), .ZN(_09780_ ) );
NAND2_X1 _16303_ ( .A1(_09780_ ), .A2(_09661_ ), .ZN(_09781_ ) );
XNOR2_X1 _16304_ ( .A(_09781_ ), .B(_09658_ ), .ZN(_09782_ ) );
NAND2_X1 _16305_ ( .A1(_09782_ ), .A2(_09354_ ), .ZN(_09783_ ) );
INV_X1 _16306_ ( .A(_09356_ ), .ZN(_09784_ ) );
OAI21_X1 _16307_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_2_A_$_MUX__A_B ), .B1(_09784_ ), .B2(\exu.addi._io_rd_T_4_$_NOT__Y_3_A_$_MUX__A_B ), .ZN(_09785_ ) );
INV_X1 _16308_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_2_A_$_MUX__A_B ), .ZN(_09786_ ) );
NAND3_X1 _16309_ ( .A1(_09356_ ), .A2(_09786_ ), .A3(_09382_ ), .ZN(_09787_ ) );
NAND2_X1 _16310_ ( .A1(_09785_ ), .A2(_09787_ ), .ZN(_09788_ ) );
OAI211_X1 _16311_ ( .A(_09783_ ), .B(fanout_net_7 ), .C1(_09354_ ), .C2(_09788_ ), .ZN(_09789_ ) );
AND2_X1 _16312_ ( .A1(_08969_ ), .A2(_09739_ ), .ZN(_09790_ ) );
NAND2_X1 _16313_ ( .A1(_09360_ ), .A2(\exu.csrrs.io_csr_rdata [28] ), .ZN(_09791_ ) );
AOI211_X1 _16314_ ( .A(_09271_ ), .B(_09790_ ), .C1(_09791_ ), .C2(_09683_ ), .ZN(_09792_ ) );
AOI211_X1 _16315_ ( .A(_09288_ ), .B(_09792_ ), .C1(_09786_ ), .C2(_09271_ ), .ZN(_09793_ ) );
INV_X1 _16316_ ( .A(_09788_ ), .ZN(_09794_ ) );
AOI21_X1 _16317_ ( .A(fanout_net_11 ), .B1(_09794_ ), .B2(exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ), .ZN(_09795_ ) );
OAI21_X1 _16318_ ( .A(_09256_ ), .B1(_09793_ ), .B2(_09795_ ), .ZN(_09796_ ) );
NAND3_X1 _16319_ ( .A1(_09789_ ), .A2(_09253_ ), .A3(_09796_ ), .ZN(_09797_ ) );
INV_X1 _16320_ ( .A(_08979_ ), .ZN(_09798_ ) );
AOI22_X1 _16321_ ( .A1(_09782_ ), .A2(_09293_ ), .B1(_09798_ ), .B2(_09794_ ), .ZN(_09799_ ) );
OAI211_X1 _16322_ ( .A(_09797_ ), .B(_09413_ ), .C1(_09253_ ), .C2(_09799_ ), .ZN(_09800_ ) );
INV_X1 _16323_ ( .A(_09782_ ), .ZN(_09801_ ) );
AOI22_X1 _16324_ ( .A1(_09801_ ), .A2(_09437_ ), .B1(_09298_ ), .B2(_09788_ ), .ZN(_09802_ ) );
AOI21_X1 _16325_ ( .A(\exu.bge.io_is ), .B1(_09800_ ), .B2(_09802_ ), .ZN(_09803_ ) );
OAI22_X1 _16326_ ( .A1(_09782_ ), .A2(_09440_ ), .B1(_08930_ ), .B2(_09794_ ), .ZN(_09804_ ) );
OAI21_X1 _16327_ ( .A(_09411_ ), .B1(_09803_ ), .B2(_09804_ ), .ZN(_09805_ ) );
AOI22_X1 _16328_ ( .A1(_09801_ ), .A2(_09443_ ), .B1(_09444_ ), .B2(_09788_ ), .ZN(_09806_ ) );
AOI21_X1 _16329_ ( .A(\exu.beq.io_is ), .B1(_09805_ ), .B2(_09806_ ), .ZN(_09807_ ) );
OAI22_X1 _16330_ ( .A1(_09782_ ), .A2(_08786_ ), .B1(_09448_ ), .B2(_09794_ ), .ZN(_09808_ ) );
OAI21_X1 _16331_ ( .A(_09410_ ), .B1(_09807_ ), .B2(_09808_ ), .ZN(_09809_ ) );
OAI21_X1 _16332_ ( .A(_09776_ ), .B1(_09782_ ), .B2(fanout_net_18 ), .ZN(_09810_ ) );
AOI21_X1 _16333_ ( .A(_09342_ ), .B1(_09810_ ), .B2(fanout_net_9 ), .ZN(_09811_ ) );
AOI22_X1 _16334_ ( .A1(_09809_ ), .A2(_09811_ ), .B1(\exu.csrrs.io_csr_rdata [29] ), .B2(_09343_ ), .ZN(_09812_ ) );
OAI211_X1 _16335_ ( .A(_09775_ ), .B(_09779_ ), .C1(_09812_ ), .C2(fanout_net_10 ), .ZN(_09813_ ) );
INV_X1 _16336_ ( .A(\ifu.pc [29] ), .ZN(_09814_ ) );
OAI21_X1 _16337_ ( .A(_09814_ ), .B1(_09402_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_09815_ ) );
NAND3_X1 _16338_ ( .A1(_09813_ ), .A2(_09466_ ), .A3(_09815_ ), .ZN(_09816_ ) );
OAI21_X1 _16339_ ( .A(\ifu.pc [29] ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09817_ ) );
BUF_X4 _16340_ ( .A(_09332_ ), .Z(_09818_ ) );
NAND2_X1 _16341_ ( .A1(_09818_ ), .A2(\icache.tag_reg_1 [24] ), .ZN(_09819_ ) );
NAND3_X1 _16342_ ( .A1(_09335_ ), .A2(\icache.tag_reg_0 [24] ), .A3(_09337_ ), .ZN(_09820_ ) );
AOI22_X1 _16343_ ( .A1(_09816_ ), .A2(_09817_ ), .B1(_09819_ ), .B2(_09820_ ), .ZN(_09821_ ) );
AND4_X1 _16344_ ( .A1(_09816_ ), .A2(_09817_ ), .A3(_09819_ ), .A4(_09820_ ), .ZN(_09822_ ) );
OAI211_X1 _16345_ ( .A(_09721_ ), .B(_09774_ ), .C1(_09821_ ), .C2(_09822_ ), .ZN(_09823_ ) );
NOR2_X1 _16346_ ( .A1(_08625_ ), .A2(_08642_ ), .ZN(_09824_ ) );
INV_X1 _16347_ ( .A(_08631_ ), .ZN(_09825_ ) );
INV_X1 _16348_ ( .A(_08632_ ), .ZN(_09826_ ) );
NOR3_X1 _16349_ ( .A1(_09824_ ), .A2(_09825_ ), .A3(_09826_ ), .ZN(_09827_ ) );
OAI21_X1 _16350_ ( .A(_08627_ ), .B1(_09827_ ), .B2(_08650_ ), .ZN(_09828_ ) );
INV_X1 _16351_ ( .A(_08644_ ), .ZN(_09829_ ) );
AND2_X1 _16352_ ( .A1(_09828_ ), .A2(_09829_ ), .ZN(_09830_ ) );
XOR2_X1 _16353_ ( .A(_09830_ ), .B(_08626_ ), .Z(_09831_ ) );
OR2_X1 _16354_ ( .A1(_09831_ ), .A2(_08786_ ), .ZN(_09832_ ) );
AND3_X1 _16355_ ( .A1(_08798_ ), .A2(\exu.auipc.io_rs1_data [14] ), .A3(_08801_ ), .ZN(_09833_ ) );
INV_X1 _16356_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_16_A_$_MUX__A_B ), .ZN(_09834_ ) );
XNOR2_X1 _16357_ ( .A(_09833_ ), .B(_09834_ ), .ZN(_09835_ ) );
NOR3_X1 _16358_ ( .A1(_09443_ ), .A2(_08984_ ), .A3(_09835_ ), .ZN(_09836_ ) );
INV_X1 _16359_ ( .A(_09831_ ), .ZN(_09837_ ) );
OR2_X1 _16360_ ( .A1(_09831_ ), .A2(_08926_ ), .ZN(_09838_ ) );
NOR3_X1 _16361_ ( .A1(_08935_ ), .A2(_08931_ ), .A3(_09835_ ), .ZN(_09839_ ) );
INV_X1 _16362_ ( .A(_09835_ ), .ZN(_09840_ ) );
OAI211_X1 _16363_ ( .A(fanout_net_6 ), .B(_09840_ ), .C1(_08921_ ), .C2(fanout_net_18 ), .ZN(_09841_ ) );
AOI21_X1 _16364_ ( .A(fanout_net_11 ), .B1(_09840_ ), .B2(exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ), .ZN(_09842_ ) );
XNOR2_X1 _16365_ ( .A(_09275_ ), .B(\exu.csrrs.io_csr_rdata [15] ), .ZN(_09843_ ) );
MUX2_X1 _16366_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_16_A_$_MUX__A_B ), .B(_09843_ ), .S(_08972_ ), .Z(_09844_ ) );
AOI211_X1 _16367_ ( .A(fanout_net_7 ), .B(_09842_ ), .C1(_09844_ ), .C2(fanout_net_11 ), .ZN(_09845_ ) );
MUX2_X1 _16368_ ( .A(_09840_ ), .B(_09837_ ), .S(_08943_ ), .Z(_09846_ ) );
AOI21_X1 _16369_ ( .A(_09845_ ), .B1(_09846_ ), .B2(fanout_net_7 ), .ZN(_09847_ ) );
OAI221_X1 _16370_ ( .A(_09841_ ), .B1(_08977_ ), .B2(_09831_ ), .C1(_09847_ ), .C2(fanout_net_6 ), .ZN(_09848_ ) );
AOI221_X4 _16371_ ( .A(_09839_ ), .B1(_08935_ ), .B2(_09837_ ), .C1(_09848_ ), .C2(_09412_ ), .ZN(_09849_ ) );
OAI221_X1 _16372_ ( .A(_09838_ ), .B1(_08930_ ), .B2(_09835_ ), .C1(_09849_ ), .C2(\exu.bge.io_is ), .ZN(_09850_ ) );
AOI221_X4 _16373_ ( .A(_09836_ ), .B1(_09443_ ), .B2(_09837_ ), .C1(_09850_ ), .C2(_08984_ ), .ZN(_09851_ ) );
OAI221_X1 _16374_ ( .A(_09832_ ), .B1(_09448_ ), .B2(_09835_ ), .C1(_09851_ ), .C2(\exu.beq.io_is ), .ZN(_09852_ ) );
NAND2_X1 _16375_ ( .A1(_09852_ ), .A2(_09409_ ), .ZN(_09853_ ) );
NAND2_X1 _16376_ ( .A1(_09831_ ), .A2(_09317_ ), .ZN(_09854_ ) );
OAI211_X1 _16377_ ( .A(_09854_ ), .B(fanout_net_9 ), .C1(_09395_ ), .C2(_09834_ ), .ZN(_09855_ ) );
AOI21_X1 _16378_ ( .A(fanout_net_8 ), .B1(_09853_ ), .B2(_09855_ ), .ZN(_09856_ ) );
AOI211_X1 _16379_ ( .A(fanout_net_10 ), .B(_09856_ ), .C1(\exu.csrrs.io_csr_rdata [15] ), .C2(_08991_ ), .ZN(_09857_ ) );
OAI21_X1 _16380_ ( .A(_09115_ ), .B1(_09094_ ), .B2(_09101_ ), .ZN(_09858_ ) );
AOI21_X1 _16381_ ( .A(_09118_ ), .B1(_09858_ ), .B2(_09117_ ), .ZN(_09859_ ) );
NOR2_X1 _16382_ ( .A1(_09859_ ), .A2(_09106_ ), .ZN(_09860_ ) );
XNOR2_X1 _16383_ ( .A(_09860_ ), .B(_09105_ ), .ZN(\exu.addi._io_rd_T_4 [15] ) );
NOR2_X1 _16384_ ( .A1(\exu.addi._io_rd_T_4 [15] ), .A2(fanout_net_18 ), .ZN(_09861_ ) );
AND2_X1 _16385_ ( .A1(fanout_net_18 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_16_A_$_MUX__A_B ), .ZN(_09862_ ) );
OAI21_X1 _16386_ ( .A(fanout_net_10 ), .B1(_09861_ ), .B2(_09862_ ), .ZN(_09863_ ) );
INV_X1 _16387_ ( .A(_09863_ ), .ZN(_09864_ ) );
OR3_X1 _16388_ ( .A1(_09857_ ), .A2(_09040_ ), .A3(_09864_ ), .ZN(_09865_ ) );
OAI21_X1 _16389_ ( .A(\ifu.pc [15] ), .B1(_09402_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_09866_ ) );
NAND3_X1 _16390_ ( .A1(_09865_ ), .A2(_09183_ ), .A3(_09866_ ), .ZN(_09867_ ) );
OR2_X1 _16391_ ( .A1(_09182_ ), .A2(\ifu.pc [15] ), .ZN(_09868_ ) );
NAND2_X1 _16392_ ( .A1(_09867_ ), .A2(_09868_ ), .ZN(_09869_ ) );
INV_X1 _16393_ ( .A(_09245_ ), .ZN(_09870_ ) );
OR2_X1 _16394_ ( .A1(_09870_ ), .A2(\icache.tag_reg_1 [10] ), .ZN(_09871_ ) );
OR2_X1 _16395_ ( .A1(_09246_ ), .A2(\icache.tag_reg_0 [10] ), .ZN(_09872_ ) );
AND3_X1 _16396_ ( .A1(_09869_ ), .A2(_09871_ ), .A3(_09872_ ), .ZN(_09873_ ) );
AOI21_X1 _16397_ ( .A(_09869_ ), .B1(_09871_ ), .B2(_09872_ ), .ZN(_09874_ ) );
NOR2_X1 _16398_ ( .A1(_08634_ ), .A2(_08653_ ), .ZN(_09875_ ) );
XNOR2_X1 _16399_ ( .A(_09875_ ), .B(_08579_ ), .ZN(_09876_ ) );
INV_X1 _16400_ ( .A(_09876_ ), .ZN(_09877_ ) );
AND2_X1 _16401_ ( .A1(_09220_ ), .A2(_09877_ ), .ZN(_09878_ ) );
AND3_X1 _16402_ ( .A1(_08798_ ), .A2(_08802_ ), .A3(_08801_ ), .ZN(_09879_ ) );
XNOR2_X1 _16403_ ( .A(_09879_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_15_A_$_MUX__A_B ), .ZN(_09880_ ) );
INV_X1 _16404_ ( .A(_09880_ ), .ZN(_09881_ ) );
AOI211_X1 _16405_ ( .A(_09252_ ), .B(_09878_ ), .C1(_09432_ ), .C2(_09881_ ), .ZN(_09882_ ) );
OR2_X1 _16406_ ( .A1(_09876_ ), .A2(_09207_ ), .ZN(_09883_ ) );
OAI211_X1 _16407_ ( .A(_09883_ ), .B(fanout_net_7 ), .C1(_09354_ ), .C2(_09880_ ), .ZN(_09884_ ) );
AND2_X1 _16408_ ( .A1(_09880_ ), .A2(exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ), .ZN(_09885_ ) );
XNOR2_X1 _16409_ ( .A(_09276_ ), .B(\exu.csrrs.io_csr_rdata [16] ), .ZN(_09886_ ) );
NOR2_X1 _16410_ ( .A1(_09886_ ), .A2(_09271_ ), .ZN(_09887_ ) );
OAI21_X1 _16411_ ( .A(fanout_net_11 ), .B1(_09191_ ), .B2(\exu.addi._io_rd_T_4_$_NOT__Y_15_A_$_MUX__A_B ), .ZN(_09888_ ) );
OAI221_X1 _16412_ ( .A(_09255_ ), .B1(fanout_net_11 ), .B2(_09885_ ), .C1(_09887_ ), .C2(_09888_ ), .ZN(_09889_ ) );
AOI21_X1 _16413_ ( .A(fanout_net_6 ), .B1(_09884_ ), .B2(_09889_ ), .ZN(_09890_ ) );
OAI21_X1 _16414_ ( .A(_09413_ ), .B1(_09882_ ), .B2(_09890_ ), .ZN(_09891_ ) );
OR2_X1 _16415_ ( .A1(_09876_ ), .A2(_09297_ ), .ZN(_09892_ ) );
OAI211_X1 _16416_ ( .A(_09892_ ), .B(\exu.bgeu.io_is ), .C1(_09437_ ), .C2(_09880_ ), .ZN(_09893_ ) );
AOI21_X1 _16417_ ( .A(\exu.bge.io_is ), .B1(_09891_ ), .B2(_09893_ ), .ZN(_09894_ ) );
OAI22_X1 _16418_ ( .A1(_08930_ ), .A2(_09881_ ), .B1(_09440_ ), .B2(_09877_ ), .ZN(_09895_ ) );
OAI21_X1 _16419_ ( .A(_09411_ ), .B1(_09894_ ), .B2(_09895_ ), .ZN(_09896_ ) );
AOI22_X1 _16420_ ( .A1(_09876_ ), .A2(_09443_ ), .B1(_09444_ ), .B2(_09880_ ), .ZN(_09897_ ) );
AOI21_X1 _16421_ ( .A(\exu.beq.io_is ), .B1(_09896_ ), .B2(_09897_ ), .ZN(_09898_ ) );
NAND2_X1 _16422_ ( .A1(_09876_ ), .A2(_08784_ ), .ZN(_09899_ ) );
OAI21_X1 _16423_ ( .A(_09899_ ), .B1(_09448_ ), .B2(_09881_ ), .ZN(_09900_ ) );
OAI21_X1 _16424_ ( .A(_08702_ ), .B1(_09898_ ), .B2(_09900_ ), .ZN(_09901_ ) );
INV_X1 _16425_ ( .A(_08699_ ), .ZN(_09902_ ) );
OR2_X1 _16426_ ( .A1(_09876_ ), .A2(_09902_ ), .ZN(_09903_ ) );
INV_X1 _16427_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_15_A_$_MUX__A_B ), .ZN(_09904_ ) );
OAI211_X1 _16428_ ( .A(_09903_ ), .B(fanout_net_9 ), .C1(_09395_ ), .C2(_09904_ ), .ZN(_09905_ ) );
AOI21_X1 _16429_ ( .A(fanout_net_8 ), .B1(_09901_ ), .B2(_09905_ ), .ZN(_09906_ ) );
AOI211_X1 _16430_ ( .A(fanout_net_10 ), .B(_09906_ ), .C1(\exu.csrrs.io_csr_rdata [16] ), .C2(_08991_ ), .ZN(_09907_ ) );
INV_X1 _16431_ ( .A(_09126_ ), .ZN(_09908_ ) );
XNOR2_X1 _16432_ ( .A(_09123_ ), .B(_09908_ ), .ZN(\exu.addi._io_rd_T_4 [16] ) );
NOR2_X1 _16433_ ( .A1(\exu.addi._io_rd_T_4 [16] ), .A2(fanout_net_18 ), .ZN(_09909_ ) );
AND2_X1 _16434_ ( .A1(fanout_net_18 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_15_A_$_MUX__A_B ), .ZN(_09910_ ) );
OAI21_X1 _16435_ ( .A(fanout_net_10 ), .B1(_09909_ ), .B2(_09910_ ), .ZN(_09911_ ) );
INV_X1 _16436_ ( .A(_09911_ ), .ZN(_09912_ ) );
OR3_X1 _16437_ ( .A1(_09907_ ), .A2(_09040_ ), .A3(_09912_ ), .ZN(_09913_ ) );
OAI21_X1 _16438_ ( .A(\ifu.pc [16] ), .B1(_09401_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_09914_ ) );
NAND3_X1 _16439_ ( .A1(_09913_ ), .A2(_09182_ ), .A3(_09914_ ), .ZN(_09915_ ) );
INV_X1 _16440_ ( .A(\ifu.pc [16] ), .ZN(_09916_ ) );
OAI21_X1 _16441_ ( .A(_09916_ ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_09917_ ) );
NAND2_X1 _16442_ ( .A1(_09915_ ), .A2(_09917_ ), .ZN(_09918_ ) );
MUX2_X1 _16443_ ( .A(\icache.tag_reg_0 [11] ), .B(\icache.tag_reg_1 [11] ), .S(_09245_ ), .Z(_09919_ ) );
XNOR2_X1 _16444_ ( .A(_09918_ ), .B(_09919_ ), .ZN(_09920_ ) );
OR3_X1 _16445_ ( .A1(_09873_ ), .A2(_09874_ ), .A3(_09920_ ), .ZN(_09921_ ) );
OAI21_X1 _16446_ ( .A(_08581_ ), .B1(_08634_ ), .B2(_08653_ ), .ZN(_09922_ ) );
NAND2_X1 _16447_ ( .A1(_09922_ ), .A2(_08671_ ), .ZN(_09923_ ) );
NAND2_X1 _16448_ ( .A1(_09923_ ), .A2(_08583_ ), .ZN(_09924_ ) );
AND2_X1 _16449_ ( .A1(_09924_ ), .A2(_08676_ ), .ZN(_09925_ ) );
XNOR2_X1 _16450_ ( .A(_09925_ ), .B(_08582_ ), .ZN(_09926_ ) );
AND2_X1 _16451_ ( .A1(_09926_ ), .A2(_08945_ ), .ZN(_09927_ ) );
NAND3_X1 _16452_ ( .A1(_08798_ ), .A2(\exu.auipc.io_rs1_data [18] ), .A3(_08803_ ), .ZN(_09928_ ) );
XNOR2_X1 _16453_ ( .A(_09928_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_12_A_$_MUX__A_B ), .ZN(_09929_ ) );
INV_X1 _16454_ ( .A(_09929_ ), .ZN(_09930_ ) );
AOI211_X1 _16455_ ( .A(_09255_ ), .B(_09927_ ), .C1(_09257_ ), .C2(_09930_ ), .ZN(_09931_ ) );
OAI21_X1 _16456_ ( .A(_09288_ ), .B1(_09929_ ), .B2(_09036_ ), .ZN(_09932_ ) );
AND3_X1 _16457_ ( .A1(_08957_ ), .A2(\exu.csrrs.io_csr_rdata [18] ), .A3(_08962_ ), .ZN(_09933_ ) );
OAI211_X1 _16458_ ( .A(_09414_ ), .B(_09582_ ), .C1(_09933_ ), .C2(\exu.csrrs.io_csr_rdata [19] ), .ZN(_09934_ ) );
OAI211_X1 _16459_ ( .A(_09934_ ), .B(fanout_net_11 ), .C1(_09191_ ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_12_A_$_MUX__A_B ), .ZN(_09935_ ) );
AOI21_X1 _16460_ ( .A(fanout_net_7 ), .B1(_09932_ ), .B2(_09935_ ), .ZN(_09936_ ) );
OAI21_X1 _16461_ ( .A(_09252_ ), .B1(_09931_ ), .B2(_09936_ ), .ZN(_09937_ ) );
NAND2_X1 _16462_ ( .A1(_09926_ ), .A2(_09220_ ), .ZN(_09938_ ) );
OAI211_X1 _16463_ ( .A(_09938_ ), .B(fanout_net_6 ), .C1(_08979_ ), .C2(_09929_ ), .ZN(_09939_ ) );
AOI21_X1 _16464_ ( .A(\exu.bgeu.io_is ), .B1(_09937_ ), .B2(_09939_ ), .ZN(_09940_ ) );
OAI211_X1 _16465_ ( .A(\exu.bgeu.io_is ), .B(_09929_ ), .C1(_09428_ ), .C2(fanout_net_18 ), .ZN(_09941_ ) );
OAI21_X1 _16466_ ( .A(_09941_ ), .B1(_09926_ ), .B2(_09297_ ), .ZN(_09942_ ) );
OAI21_X1 _16467_ ( .A(_09251_ ), .B1(_09940_ ), .B2(_09942_ ), .ZN(_09943_ ) );
BUF_X2 _16468_ ( .A(_08921_ ), .Z(_09944_ ) );
AOI211_X1 _16469_ ( .A(_09250_ ), .B(_09930_ ), .C1(_09944_ ), .C2(_09192_ ), .ZN(_09945_ ) );
INV_X1 _16470_ ( .A(_09926_ ), .ZN(_09946_ ) );
AOI21_X1 _16471_ ( .A(_09945_ ), .B1(_09946_ ), .B2(_09303_ ), .ZN(_09947_ ) );
AOI21_X1 _16472_ ( .A(\exu.bne.io_is ), .B1(_09943_ ), .B2(_09947_ ), .ZN(_09948_ ) );
OAI22_X1 _16473_ ( .A1(_09926_ ), .A2(_09306_ ), .B1(_09309_ ), .B2(_09930_ ), .ZN(_09949_ ) );
OAI21_X1 _16474_ ( .A(_09249_ ), .B1(_09948_ ), .B2(_09949_ ), .ZN(_09950_ ) );
AOI22_X1 _16475_ ( .A1(_09946_ ), .A2(_09312_ ), .B1(_09313_ ), .B2(_09929_ ), .ZN(_09951_ ) );
AOI21_X1 _16476_ ( .A(fanout_net_9 ), .B1(_09950_ ), .B2(_09951_ ), .ZN(_09952_ ) );
AND2_X1 _16477_ ( .A1(fanout_net_9 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_12_A_$_MUX__A_B ), .ZN(_09953_ ) );
MUX2_X1 _16478_ ( .A(_09953_ ), .B(_09946_ ), .S(_09317_ ), .Z(_09954_ ) );
NOR3_X1 _16479_ ( .A1(_09952_ ), .A2(_09342_ ), .A3(_09954_ ), .ZN(_09955_ ) );
AOI211_X1 _16480_ ( .A(fanout_net_10 ), .B(_09955_ ), .C1(\exu.csrrs.io_csr_rdata [19] ), .C2(_09343_ ), .ZN(_09956_ ) );
AOI21_X1 _16481_ ( .A(_09908_ ), .B1(_09116_ ), .B2(_09122_ ), .ZN(_09957_ ) );
OR2_X1 _16482_ ( .A1(_09957_ ), .A2(_09124_ ), .ZN(_09958_ ) );
AOI21_X1 _16483_ ( .A(_09127_ ), .B1(_09958_ ), .B2(_09131_ ), .ZN(_09959_ ) );
NOR2_X1 _16484_ ( .A1(_09959_ ), .A2(_09133_ ), .ZN(_09960_ ) );
NOR2_X1 _16485_ ( .A1(_09960_ ), .A2(_09046_ ), .ZN(_09961_ ) );
XNOR2_X1 _16486_ ( .A(_09961_ ), .B(_09045_ ), .ZN(\exu.addi._io_rd_T_4 [19] ) );
OR2_X1 _16487_ ( .A1(\exu.addi._io_rd_T_4 [19] ), .A2(fanout_net_18 ), .ZN(_09962_ ) );
NAND2_X1 _16488_ ( .A1(fanout_net_18 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_12_A_$_MUX__A_B ), .ZN(_09963_ ) );
AOI21_X1 _16489_ ( .A(_09042_ ), .B1(_09962_ ), .B2(_09963_ ), .ZN(_09964_ ) );
OR3_X1 _16490_ ( .A1(_09956_ ), .A2(_09040_ ), .A3(_09964_ ), .ZN(_09965_ ) );
OAI21_X1 _16491_ ( .A(\ifu.pc [19] ), .B1(_09401_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_09966_ ) );
NAND3_X1 _16492_ ( .A1(_09965_ ), .A2(_09182_ ), .A3(_09966_ ), .ZN(_09967_ ) );
OR2_X1 _16493_ ( .A1(_09182_ ), .A2(\ifu.pc [19] ), .ZN(_09968_ ) );
NAND2_X1 _16494_ ( .A1(_09967_ ), .A2(_09968_ ), .ZN(_09969_ ) );
MUX2_X1 _16495_ ( .A(\icache.tag_reg_0 [14] ), .B(\icache.tag_reg_1 [14] ), .S(_09245_ ), .Z(_09970_ ) );
XOR2_X1 _16496_ ( .A(_09969_ ), .B(_09970_ ), .Z(_09971_ ) );
XNOR2_X1 _16497_ ( .A(_09923_ ), .B(_08672_ ), .ZN(_09972_ ) );
NOR2_X1 _16498_ ( .A1(_09972_ ), .A2(_09257_ ), .ZN(_09973_ ) );
INV_X1 _16499_ ( .A(\exu.auipc.io_rs1_data [18] ), .ZN(_09974_ ) );
XNOR2_X1 _16500_ ( .A(_08804_ ), .B(_09974_ ), .ZN(_09975_ ) );
INV_X1 _16501_ ( .A(_09975_ ), .ZN(_09976_ ) );
AOI211_X1 _16502_ ( .A(_09255_ ), .B(_09973_ ), .C1(_09257_ ), .C2(_09976_ ), .ZN(_09977_ ) );
AOI21_X1 _16503_ ( .A(\exu.csrrs.io_csr_rdata [18] ), .B1(_08957_ ), .B2(_08962_ ), .ZN(_09978_ ) );
NOR3_X1 _16504_ ( .A1(_09933_ ), .A2(_09978_ ), .A3(_09271_ ), .ZN(_09979_ ) );
INV_X1 _16505_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_13_A_$_MUX__A_B ), .ZN(_09980_ ) );
AOI211_X1 _16506_ ( .A(_09288_ ), .B(_09979_ ), .C1(fanout_net_18 ), .C2(_09980_ ), .ZN(_09981_ ) );
NAND2_X1 _16507_ ( .A1(_09975_ ), .A2(exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ), .ZN(_09982_ ) );
AOI211_X1 _16508_ ( .A(fanout_net_7 ), .B(_09981_ ), .C1(_09288_ ), .C2(_09982_ ), .ZN(_09983_ ) );
OR3_X1 _16509_ ( .A1(_09977_ ), .A2(fanout_net_6 ), .A3(_09983_ ), .ZN(_09984_ ) );
NOR2_X1 _16510_ ( .A1(_09972_ ), .A2(_09432_ ), .ZN(_09985_ ) );
AOI21_X1 _16511_ ( .A(_09985_ ), .B1(_09798_ ), .B2(_09976_ ), .ZN(_09986_ ) );
OAI211_X1 _16512_ ( .A(_09984_ ), .B(_09413_ ), .C1(_09253_ ), .C2(_09986_ ), .ZN(_09987_ ) );
OR2_X1 _16513_ ( .A1(_09972_ ), .A2(_09297_ ), .ZN(_09988_ ) );
OAI211_X1 _16514_ ( .A(_09988_ ), .B(\exu.bgeu.io_is ), .C1(_09437_ ), .C2(_09975_ ), .ZN(_09989_ ) );
AOI21_X1 _16515_ ( .A(\exu.bge.io_is ), .B1(_09987_ ), .B2(_09989_ ), .ZN(_09990_ ) );
NOR4_X1 _16516_ ( .A1(_09972_ ), .A2(fanout_net_18 ), .A3(_09251_ ), .A4(_08920_ ), .ZN(_09991_ ) );
AOI211_X1 _16517_ ( .A(_09251_ ), .B(_09991_ ), .C1(_09440_ ), .C2(_09976_ ), .ZN(_09992_ ) );
OAI21_X1 _16518_ ( .A(_09411_ ), .B1(_09990_ ), .B2(_09992_ ), .ZN(_09993_ ) );
AOI22_X1 _16519_ ( .A1(_09972_ ), .A2(_09443_ ), .B1(_09444_ ), .B2(_09975_ ), .ZN(_09994_ ) );
AOI21_X1 _16520_ ( .A(\exu.beq.io_is ), .B1(_09993_ ), .B2(_09994_ ), .ZN(_09995_ ) );
NAND2_X1 _16521_ ( .A1(_09972_ ), .A2(_09312_ ), .ZN(_09996_ ) );
OAI21_X1 _16522_ ( .A(_09996_ ), .B1(_09448_ ), .B2(_09976_ ), .ZN(_09997_ ) );
OAI21_X1 _16523_ ( .A(_09409_ ), .B1(_09995_ ), .B2(_09997_ ), .ZN(_09998_ ) );
BUF_X2 _16524_ ( .A(_09902_ ), .Z(_09999_ ) );
OR2_X1 _16525_ ( .A1(_09972_ ), .A2(_09999_ ), .ZN(_10000_ ) );
OAI211_X1 _16526_ ( .A(_10000_ ), .B(fanout_net_9 ), .C1(_09396_ ), .C2(_09980_ ), .ZN(_10001_ ) );
AOI21_X1 _16527_ ( .A(fanout_net_8 ), .B1(_09998_ ), .B2(_10001_ ), .ZN(_10002_ ) );
AND3_X1 _16528_ ( .A1(_09396_ ), .A2(fanout_net_8 ), .A3(\exu.csrrs.io_csr_rdata [18] ), .ZN(_10003_ ) );
OAI21_X1 _16529_ ( .A(_09321_ ), .B1(_10002_ ), .B2(_10003_ ), .ZN(_10004_ ) );
XNOR2_X1 _16530_ ( .A(_09959_ ), .B(_09048_ ), .ZN(\exu.addi._io_rd_T_4 [18] ) );
OR2_X1 _16531_ ( .A1(\exu.addi._io_rd_T_4 [18] ), .A2(_09177_ ), .ZN(_10005_ ) );
OAI211_X1 _16532_ ( .A(_10005_ ), .B(fanout_net_10 ), .C1(_09462_ ), .C2(_09980_ ), .ZN(_10006_ ) );
NAND2_X1 _16533_ ( .A1(_10004_ ), .A2(_10006_ ), .ZN(_10007_ ) );
NAND2_X1 _16534_ ( .A1(_10007_ ), .A2(_09185_ ), .ZN(_10008_ ) );
OAI21_X1 _16535_ ( .A(\ifu.pc [18] ), .B1(_09402_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_10009_ ) );
NAND3_X1 _16536_ ( .A1(_10008_ ), .A2(_09183_ ), .A3(_10009_ ), .ZN(_10010_ ) );
INV_X1 _16537_ ( .A(\ifu.pc [18] ), .ZN(_10011_ ) );
OAI21_X1 _16538_ ( .A(_10011_ ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10012_ ) );
NAND2_X1 _16539_ ( .A1(_10010_ ), .A2(_10012_ ), .ZN(_10013_ ) );
NAND2_X1 _16540_ ( .A1(_09246_ ), .A2(\icache.tag_reg_1 [13] ), .ZN(_10014_ ) );
NAND3_X1 _16541_ ( .A1(_09335_ ), .A2(\icache.tag_reg_0 [13] ), .A3(_09337_ ), .ZN(_10015_ ) );
AND2_X1 _16542_ ( .A1(_10014_ ), .A2(_10015_ ), .ZN(_10016_ ) );
XNOR2_X1 _16543_ ( .A(_10013_ ), .B(_10016_ ), .ZN(_10017_ ) );
XNOR2_X1 _16544_ ( .A(_09475_ ), .B(_08658_ ), .ZN(_10018_ ) );
OR2_X1 _16545_ ( .A1(_10018_ ), .A2(_09257_ ), .ZN(_10019_ ) );
XNOR2_X1 _16546_ ( .A(_09573_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_11_A_$_MUX__A_B ), .ZN(_10020_ ) );
OAI211_X1 _16547_ ( .A(_10019_ ), .B(fanout_net_7 ), .C1(_09354_ ), .C2(_10020_ ), .ZN(_10021_ ) );
AOI21_X1 _16548_ ( .A(fanout_net_11 ), .B1(_10020_ ), .B2(exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ), .ZN(_10022_ ) );
AND3_X1 _16549_ ( .A1(_08957_ ), .A2(_08964_ ), .A3(_08962_ ), .ZN(_10023_ ) );
NAND2_X1 _16550_ ( .A1(_10023_ ), .A2(\exu.csrrs.io_csr_rdata [20] ), .ZN(_10024_ ) );
NAND2_X1 _16551_ ( .A1(_09582_ ), .A2(_09583_ ), .ZN(_10025_ ) );
AOI21_X1 _16552_ ( .A(_09271_ ), .B1(_10024_ ), .B2(_10025_ ), .ZN(_10026_ ) );
AND3_X1 _16553_ ( .A1(fanout_net_18 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_11_A_$_MUX__A_B ), .A3(fanout_net_11 ), .ZN(_10027_ ) );
OR4_X1 _16554_ ( .A1(fanout_net_7 ), .A2(_10022_ ), .A3(_10026_ ), .A4(_10027_ ), .ZN(_10028_ ) );
AOI21_X1 _16555_ ( .A(fanout_net_6 ), .B1(_10021_ ), .B2(_10028_ ), .ZN(_10029_ ) );
NOR2_X1 _16556_ ( .A1(_10018_ ), .A2(_09432_ ), .ZN(_10030_ ) );
INV_X1 _16557_ ( .A(_10020_ ), .ZN(_10031_ ) );
AOI211_X1 _16558_ ( .A(_09252_ ), .B(_10030_ ), .C1(_09432_ ), .C2(_10031_ ), .ZN(_10032_ ) );
OAI21_X1 _16559_ ( .A(_09413_ ), .B1(_10029_ ), .B2(_10032_ ), .ZN(_10033_ ) );
AOI22_X1 _16560_ ( .A1(_10018_ ), .A2(_09437_ ), .B1(_09298_ ), .B2(_10020_ ), .ZN(_10034_ ) );
AOI21_X1 _16561_ ( .A(\exu.bge.io_is ), .B1(_10033_ ), .B2(_10034_ ), .ZN(_10035_ ) );
NAND2_X1 _16562_ ( .A1(_10018_ ), .A2(_09303_ ), .ZN(_10036_ ) );
OAI21_X1 _16563_ ( .A(_10036_ ), .B1(_08930_ ), .B2(_10031_ ), .ZN(_10037_ ) );
OAI21_X1 _16564_ ( .A(_09411_ ), .B1(_10035_ ), .B2(_10037_ ), .ZN(_10038_ ) );
AOI22_X1 _16565_ ( .A1(_10018_ ), .A2(_09443_ ), .B1(_09444_ ), .B2(_10020_ ), .ZN(_10039_ ) );
AOI21_X1 _16566_ ( .A(\exu.beq.io_is ), .B1(_10038_ ), .B2(_10039_ ), .ZN(_10040_ ) );
NAND2_X1 _16567_ ( .A1(_10018_ ), .A2(_09312_ ), .ZN(_10041_ ) );
OAI21_X1 _16568_ ( .A(_10041_ ), .B1(_09448_ ), .B2(_10031_ ), .ZN(_10042_ ) );
OAI21_X1 _16569_ ( .A(_09409_ ), .B1(_10040_ ), .B2(_10042_ ), .ZN(_10043_ ) );
OR2_X1 _16570_ ( .A1(_10018_ ), .A2(_09999_ ), .ZN(_10044_ ) );
OAI211_X1 _16571_ ( .A(_10044_ ), .B(fanout_net_9 ), .C1(_09395_ ), .C2(_09574_ ), .ZN(_10045_ ) );
AOI21_X1 _16572_ ( .A(fanout_net_8 ), .B1(_10043_ ), .B2(_10045_ ), .ZN(_10046_ ) );
AOI211_X1 _16573_ ( .A(fanout_net_10 ), .B(_10046_ ), .C1(\exu.csrrs.io_csr_rdata [20] ), .C2(_08991_ ), .ZN(_10047_ ) );
XOR2_X1 _16574_ ( .A(_09138_ ), .B(_09150_ ), .Z(\exu.addi._io_rd_T_4 [20] ) );
NOR2_X1 _16575_ ( .A1(\exu.addi._io_rd_T_4 [20] ), .A2(fanout_net_18 ), .ZN(_10048_ ) );
AND2_X1 _16576_ ( .A1(fanout_net_18 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_11_A_$_MUX__A_B ), .ZN(_10049_ ) );
OAI21_X1 _16577_ ( .A(fanout_net_10 ), .B1(_10048_ ), .B2(_10049_ ), .ZN(_10050_ ) );
INV_X1 _16578_ ( .A(_10050_ ), .ZN(_10051_ ) );
OR3_X1 _16579_ ( .A1(_10047_ ), .A2(_09040_ ), .A3(_10051_ ), .ZN(_10052_ ) );
OAI21_X1 _16580_ ( .A(\ifu.pc [20] ), .B1(_09402_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_10053_ ) );
NAND3_X1 _16581_ ( .A1(_10052_ ), .A2(_09183_ ), .A3(_10053_ ), .ZN(_10054_ ) );
INV_X1 _16582_ ( .A(\ifu.pc [20] ), .ZN(_10055_ ) );
OAI21_X1 _16583_ ( .A(_10055_ ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10056_ ) );
NAND2_X1 _16584_ ( .A1(_10054_ ), .A2(_10056_ ), .ZN(_10057_ ) );
NAND2_X1 _16585_ ( .A1(_09246_ ), .A2(\icache.tag_reg_1 [15] ), .ZN(_10058_ ) );
NAND3_X1 _16586_ ( .A1(_09334_ ), .A2(\icache.tag_reg_0 [15] ), .A3(_09336_ ), .ZN(_10059_ ) );
AND2_X1 _16587_ ( .A1(_10058_ ), .A2(_10059_ ), .ZN(_10060_ ) );
XNOR2_X1 _16588_ ( .A(_10057_ ), .B(_10060_ ), .ZN(_10061_ ) );
AND2_X1 _16589_ ( .A1(fanout_net_11 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_14_A_$_MUX__A_B ), .ZN(_10062_ ) );
XNOR2_X1 _16590_ ( .A(_09277_ ), .B(\exu.csrrs.io_csr_rdata [17] ), .ZN(_10063_ ) );
MUX2_X1 _16591_ ( .A(_10062_ ), .B(_10063_ ), .S(_09414_ ), .Z(_10064_ ) );
NAND2_X1 _16592_ ( .A1(_09879_ ), .A2(_09904_ ), .ZN(_10065_ ) );
XNOR2_X1 _16593_ ( .A(_10065_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_14_A_$_MUX__A_B ), .ZN(_10066_ ) );
NOR2_X1 _16594_ ( .A1(_10066_ ), .A2(_09036_ ), .ZN(_10067_ ) );
OAI21_X1 _16595_ ( .A(_09255_ ), .B1(_10067_ ), .B2(fanout_net_11 ), .ZN(_10068_ ) );
NOR2_X1 _16596_ ( .A1(\exu.addi.io_imm [16] ), .A2(\exu.auipc.io_rs1_data [16] ), .ZN(_10069_ ) );
NOR3_X1 _16597_ ( .A1(_09875_ ), .A2(_08669_ ), .A3(_10069_ ), .ZN(_10070_ ) );
NOR2_X1 _16598_ ( .A1(_10070_ ), .A2(_08669_ ), .ZN(_10071_ ) );
XNOR2_X1 _16599_ ( .A(_10071_ ), .B(_08580_ ), .ZN(_10072_ ) );
INV_X1 _16600_ ( .A(_10066_ ), .ZN(_10073_ ) );
AOI22_X1 _16601_ ( .A1(_10072_ ), .A2(_09354_ ), .B1(_09535_ ), .B2(_10073_ ), .ZN(_10074_ ) );
OAI221_X1 _16602_ ( .A(_09252_ ), .B1(_10064_ ), .B2(_10068_ ), .C1(_10074_ ), .C2(_09256_ ), .ZN(_10075_ ) );
NAND2_X1 _16603_ ( .A1(_10072_ ), .A2(_09220_ ), .ZN(_10076_ ) );
OAI211_X1 _16604_ ( .A(_10076_ ), .B(fanout_net_6 ), .C1(_09293_ ), .C2(_10066_ ), .ZN(_10077_ ) );
AOI21_X1 _16605_ ( .A(\exu.bgeu.io_is ), .B1(_10075_ ), .B2(_10077_ ), .ZN(_10078_ ) );
OAI22_X1 _16606_ ( .A1(_10072_ ), .A2(_09297_ ), .B1(_09299_ ), .B2(_10073_ ), .ZN(_10079_ ) );
OAI21_X1 _16607_ ( .A(_09251_ ), .B1(_10078_ ), .B2(_10079_ ), .ZN(_10080_ ) );
NAND2_X1 _16608_ ( .A1(_10072_ ), .A2(_09303_ ), .ZN(_10081_ ) );
OAI211_X1 _16609_ ( .A(_10081_ ), .B(\exu.bge.io_is ), .C1(_09303_ ), .C2(_10066_ ), .ZN(_10082_ ) );
AOI21_X1 _16610_ ( .A(\exu.bne.io_is ), .B1(_10080_ ), .B2(_10082_ ), .ZN(_10083_ ) );
OAI22_X1 _16611_ ( .A1(_10072_ ), .A2(_09306_ ), .B1(_09309_ ), .B2(_10073_ ), .ZN(_10084_ ) );
OAI21_X1 _16612_ ( .A(_09249_ ), .B1(_10083_ ), .B2(_10084_ ), .ZN(_10085_ ) );
INV_X1 _16613_ ( .A(_10072_ ), .ZN(_10086_ ) );
AOI22_X1 _16614_ ( .A1(_10086_ ), .A2(_09312_ ), .B1(_09313_ ), .B2(_10066_ ), .ZN(_10087_ ) );
AOI21_X1 _16615_ ( .A(fanout_net_9 ), .B1(_10085_ ), .B2(_10087_ ), .ZN(_10088_ ) );
AND2_X1 _16616_ ( .A1(fanout_net_9 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_14_A_$_MUX__A_B ), .ZN(_10089_ ) );
MUX2_X1 _16617_ ( .A(_10089_ ), .B(_10086_ ), .S(_09317_ ), .Z(_10090_ ) );
NOR3_X1 _16618_ ( .A1(_10088_ ), .A2(_09342_ ), .A3(_10090_ ), .ZN(_10091_ ) );
AOI211_X1 _16619_ ( .A(fanout_net_10 ), .B(_10091_ ), .C1(\exu.csrrs.io_csr_rdata [17] ), .C2(_09343_ ), .ZN(_10092_ ) );
XNOR2_X1 _16620_ ( .A(_09958_ ), .B(_09129_ ), .ZN(_10093_ ) );
AND2_X1 _16621_ ( .A1(_10093_ ), .A2(_09396_ ), .ZN(_10094_ ) );
AND2_X1 _16622_ ( .A1(fanout_net_18 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_14_A_$_MUX__A_B ), .ZN(_10095_ ) );
OAI21_X1 _16623_ ( .A(fanout_net_10 ), .B1(_10094_ ), .B2(_10095_ ), .ZN(_10096_ ) );
INV_X1 _16624_ ( .A(_10096_ ), .ZN(_10097_ ) );
OAI21_X1 _16625_ ( .A(_09185_ ), .B1(_10092_ ), .B2(_10097_ ), .ZN(_10098_ ) );
INV_X1 _16626_ ( .A(\ifu.pc [17] ), .ZN(_10099_ ) );
OAI21_X1 _16627_ ( .A(_10099_ ), .B1(_09401_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_10100_ ) );
NAND2_X1 _16628_ ( .A1(_10098_ ), .A2(_10100_ ), .ZN(_10101_ ) );
NAND2_X1 _16629_ ( .A1(_10101_ ), .A2(_09183_ ), .ZN(_10102_ ) );
OAI21_X1 _16630_ ( .A(_10099_ ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10103_ ) );
NAND2_X1 _16631_ ( .A1(_10102_ ), .A2(_10103_ ), .ZN(_10104_ ) );
NAND2_X1 _16632_ ( .A1(_09246_ ), .A2(\icache.tag_reg_1 [12] ), .ZN(_10105_ ) );
NAND3_X1 _16633_ ( .A1(_09334_ ), .A2(\icache.tag_reg_0 [12] ), .A3(_09336_ ), .ZN(_10106_ ) );
AND2_X1 _16634_ ( .A1(_10105_ ), .A2(_10106_ ), .ZN(_10107_ ) );
XNOR2_X1 _16635_ ( .A(_10104_ ), .B(_10107_ ), .ZN(_10108_ ) );
NAND4_X1 _16636_ ( .A1(_09971_ ), .A2(_10017_ ), .A3(_10061_ ), .A4(_10108_ ), .ZN(_10109_ ) );
AOI21_X1 _16637_ ( .A(_09220_ ), .B1(_08947_ ), .B2(_08943_ ), .ZN(_10110_ ) );
INV_X1 _16638_ ( .A(_10110_ ), .ZN(_10111_ ) );
AOI21_X1 _16639_ ( .A(_08935_ ), .B1(_10111_ ), .B2(_09412_ ), .ZN(_10112_ ) );
INV_X1 _16640_ ( .A(_10112_ ), .ZN(_10113_ ) );
OR3_X1 _16641_ ( .A1(_09827_ ), .A2(_08627_ ), .A3(_08650_ ), .ZN(_10114_ ) );
AND2_X1 _16642_ ( .A1(_10114_ ), .A2(_09828_ ), .ZN(_10115_ ) );
NAND2_X1 _16643_ ( .A1(fanout_net_11 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_17_A_$_MUX__A_B ), .ZN(_10116_ ) );
XOR2_X1 _16644_ ( .A(_09274_ ), .B(\exu.csrrs.io_csr_rdata [14] ), .Z(_10117_ ) );
MUX2_X1 _16645_ ( .A(_10116_ ), .B(_10117_ ), .S(_09414_ ), .Z(_10118_ ) );
AND2_X1 _16646_ ( .A1(_08798_ ), .A2(_08801_ ), .ZN(_10119_ ) );
INV_X1 _16647_ ( .A(\exu.auipc.io_rs1_data [14] ), .ZN(_10120_ ) );
XNOR2_X1 _16648_ ( .A(_10119_ ), .B(_10120_ ), .ZN(_10121_ ) );
AOI21_X1 _16649_ ( .A(fanout_net_11 ), .B1(_10121_ ), .B2(exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ), .ZN(_10122_ ) );
NOR4_X1 _16650_ ( .A1(_10122_ ), .A2(\exu.bgeu.io_is ), .A3(fanout_net_6 ), .A4(fanout_net_7 ), .ZN(_10123_ ) );
AOI22_X1 _16651_ ( .A1(_10113_ ), .A2(_10115_ ), .B1(_10118_ ), .B2(_10123_ ), .ZN(_10124_ ) );
OAI21_X1 _16652_ ( .A(fanout_net_6 ), .B1(_09944_ ), .B2(fanout_net_18 ), .ZN(_10125_ ) );
NAND3_X1 _16653_ ( .A1(_09207_ ), .A2(_09222_ ), .A3(fanout_net_7 ), .ZN(_10126_ ) );
AOI21_X1 _16654_ ( .A(\exu.bgeu.io_is ), .B1(_10125_ ), .B2(_10126_ ), .ZN(_10127_ ) );
OAI21_X1 _16655_ ( .A(_10121_ ), .B1(_10127_ ), .B2(_09298_ ), .ZN(_10128_ ) );
AOI21_X1 _16656_ ( .A(\exu.bge.io_is ), .B1(_10124_ ), .B2(_10128_ ), .ZN(_10129_ ) );
AOI21_X1 _16657_ ( .A(_08926_ ), .B1(_09828_ ), .B2(_10114_ ), .ZN(_10130_ ) );
INV_X1 _16658_ ( .A(_10121_ ), .ZN(_10131_ ) );
AOI211_X1 _16659_ ( .A(_09250_ ), .B(_10130_ ), .C1(_08926_ ), .C2(_10131_ ), .ZN(_10132_ ) );
OAI21_X1 _16660_ ( .A(_08984_ ), .B1(_10129_ ), .B2(_10132_ ), .ZN(_10133_ ) );
AOI22_X1 _16661_ ( .A1(_10115_ ), .A2(_09443_ ), .B1(_09307_ ), .B2(_10121_ ), .ZN(_10134_ ) );
AOI21_X1 _16662_ ( .A(\exu.beq.io_is ), .B1(_10133_ ), .B2(_10134_ ), .ZN(_10135_ ) );
NAND3_X1 _16663_ ( .A1(_10114_ ), .A2(_08784_ ), .A3(_09828_ ), .ZN(_10136_ ) );
OAI21_X1 _16664_ ( .A(_10136_ ), .B1(_08790_ ), .B2(_10131_ ), .ZN(_10137_ ) );
OAI21_X1 _16665_ ( .A(_08702_ ), .B1(_10135_ ), .B2(_10137_ ), .ZN(_10138_ ) );
AND2_X1 _16666_ ( .A1(fanout_net_18 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_17_A_$_MUX__A_B ), .ZN(_10139_ ) );
INV_X1 _16667_ ( .A(_10139_ ), .ZN(_10140_ ) );
OAI211_X1 _16668_ ( .A(fanout_net_9 ), .B(_10140_ ), .C1(_10115_ ), .C2(fanout_net_18 ), .ZN(_10141_ ) );
AOI21_X1 _16669_ ( .A(fanout_net_8 ), .B1(_10138_ ), .B2(_10141_ ), .ZN(_10142_ ) );
AOI211_X1 _16670_ ( .A(fanout_net_10 ), .B(_10142_ ), .C1(\exu.csrrs.io_csr_rdata [14] ), .C2(_08990_ ), .ZN(_10143_ ) );
AND3_X1 _16671_ ( .A1(_09858_ ), .A2(_09118_ ), .A3(_09117_ ), .ZN(_10144_ ) );
NOR2_X1 _16672_ ( .A1(_10144_ ), .A2(_09859_ ), .ZN(\exu.addi._io_rd_T_4 [14] ) );
NOR2_X1 _16673_ ( .A1(\exu.addi._io_rd_T_4 [14] ), .A2(fanout_net_18 ), .ZN(_10145_ ) );
OAI21_X1 _16674_ ( .A(fanout_net_10 ), .B1(_10145_ ), .B2(_10139_ ), .ZN(_10146_ ) );
INV_X1 _16675_ ( .A(_10146_ ), .ZN(_10147_ ) );
OR3_X1 _16676_ ( .A1(_10143_ ), .A2(_09039_ ), .A3(_10147_ ), .ZN(_10148_ ) );
OAI21_X1 _16677_ ( .A(\ifu.pc [14] ), .B1(_09401_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_10149_ ) );
NAND3_X1 _16678_ ( .A1(_10148_ ), .A2(_09181_ ), .A3(_10149_ ), .ZN(_10150_ ) );
INV_X1 _16679_ ( .A(\ifu.pc [14] ), .ZN(_10151_ ) );
OAI21_X1 _16680_ ( .A(_10151_ ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10152_ ) );
NAND2_X1 _16681_ ( .A1(_10150_ ), .A2(_10152_ ), .ZN(_10153_ ) );
MUX2_X1 _16682_ ( .A(\icache.tag_reg_0 [9] ), .B(\icache.tag_reg_1 [9] ), .S(_09246_ ), .Z(_10154_ ) );
XOR2_X1 _16683_ ( .A(_10153_ ), .B(_10154_ ), .Z(_10155_ ) );
NOR2_X1 _16684_ ( .A1(_09824_ ), .A2(_09826_ ), .ZN(_10156_ ) );
OR3_X1 _16685_ ( .A1(_10156_ ), .A2(_09825_ ), .A3(_08646_ ), .ZN(_10157_ ) );
OAI21_X1 _16686_ ( .A(_09825_ ), .B1(_10156_ ), .B2(_08646_ ), .ZN(_10158_ ) );
AOI21_X1 _16687_ ( .A(_08786_ ), .B1(_10157_ ), .B2(_10158_ ), .ZN(_10159_ ) );
INV_X1 _16688_ ( .A(_08798_ ), .ZN(_10160_ ) );
NOR2_X1 _16689_ ( .A1(_10160_ ), .A2(_08799_ ), .ZN(_10161_ ) );
INV_X1 _16690_ ( .A(_10161_ ), .ZN(_10162_ ) );
NOR2_X1 _16691_ ( .A1(_10162_ ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_19_A_$_MUX__A_B ), .ZN(_10163_ ) );
INV_X1 _16692_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_18_A_$_MUX__A_B ), .ZN(_10164_ ) );
XNOR2_X1 _16693_ ( .A(_10163_ ), .B(_10164_ ), .ZN(_10165_ ) );
INV_X1 _16694_ ( .A(_10165_ ), .ZN(_10166_ ) );
NAND3_X1 _16695_ ( .A1(_09207_ ), .A2(fanout_net_7 ), .A3(_10166_ ), .ZN(_10167_ ) );
OAI21_X1 _16696_ ( .A(_09211_ ), .B1(_10165_ ), .B2(_09036_ ), .ZN(_10168_ ) );
INV_X1 _16697_ ( .A(_09274_ ), .ZN(_10169_ ) );
AND4_X1 _16698_ ( .A1(\exu.csrrs.io_csr_rdata [11] ), .A2(_08957_ ), .A3(\exu.csrrs.io_csr_rdata [10] ), .A4(\exu.csrrs.io_csr_rdata [12] ), .ZN(_10170_ ) );
OAI211_X1 _16699_ ( .A(_10169_ ), .B(_08972_ ), .C1(\exu.csrrs.io_csr_rdata [13] ), .C2(_10170_ ), .ZN(_10171_ ) );
AND2_X1 _16700_ ( .A1(fanout_net_11 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_18_A_$_MUX__A_B ), .ZN(_10172_ ) );
OAI21_X1 _16701_ ( .A(_10171_ ), .B1(_09414_ ), .B2(_10172_ ), .ZN(_10173_ ) );
NAND3_X1 _16702_ ( .A1(_10168_ ), .A2(_10173_ ), .A3(_09254_ ), .ZN(_10174_ ) );
AOI21_X1 _16703_ ( .A(fanout_net_6 ), .B1(_10167_ ), .B2(_10174_ ), .ZN(_10175_ ) );
AOI211_X1 _16704_ ( .A(_09222_ ), .B(_10165_ ), .C1(_08920_ ), .C2(_09190_ ), .ZN(_10176_ ) );
OAI21_X1 _16705_ ( .A(_09412_ ), .B1(_10175_ ), .B2(_10176_ ), .ZN(_10177_ ) );
AND2_X1 _16706_ ( .A1(_10157_ ), .A2(_10158_ ), .ZN(_10178_ ) );
OAI21_X1 _16707_ ( .A(_10177_ ), .B1(_10112_ ), .B2(_10178_ ), .ZN(_10179_ ) );
AND2_X1 _16708_ ( .A1(_10179_ ), .A2(_09250_ ), .ZN(_10180_ ) );
NOR2_X1 _16709_ ( .A1(_10178_ ), .A2(_09440_ ), .ZN(_10181_ ) );
OAI21_X1 _16710_ ( .A(_08984_ ), .B1(_10180_ ), .B2(_10181_ ), .ZN(_10182_ ) );
MUX2_X1 _16711_ ( .A(_09298_ ), .B(_08926_ ), .S(\exu.bge.io_is ), .Z(_10183_ ) );
AOI21_X1 _16712_ ( .A(_09307_ ), .B1(_10183_ ), .B2(_08984_ ), .ZN(_10184_ ) );
OAI221_X1 _16713_ ( .A(_10182_ ), .B1(_09306_ ), .B2(_10178_ ), .C1(_10165_ ), .C2(_10184_ ), .ZN(_10185_ ) );
AOI221_X4 _16714_ ( .A(_10159_ ), .B1(_09313_ ), .B2(_10166_ ), .C1(_10185_ ), .C2(_09249_ ), .ZN(_10186_ ) );
NOR2_X1 _16715_ ( .A1(_10186_ ), .A2(fanout_net_9 ), .ZN(_10187_ ) );
AND3_X1 _16716_ ( .A1(_10157_ ), .A2(_08700_ ), .A3(_10158_ ), .ZN(_10188_ ) );
AOI211_X1 _16717_ ( .A(_08702_ ), .B(_10188_ ), .C1(fanout_net_18 ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_18_A_$_MUX__A_B ), .ZN(_10189_ ) );
OAI21_X1 _16718_ ( .A(_08989_ ), .B1(_10187_ ), .B2(_10189_ ), .ZN(_10190_ ) );
NAND3_X1 _16719_ ( .A1(_09396_ ), .A2(fanout_net_8 ), .A3(\exu.csrrs.io_csr_rdata [13] ), .ZN(_10191_ ) );
NAND3_X1 _16720_ ( .A1(_10190_ ), .A2(_09042_ ), .A3(_10191_ ), .ZN(_10192_ ) );
AND2_X1 _16721_ ( .A1(_09102_ ), .A2(_09114_ ), .ZN(_10193_ ) );
NOR2_X1 _16722_ ( .A1(_10193_ ), .A2(_09112_ ), .ZN(_10194_ ) );
XNOR2_X1 _16723_ ( .A(_10194_ ), .B(_09111_ ), .ZN(\exu.addi._io_rd_T_4 [13] ) );
MUX2_X1 _16724_ ( .A(_10164_ ), .B(\exu.addi._io_rd_T_4 [13] ), .S(_09395_ ), .Z(_10195_ ) );
OR2_X1 _16725_ ( .A1(_10195_ ), .A2(_09042_ ), .ZN(_10196_ ) );
NAND3_X1 _16726_ ( .A1(_10192_ ), .A2(_09185_ ), .A3(_10196_ ), .ZN(_10197_ ) );
OAI21_X1 _16727_ ( .A(\ifu.pc [13] ), .B1(_09401_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_10198_ ) );
NAND3_X1 _16728_ ( .A1(_10197_ ), .A2(_09182_ ), .A3(_10198_ ), .ZN(_10199_ ) );
INV_X1 _16729_ ( .A(\ifu.pc [13] ), .ZN(_10200_ ) );
OAI21_X1 _16730_ ( .A(_10200_ ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10201_ ) );
NAND2_X1 _16731_ ( .A1(_10199_ ), .A2(_10201_ ), .ZN(_10202_ ) );
NOR2_X1 _16732_ ( .A1(_09246_ ), .A2(\icache.tag_reg_0 [8] ), .ZN(_10203_ ) );
AOI21_X1 _16733_ ( .A(\icache.tag_reg_1 [8] ), .B1(_09334_ ), .B2(_09336_ ), .ZN(_10204_ ) );
OR2_X1 _16734_ ( .A1(_10203_ ), .A2(_10204_ ), .ZN(_10205_ ) );
XNOR2_X1 _16735_ ( .A(_10202_ ), .B(_10205_ ), .ZN(_10206_ ) );
NAND2_X1 _16736_ ( .A1(_10155_ ), .A2(_10206_ ), .ZN(_10207_ ) );
NOR3_X1 _16737_ ( .A1(_08622_ ), .A2(_08618_ ), .A3(_08640_ ), .ZN(_10208_ ) );
XNOR2_X1 _16738_ ( .A(_10208_ ), .B(_08624_ ), .ZN(_10209_ ) );
OR2_X1 _16739_ ( .A1(_10110_ ), .A2(_10209_ ), .ZN(_10210_ ) );
INV_X1 _16740_ ( .A(\exu.auipc.io_rs1_data [10] ), .ZN(_10211_ ) );
XNOR2_X1 _16741_ ( .A(_08798_ ), .B(_10211_ ), .ZN(_10212_ ) );
AOI211_X1 _16742_ ( .A(_09255_ ), .B(_10212_ ), .C1(_09428_ ), .C2(_09191_ ), .ZN(_10213_ ) );
NOR2_X1 _16743_ ( .A1(_08957_ ), .A2(\exu.csrrs.io_csr_rdata [10] ), .ZN(_10214_ ) );
OR3_X1 _16744_ ( .A1(_10214_ ), .A2(_09214_ ), .A3(_09272_ ), .ZN(_10215_ ) );
OAI211_X1 _16745_ ( .A(_10215_ ), .B(fanout_net_11 ), .C1(\exu.addi._io_rd_T_4_$_NOT__Y_21_A_$_MUX__A_B ), .C2(_09414_ ), .ZN(_10216_ ) );
INV_X1 _16746_ ( .A(_10212_ ), .ZN(_10217_ ) );
OAI21_X1 _16747_ ( .A(_09211_ ), .B1(_10217_ ), .B2(_09036_ ), .ZN(_10218_ ) );
AOI21_X1 _16748_ ( .A(fanout_net_7 ), .B1(_10216_ ), .B2(_10218_ ), .ZN(_10219_ ) );
OAI21_X1 _16749_ ( .A(_09252_ ), .B1(_10213_ ), .B2(_10219_ ), .ZN(_10220_ ) );
OAI211_X1 _16750_ ( .A(fanout_net_6 ), .B(_10217_ ), .C1(_09944_ ), .C2(fanout_net_18 ), .ZN(_10221_ ) );
NAND4_X1 _16751_ ( .A1(_10210_ ), .A2(_09413_ ), .A3(_10220_ ), .A4(_10221_ ), .ZN(_10222_ ) );
OR2_X1 _16752_ ( .A1(_10209_ ), .A2(_08936_ ), .ZN(_10223_ ) );
OAI211_X1 _16753_ ( .A(_10223_ ), .B(\exu.bgeu.io_is ), .C1(_09437_ ), .C2(_10212_ ), .ZN(_10224_ ) );
NAND3_X1 _16754_ ( .A1(_10222_ ), .A2(_09251_ ), .A3(_10224_ ), .ZN(_10225_ ) );
NAND3_X1 _16755_ ( .A1(_09944_ ), .A2(_08923_ ), .A3(_10209_ ), .ZN(_10226_ ) );
OAI211_X1 _16756_ ( .A(\exu.bge.io_is ), .B(_10226_ ), .C1(_08925_ ), .C2(_10217_ ), .ZN(_10227_ ) );
AOI21_X1 _16757_ ( .A(\exu.bne.io_is ), .B1(_10225_ ), .B2(_10227_ ), .ZN(_10228_ ) );
AND2_X1 _16758_ ( .A1(_10209_ ), .A2(_08815_ ), .ZN(_10229_ ) );
AOI211_X1 _16759_ ( .A(_08984_ ), .B(_10229_ ), .C1(_09306_ ), .C2(_10212_ ), .ZN(_10230_ ) );
OAI21_X1 _16760_ ( .A(_09249_ ), .B1(_10228_ ), .B2(_10230_ ), .ZN(_10231_ ) );
NAND2_X1 _16761_ ( .A1(_10209_ ), .A2(_09231_ ), .ZN(_10232_ ) );
OAI211_X1 _16762_ ( .A(_10232_ ), .B(\exu.beq.io_is ), .C1(_09231_ ), .C2(_10217_ ), .ZN(_10233_ ) );
AOI21_X1 _16763_ ( .A(fanout_net_9 ), .B1(_10231_ ), .B2(_10233_ ), .ZN(_10234_ ) );
OAI21_X1 _16764_ ( .A(fanout_net_9 ), .B1(_09192_ ), .B2(\exu.addi._io_rd_T_4_$_NOT__Y_21_A_$_MUX__A_B ), .ZN(_10235_ ) );
AOI21_X1 _16765_ ( .A(_10235_ ), .B1(_10209_ ), .B2(_08700_ ), .ZN(_10236_ ) );
NOR3_X1 _16766_ ( .A1(_10234_ ), .A2(fanout_net_8 ), .A3(_10236_ ), .ZN(_10237_ ) );
AOI211_X1 _16767_ ( .A(fanout_net_10 ), .B(_10237_ ), .C1(\exu.csrrs.io_csr_rdata [10] ), .C2(_08991_ ), .ZN(_10238_ ) );
NAND3_X1 _16768_ ( .A1(fanout_net_18 ), .A2(fanout_net_10 ), .A3(\exu.addi._io_rd_T_4_$_NOT__Y_21_A_$_MUX__A_B ), .ZN(_10239_ ) );
OR3_X1 _16769_ ( .A1(_09078_ ), .A2(_09079_ ), .A3(_09086_ ), .ZN(_10240_ ) );
INV_X1 _16770_ ( .A(_09089_ ), .ZN(_10241_ ) );
AND3_X1 _16771_ ( .A1(_10240_ ), .A2(_10241_ ), .A3(_09096_ ), .ZN(_10242_ ) );
AOI21_X1 _16772_ ( .A(_10241_ ), .B1(_10240_ ), .B2(_09096_ ), .ZN(_10243_ ) );
NOR2_X1 _16773_ ( .A1(_10242_ ), .A2(_10243_ ), .ZN(\exu.addi._io_rd_T_4 [10] ) );
OAI21_X1 _16774_ ( .A(_10239_ ), .B1(\exu.addi._io_rd_T_4 [10] ), .B2(_09177_ ), .ZN(_10244_ ) );
OR3_X1 _16775_ ( .A1(_10238_ ), .A2(_09039_ ), .A3(_10244_ ), .ZN(_10245_ ) );
INV_X1 _16776_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_7_A_$_MUX__Y_B ), .ZN(_10246_ ) );
OAI21_X1 _16777_ ( .A(_10246_ ), .B1(_09401_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_10247_ ) );
NAND3_X1 _16778_ ( .A1(_10245_ ), .A2(_09181_ ), .A3(_10247_ ), .ZN(_10248_ ) );
OAI21_X1 _16779_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_7_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10249_ ) );
AND2_X1 _16780_ ( .A1(_10248_ ), .A2(_10249_ ), .ZN(_10250_ ) );
NAND2_X1 _16781_ ( .A1(_09246_ ), .A2(\icache.tag_reg_1 [5] ), .ZN(_10251_ ) );
NAND3_X1 _16782_ ( .A1(_09334_ ), .A2(\icache.tag_reg_0 [5] ), .A3(_09336_ ), .ZN(_10252_ ) );
AND3_X1 _16783_ ( .A1(_10250_ ), .A2(_10251_ ), .A3(_10252_ ), .ZN(_10253_ ) );
AOI21_X1 _16784_ ( .A(_10250_ ), .B1(_10251_ ), .B2(_10252_ ), .ZN(_10254_ ) );
OAI21_X1 _16785_ ( .A(_08617_ ), .B1(_08603_ ), .B2(_08614_ ), .ZN(_10255_ ) );
NAND2_X1 _16786_ ( .A1(_10255_ ), .A2(_08639_ ), .ZN(_10256_ ) );
XOR2_X1 _16787_ ( .A(_10256_ ), .B(_08620_ ), .Z(_10257_ ) );
OR2_X1 _16788_ ( .A1(_10257_ ), .A2(_08786_ ), .ZN(_10258_ ) );
INV_X1 _16789_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_23_A_$_MUX__A_B ), .ZN(_10259_ ) );
AND2_X1 _16790_ ( .A1(_08795_ ), .A2(_10259_ ), .ZN(_10260_ ) );
INV_X1 _16791_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_22_A_$_MUX__A_B ), .ZN(_10261_ ) );
XNOR2_X1 _16792_ ( .A(_10260_ ), .B(_10261_ ), .ZN(_10262_ ) );
INV_X1 _16793_ ( .A(_10262_ ), .ZN(_10263_ ) );
NOR2_X1 _16794_ ( .A1(_10257_ ), .A2(_09202_ ), .ZN(_10264_ ) );
INV_X1 _16795_ ( .A(_10257_ ), .ZN(_10265_ ) );
NAND3_X1 _16796_ ( .A1(_09944_ ), .A2(_08923_ ), .A3(_10265_ ), .ZN(_10266_ ) );
NOR3_X1 _16797_ ( .A1(_09428_ ), .A2(_10257_ ), .A3(_08933_ ), .ZN(_10267_ ) );
OAI21_X1 _16798_ ( .A(fanout_net_7 ), .B1(_08943_ ), .B2(_10262_ ), .ZN(_10268_ ) );
AND3_X1 _16799_ ( .A1(_08918_ ), .A2(_10257_ ), .A3(_08941_ ), .ZN(_10269_ ) );
NOR2_X1 _16800_ ( .A1(_10262_ ), .A2(_09035_ ), .ZN(_10270_ ) );
XNOR2_X1 _16801_ ( .A(_08955_ ), .B(\exu.csrrs.io_csr_rdata [9] ), .ZN(_10271_ ) );
MUX2_X1 _16802_ ( .A(_10261_ ), .B(_10271_ ), .S(_08972_ ), .Z(_10272_ ) );
MUX2_X1 _16803_ ( .A(_10270_ ), .B(_10272_ ), .S(fanout_net_11 ), .Z(_10273_ ) );
OAI22_X1 _16804_ ( .A1(_10268_ ), .A2(_10269_ ), .B1(fanout_net_7 ), .B2(_10273_ ), .ZN(_10274_ ) );
MUX2_X1 _16805_ ( .A(_10262_ ), .B(_10265_ ), .S(_08976_ ), .Z(_10275_ ) );
MUX2_X1 _16806_ ( .A(_10274_ ), .B(_10275_ ), .S(fanout_net_6 ), .Z(_10276_ ) );
AOI221_X4 _16807_ ( .A(_10267_ ), .B1(_08938_ ), .B2(_10262_ ), .C1(_10276_ ), .C2(_08931_ ), .ZN(_10277_ ) );
OAI221_X1 _16808_ ( .A(_10266_ ), .B1(_08930_ ), .B2(_10263_ ), .C1(_10277_ ), .C2(\exu.bge.io_is ), .ZN(_10278_ ) );
AOI221_X1 _16809_ ( .A(_10264_ ), .B1(_09307_ ), .B2(_10262_ ), .C1(_10278_ ), .C2(_08984_ ), .ZN(_10279_ ) );
OAI221_X1 _16810_ ( .A(_10258_ ), .B1(_08790_ ), .B2(_10263_ ), .C1(_10279_ ), .C2(\exu.beq.io_is ), .ZN(_10280_ ) );
NAND2_X1 _16811_ ( .A1(_10280_ ), .A2(_08702_ ), .ZN(_10281_ ) );
NAND2_X1 _16812_ ( .A1(fanout_net_9 ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_22_A_$_MUX__A_B ), .ZN(_10282_ ) );
MUX2_X1 _16813_ ( .A(_10282_ ), .B(_10257_ ), .S(_08700_ ), .Z(_10283_ ) );
NAND3_X1 _16814_ ( .A1(_10281_ ), .A2(_08989_ ), .A3(_10283_ ), .ZN(_10284_ ) );
OAI211_X1 _16815_ ( .A(_10284_ ), .B(_09042_ ), .C1(_08956_ ), .C2(_09456_ ), .ZN(_10285_ ) );
INV_X1 _16816_ ( .A(_09082_ ), .ZN(_10286_ ) );
NOR3_X1 _16817_ ( .A1(_09078_ ), .A2(_09079_ ), .A3(_10286_ ), .ZN(_10287_ ) );
NOR2_X1 _16818_ ( .A1(_10287_ ), .A2(_09080_ ), .ZN(_10288_ ) );
XNOR2_X1 _16819_ ( .A(_10288_ ), .B(_09085_ ), .ZN(\exu.addi._io_rd_T_4 [9] ) );
NAND2_X1 _16820_ ( .A1(\exu.addi._io_rd_T_4 [9] ), .A2(_09174_ ), .ZN(_10289_ ) );
OAI211_X1 _16821_ ( .A(_10289_ ), .B(\exu.io_in_bits_jalr ), .C1(_09396_ ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_22_A_$_MUX__A_B ), .ZN(_10290_ ) );
AND3_X1 _16822_ ( .A1(_10285_ ), .A2(_09184_ ), .A3(_10290_ ), .ZN(_10291_ ) );
INV_X1 _16823_ ( .A(_09181_ ), .ZN(\ifu._start_T ) );
NOR2_X1 _16824_ ( .A1(_09185_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_8_A_$_MUX__Y_B ), .ZN(_10292_ ) );
OR3_X4 _16825_ ( .A1(_10291_ ), .A2(\ifu._start_T ), .A3(_10292_ ), .ZN(_10293_ ) );
OAI21_X1 _16826_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_8_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10294_ ) );
NOR2_X1 _16827_ ( .A1(_09245_ ), .A2(\icache.tag_reg_0 [4] ), .ZN(_10295_ ) );
AOI21_X1 _16828_ ( .A(\icache.tag_reg_1 [4] ), .B1(_09334_ ), .B2(_09336_ ), .ZN(_10296_ ) );
NOR2_X1 _16829_ ( .A1(_10295_ ), .A2(_10296_ ), .ZN(_10297_ ) );
NAND3_X1 _16830_ ( .A1(_10293_ ), .A2(_10294_ ), .A3(_10297_ ), .ZN(_10298_ ) );
AND2_X1 _16831_ ( .A1(_10293_ ), .A2(_10294_ ), .ZN(_10299_ ) );
OR2_X1 _16832_ ( .A1(_10299_ ), .A2(_10297_ ), .ZN(_10300_ ) );
AOI211_X1 _16833_ ( .A(_10253_ ), .B(_10254_ ), .C1(_10298_ ), .C2(_10300_ ), .ZN(_10301_ ) );
NOR2_X1 _16834_ ( .A1(\exu.auipc.io_rs1_data [10] ), .A2(\exu.addi.io_imm [10] ), .ZN(_10302_ ) );
NOR3_X1 _16835_ ( .A1(_10208_ ), .A2(_08636_ ), .A3(_10302_ ), .ZN(_10303_ ) );
INV_X1 _16836_ ( .A(_08623_ ), .ZN(_10304_ ) );
OR3_X1 _16837_ ( .A1(_10303_ ), .A2(_10304_ ), .A3(_08636_ ), .ZN(_10305_ ) );
OAI21_X1 _16838_ ( .A(_10304_ ), .B1(_10303_ ), .B2(_08636_ ), .ZN(_10306_ ) );
AND3_X1 _16839_ ( .A1(_10305_ ), .A2(_08815_ ), .A3(_10306_ ), .ZN(_10307_ ) );
OAI21_X1 _16840_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_20_A_$_MUX__A_B ), .B1(_10160_ ), .B2(_10211_ ), .ZN(_10308_ ) );
INV_X1 _16841_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_20_A_$_MUX__A_B ), .ZN(_10309_ ) );
NAND3_X1 _16842_ ( .A1(_08798_ ), .A2(\exu.auipc.io_rs1_data [10] ), .A3(_10309_ ), .ZN(_10310_ ) );
NAND2_X1 _16843_ ( .A1(_10308_ ), .A2(_10310_ ), .ZN(_10311_ ) );
INV_X1 _16844_ ( .A(_10311_ ), .ZN(_10312_ ) );
NOR3_X1 _16845_ ( .A1(_09443_ ), .A2(_08984_ ), .A3(_10312_ ), .ZN(_10313_ ) );
NAND2_X1 _16846_ ( .A1(_10305_ ), .A2(_10306_ ), .ZN(_10314_ ) );
NOR2_X1 _16847_ ( .A1(_10112_ ), .A2(_10314_ ), .ZN(_10315_ ) );
NAND3_X1 _16848_ ( .A1(_09207_ ), .A2(fanout_net_7 ), .A3(_10311_ ), .ZN(_10316_ ) );
AND2_X1 _16849_ ( .A1(_09272_ ), .A2(\exu.csrrs.io_csr_rdata [11] ), .ZN(_10317_ ) );
OR2_X1 _16850_ ( .A1(_10317_ ), .A2(_09214_ ), .ZN(_10318_ ) );
INV_X1 _16851_ ( .A(_09272_ ), .ZN(_10319_ ) );
AOI21_X1 _16852_ ( .A(_10318_ ), .B1(_08960_ ), .B2(_10319_ ), .ZN(_10320_ ) );
AOI211_X1 _16853_ ( .A(_09211_ ), .B(_10320_ ), .C1(fanout_net_18 ), .C2(_10309_ ), .ZN(_10321_ ) );
AOI21_X1 _16854_ ( .A(fanout_net_11 ), .B1(_10312_ ), .B2(exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ), .ZN(_10322_ ) );
OAI21_X1 _16855_ ( .A(_09255_ ), .B1(_10321_ ), .B2(_10322_ ), .ZN(_10323_ ) );
AOI211_X1 _16856_ ( .A(\exu.bgeu.io_is ), .B(fanout_net_6 ), .C1(_10316_ ), .C2(_10323_ ), .ZN(_10324_ ) );
OAI21_X1 _16857_ ( .A(_09250_ ), .B1(_10315_ ), .B2(_10324_ ), .ZN(_10325_ ) );
OAI211_X1 _16858_ ( .A(_09412_ ), .B(fanout_net_6 ), .C1(_09944_ ), .C2(fanout_net_18 ), .ZN(_10326_ ) );
AOI21_X1 _16859_ ( .A(\exu.bge.io_is ), .B1(_10326_ ), .B2(_09299_ ), .ZN(_10327_ ) );
OAI21_X1 _16860_ ( .A(_10311_ ), .B1(_10327_ ), .B2(_08928_ ), .ZN(_10328_ ) );
OAI211_X1 _16861_ ( .A(_10325_ ), .B(_10328_ ), .C1(_09440_ ), .C2(_10314_ ), .ZN(_10329_ ) );
AOI211_X1 _16862_ ( .A(_10307_ ), .B(_10313_ ), .C1(_10329_ ), .C2(_09411_ ), .ZN(_10330_ ) );
INV_X1 _16863_ ( .A(_09231_ ), .ZN(_10331_ ) );
AOI21_X1 _16864_ ( .A(_10331_ ), .B1(_10305_ ), .B2(_10306_ ), .ZN(_10332_ ) );
OAI21_X1 _16865_ ( .A(\exu.beq.io_is ), .B1(_09231_ ), .B2(_10311_ ), .ZN(_10333_ ) );
OAI22_X1 _16866_ ( .A1(_10330_ ), .A2(\exu.beq.io_is ), .B1(_10332_ ), .B2(_10333_ ), .ZN(_10334_ ) );
AND2_X1 _16867_ ( .A1(_10334_ ), .A2(_08702_ ), .ZN(_10335_ ) );
OAI21_X1 _16868_ ( .A(fanout_net_9 ), .B1(_09395_ ), .B2(\exu.addi._io_rd_T_4_$_NOT__Y_20_A_$_MUX__A_B ), .ZN(_10336_ ) );
AOI21_X1 _16869_ ( .A(_10336_ ), .B1(_10314_ ), .B2(_09317_ ), .ZN(_10337_ ) );
NOR3_X1 _16870_ ( .A1(_10335_ ), .A2(fanout_net_8 ), .A3(_10337_ ), .ZN(_10338_ ) );
AOI211_X1 _16871_ ( .A(\exu.io_in_bits_jalr ), .B(_10338_ ), .C1(\exu.csrrs.io_csr_rdata [11] ), .C2(_08991_ ), .ZN(_10339_ ) );
NAND3_X1 _16872_ ( .A1(fanout_net_18 ), .A2(\exu.io_in_bits_jalr ), .A3(\exu.addi._io_rd_T_4_$_NOT__Y_20_A_$_MUX__A_B ), .ZN(_10340_ ) );
NOR2_X1 _16873_ ( .A1(_10243_ ), .A2(_09087_ ), .ZN(_10341_ ) );
INV_X1 _16874_ ( .A(_09092_ ), .ZN(_10342_ ) );
XNOR2_X1 _16875_ ( .A(_10341_ ), .B(_10342_ ), .ZN(_10343_ ) );
INV_X1 _16876_ ( .A(_10343_ ), .ZN(\exu.addi._io_rd_T_4 [11] ) );
OAI21_X1 _16877_ ( .A(_10340_ ), .B1(\exu.addi._io_rd_T_4 [11] ), .B2(_09177_ ), .ZN(_10344_ ) );
OR3_X1 _16878_ ( .A1(_10339_ ), .A2(_09039_ ), .A3(_10344_ ), .ZN(_10345_ ) );
OR2_X1 _16879_ ( .A1(_09185_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_6_A_$_MUX__Y_B ), .ZN(_10346_ ) );
NAND3_X1 _16880_ ( .A1(_10345_ ), .A2(_09182_ ), .A3(_10346_ ), .ZN(_10347_ ) );
OAI21_X1 _16881_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_6_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10348_ ) );
NAND2_X1 _16882_ ( .A1(_10347_ ), .A2(_10348_ ), .ZN(_10349_ ) );
NOR2_X1 _16883_ ( .A1(_09246_ ), .A2(\icache.tag_reg_0 [6] ), .ZN(_10350_ ) );
AOI21_X1 _16884_ ( .A(\icache.tag_reg_1 [6] ), .B1(_09334_ ), .B2(_09336_ ), .ZN(_10351_ ) );
OR2_X1 _16885_ ( .A1(_10350_ ), .A2(_10351_ ), .ZN(_10352_ ) );
XNOR2_X1 _16886_ ( .A(_10349_ ), .B(_10352_ ), .ZN(_10353_ ) );
XNOR2_X1 _16887_ ( .A(_09824_ ), .B(_08632_ ), .ZN(_10354_ ) );
AND2_X1 _16888_ ( .A1(_10354_ ), .A2(_08945_ ), .ZN(_10355_ ) );
XNOR2_X1 _16889_ ( .A(_10161_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_19_A_$_MUX__A_B ), .ZN(_10356_ ) );
AOI211_X1 _16890_ ( .A(_09255_ ), .B(_10355_ ), .C1(_09207_ ), .C2(_10356_ ), .ZN(_10357_ ) );
INV_X1 _16891_ ( .A(_10317_ ), .ZN(_10358_ ) );
AOI21_X1 _16892_ ( .A(_09214_ ), .B1(_10358_ ), .B2(\exu.addi._io_rd_T_4_$_NOT__Y_17_A_$_MUX__A_B_$_MUX__B_1_A_$_XOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_NOR__B_Y_$_XOR__A_B ), .ZN(_10359_ ) );
OAI21_X1 _16893_ ( .A(_10359_ ), .B1(\exu.addi._io_rd_T_4_$_NOT__Y_17_A_$_MUX__A_B_$_MUX__B_1_A_$_XOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_NOR__B_Y_$_XOR__A_B ), .B2(_10358_ ), .ZN(_10360_ ) );
OAI211_X1 _16894_ ( .A(_10360_ ), .B(fanout_net_11 ), .C1(_09190_ ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_19_A_$_MUX__A_B ), .ZN(_10361_ ) );
INV_X1 _16895_ ( .A(_10356_ ), .ZN(_10362_ ) );
OAI21_X1 _16896_ ( .A(_09288_ ), .B1(_10362_ ), .B2(_09036_ ), .ZN(_10363_ ) );
AOI21_X1 _16897_ ( .A(fanout_net_7 ), .B1(_10361_ ), .B2(_10363_ ), .ZN(_10364_ ) );
OAI21_X1 _16898_ ( .A(_09252_ ), .B1(_10357_ ), .B2(_10364_ ), .ZN(_10365_ ) );
NAND3_X1 _16899_ ( .A1(_10354_ ), .A2(_08920_ ), .A3(_08975_ ), .ZN(_10366_ ) );
OAI211_X1 _16900_ ( .A(_10366_ ), .B(fanout_net_6 ), .C1(_09220_ ), .C2(_10362_ ), .ZN(_10367_ ) );
AOI21_X1 _16901_ ( .A(\exu.bgeu.io_is ), .B1(_10365_ ), .B2(_10367_ ), .ZN(_10368_ ) );
AND2_X1 _16902_ ( .A1(_10354_ ), .A2(_08935_ ), .ZN(_10369_ ) );
AOI211_X1 _16903_ ( .A(_09413_ ), .B(_10369_ ), .C1(_09297_ ), .C2(_10356_ ), .ZN(_10370_ ) );
OAI21_X1 _16904_ ( .A(_09250_ ), .B1(_10368_ ), .B2(_10370_ ), .ZN(_10371_ ) );
NAND3_X1 _16905_ ( .A1(_10354_ ), .A2(_09944_ ), .A3(_08923_ ), .ZN(_10372_ ) );
OAI211_X1 _16906_ ( .A(\exu.bge.io_is ), .B(_10372_ ), .C1(_08925_ ), .C2(_10362_ ), .ZN(_10373_ ) );
AOI21_X1 _16907_ ( .A(\exu.bne.io_is ), .B1(_10371_ ), .B2(_10373_ ), .ZN(_10374_ ) );
OAI22_X1 _16908_ ( .A1(_10354_ ), .A2(_09202_ ), .B1(_09309_ ), .B2(_10356_ ), .ZN(_10375_ ) );
OAI21_X1 _16909_ ( .A(_08788_ ), .B1(_10374_ ), .B2(_10375_ ), .ZN(_10376_ ) );
NAND2_X1 _16910_ ( .A1(_10354_ ), .A2(_09231_ ), .ZN(_10377_ ) );
OAI211_X1 _16911_ ( .A(_10377_ ), .B(\exu.beq.io_is ), .C1(_09231_ ), .C2(_10362_ ), .ZN(_10378_ ) );
AOI21_X1 _16912_ ( .A(fanout_net_9 ), .B1(_10376_ ), .B2(_10378_ ), .ZN(_10379_ ) );
OAI21_X1 _16913_ ( .A(\exu.io_in_bits_jal ), .B1(_09192_ ), .B2(\exu.addi._io_rd_T_4_$_NOT__Y_19_A_$_MUX__A_B ), .ZN(_10380_ ) );
AOI21_X1 _16914_ ( .A(_10380_ ), .B1(_10354_ ), .B2(_08700_ ), .ZN(_10381_ ) );
NOR3_X1 _16915_ ( .A1(_10379_ ), .A2(fanout_net_8 ), .A3(_10381_ ), .ZN(_10382_ ) );
AOI211_X1 _16916_ ( .A(\exu.io_in_bits_jalr ), .B(_10382_ ), .C1(\exu.csrrs.io_csr_rdata [12] ), .C2(_08991_ ), .ZN(_10383_ ) );
NAND3_X1 _16917_ ( .A1(fanout_net_18 ), .A2(\exu.io_in_bits_jalr ), .A3(\exu.addi._io_rd_T_4_$_NOT__Y_19_A_$_MUX__A_B ), .ZN(_10384_ ) );
XOR2_X1 _16918_ ( .A(_09102_ ), .B(_09114_ ), .Z(\exu.addi._io_rd_T_4 [12] ) );
OAI21_X1 _16919_ ( .A(_10384_ ), .B1(\exu.addi._io_rd_T_4 [12] ), .B2(_09176_ ), .ZN(_10385_ ) );
OR3_X1 _16920_ ( .A1(_10383_ ), .A2(_09039_ ), .A3(_10385_ ), .ZN(_10386_ ) );
OR2_X1 _16921_ ( .A1(_09185_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_5_A_$_MUX__Y_B ), .ZN(_10387_ ) );
NAND3_X1 _16922_ ( .A1(_10386_ ), .A2(_09181_ ), .A3(_10387_ ), .ZN(_10388_ ) );
OAI21_X1 _16923_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_5_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10389_ ) );
AND2_X1 _16924_ ( .A1(_10388_ ), .A2(_10389_ ), .ZN(_10390_ ) );
MUX2_X1 _16925_ ( .A(\icache.tag_reg_0 [7] ), .B(\icache.tag_reg_1 [7] ), .S(_09245_ ), .Z(_10391_ ) );
XNOR2_X1 _16926_ ( .A(_10390_ ), .B(_10391_ ), .ZN(_10392_ ) );
NAND3_X1 _16927_ ( .A1(_09192_ ), .A2(fanout_net_8 ), .A3(\exu.csrrs.io_csr_rdata [6] ), .ZN(_10393_ ) );
AND2_X1 _16928_ ( .A1(_08598_ ), .A2(_08585_ ), .ZN(_10394_ ) );
OAI21_X1 _16929_ ( .A(_08611_ ), .B1(_10394_ ), .B2(_08609_ ), .ZN(_10395_ ) );
XNOR2_X1 _16930_ ( .A(_10395_ ), .B(_08600_ ), .ZN(_10396_ ) );
OR3_X1 _16931_ ( .A1(_09428_ ), .A2(_08933_ ), .A3(_10396_ ), .ZN(_10397_ ) );
XNOR2_X1 _16932_ ( .A(_08793_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_25_A_$_MUX__A_B ), .ZN(_10398_ ) );
OAI211_X1 _16933_ ( .A(_10397_ ), .B(\exu.bgeu.io_is ), .C1(_09437_ ), .C2(_10398_ ), .ZN(_10399_ ) );
INV_X1 _16934_ ( .A(_10398_ ), .ZN(_10400_ ) );
OAI211_X1 _16935_ ( .A(fanout_net_6 ), .B(_10400_ ), .C1(_08921_ ), .C2(fanout_net_18 ), .ZN(_10401_ ) );
OAI211_X1 _16936_ ( .A(_10401_ ), .B(_09412_ ), .C1(_09432_ ), .C2(_10396_ ), .ZN(_10402_ ) );
NAND4_X1 _16937_ ( .A1(_08866_ ), .A2(_08917_ ), .A3(_08941_ ), .A4(_10396_ ), .ZN(_10403_ ) );
OAI211_X1 _16938_ ( .A(fanout_net_7 ), .B(_10403_ ), .C1(_08945_ ), .C2(_10400_ ), .ZN(_10404_ ) );
NAND3_X1 _16939_ ( .A1(fanout_net_18 ), .A2(fanout_net_11 ), .A3(\exu.addi._io_rd_T_4_$_NOT__Y_25_A_$_MUX__A_B ), .ZN(_10405_ ) );
AND2_X1 _16940_ ( .A1(_08951_ ), .A2(\exu.csrrs.io_csr_rdata [5] ), .ZN(_10406_ ) );
XNOR2_X1 _16941_ ( .A(_10406_ ), .B(\ifu.io_out_bits_pc_$_NOT__Y_11_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ), .ZN(_10407_ ) );
AND2_X1 _16942_ ( .A1(_10398_ ), .A2(exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ), .ZN(_10408_ ) );
OAI221_X1 _16943_ ( .A(_10405_ ), .B1(_09271_ ), .B2(_10407_ ), .C1(_10408_ ), .C2(\exu.io_in_bits_mret ), .ZN(_10409_ ) );
NAND2_X1 _16944_ ( .A1(_10409_ ), .A2(_09254_ ), .ZN(_10410_ ) );
AOI21_X1 _16945_ ( .A(fanout_net_6 ), .B1(_10404_ ), .B2(_10410_ ), .ZN(_10411_ ) );
OAI211_X1 _16946_ ( .A(_09250_ ), .B(_10399_ ), .C1(_10402_ ), .C2(_10411_ ), .ZN(_10412_ ) );
NAND3_X1 _16947_ ( .A1(_09944_ ), .A2(_08923_ ), .A3(_10396_ ), .ZN(_10413_ ) );
OAI211_X1 _16948_ ( .A(\exu.bge.io_is ), .B(_10413_ ), .C1(_08925_ ), .C2(_10400_ ), .ZN(_10414_ ) );
AOI21_X1 _16949_ ( .A(\exu.bne.io_is ), .B1(_10412_ ), .B2(_10414_ ), .ZN(_10415_ ) );
OAI22_X1 _16950_ ( .A1(_10396_ ), .A2(_09202_ ), .B1(_09309_ ), .B2(_10398_ ), .ZN(_10416_ ) );
OAI21_X1 _16951_ ( .A(_08788_ ), .B1(_10415_ ), .B2(_10416_ ), .ZN(_10417_ ) );
INV_X1 _16952_ ( .A(_10396_ ), .ZN(_10418_ ) );
AOI22_X1 _16953_ ( .A1(_10418_ ), .A2(_08784_ ), .B1(_09313_ ), .B2(_10400_ ), .ZN(_10419_ ) );
AOI21_X1 _16954_ ( .A(\exu.io_in_bits_jal ), .B1(_10417_ ), .B2(_10419_ ), .ZN(_10420_ ) );
INV_X1 _16955_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_25_A_$_MUX__A_B ), .ZN(_10421_ ) );
MUX2_X1 _16956_ ( .A(_10421_ ), .B(_10396_ ), .S(_08700_ ), .Z(_10422_ ) );
OAI21_X1 _16957_ ( .A(_08989_ ), .B1(_10422_ ), .B2(_08698_ ), .ZN(_10423_ ) );
OAI211_X1 _16958_ ( .A(_09042_ ), .B(_10393_ ), .C1(_10420_ ), .C2(_10423_ ), .ZN(_10424_ ) );
NOR2_X1 _16959_ ( .A1(_09074_ ), .A2(_09075_ ), .ZN(_10425_ ) );
XNOR2_X1 _16960_ ( .A(_09073_ ), .B(_10425_ ), .ZN(\exu.addi._io_rd_T_4 [6] ) );
NAND2_X1 _16961_ ( .A1(\exu.addi._io_rd_T_4 [6] ), .A2(_09174_ ), .ZN(_10426_ ) );
OAI211_X1 _16962_ ( .A(_10426_ ), .B(\exu.io_in_bits_jalr ), .C1(_09192_ ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_25_A_$_MUX__A_B ), .ZN(_10427_ ) );
NAND3_X1 _16963_ ( .A1(_10424_ ), .A2(_09184_ ), .A3(_10427_ ), .ZN(_10428_ ) );
INV_X1 _16964_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_11_A_$_MUX__Y_B ), .ZN(_10429_ ) );
OAI21_X1 _16965_ ( .A(_10429_ ), .B1(_09037_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_10430_ ) );
NAND3_X1 _16966_ ( .A1(_10428_ ), .A2(_09181_ ), .A3(_10430_ ), .ZN(_10431_ ) );
OAI21_X1 _16967_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_11_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10432_ ) );
AND2_X1 _16968_ ( .A1(_10431_ ), .A2(_10432_ ), .ZN(_10433_ ) );
NOR2_X1 _16969_ ( .A1(_09245_ ), .A2(\icache.tag_reg_0 [1] ), .ZN(_10434_ ) );
AOI21_X1 _16970_ ( .A(\icache.tag_reg_1 [1] ), .B1(_09334_ ), .B2(_09336_ ), .ZN(_10435_ ) );
OAI21_X1 _16971_ ( .A(_10433_ ), .B1(_10434_ ), .B2(_10435_ ), .ZN(_10436_ ) );
INV_X1 _16972_ ( .A(_10394_ ), .ZN(_10437_ ) );
NAND2_X1 _16973_ ( .A1(_10437_ ), .A2(_08606_ ), .ZN(_10438_ ) );
XOR2_X1 _16974_ ( .A(_10438_ ), .B(_08602_ ), .Z(_10439_ ) );
OR2_X1 _16975_ ( .A1(_10439_ ), .A2(_08785_ ), .ZN(_10440_ ) );
XNOR2_X1 _16976_ ( .A(_09195_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_26_A_$_MUX__A_B ), .ZN(_10441_ ) );
INV_X1 _16977_ ( .A(_10441_ ), .ZN(_10442_ ) );
NOR2_X1 _16978_ ( .A1(_10439_ ), .A2(_09202_ ), .ZN(_10443_ ) );
INV_X1 _16979_ ( .A(_10439_ ), .ZN(_10444_ ) );
NAND3_X1 _16980_ ( .A1(_08921_ ), .A2(_08923_ ), .A3(_10444_ ), .ZN(_10445_ ) );
NOR3_X1 _16981_ ( .A1(_08918_ ), .A2(_08933_ ), .A3(_10439_ ), .ZN(_10446_ ) );
NAND3_X1 _16982_ ( .A1(_08920_ ), .A2(_08975_ ), .A3(_10439_ ), .ZN(_10447_ ) );
OAI211_X1 _16983_ ( .A(fanout_net_6 ), .B(_10447_ ), .C1(_08976_ ), .C2(_10441_ ), .ZN(_10448_ ) );
NOR2_X1 _16984_ ( .A1(_08951_ ), .A2(\exu.csrrs.io_csr_rdata [5] ), .ZN(_10449_ ) );
OR3_X1 _16985_ ( .A1(_10406_ ), .A2(_10449_ ), .A3(_09214_ ), .ZN(_10450_ ) );
OAI211_X1 _16986_ ( .A(_10450_ ), .B(\exu.io_in_bits_mret ), .C1(_08978_ ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_26_A_$_MUX__A_B ), .ZN(_10451_ ) );
OAI21_X1 _16987_ ( .A(_08949_ ), .B1(_10441_ ), .B2(_09035_ ), .ZN(_10452_ ) );
AOI21_X1 _16988_ ( .A(fanout_net_7 ), .B1(_10451_ ), .B2(_10452_ ), .ZN(_10453_ ) );
MUX2_X1 _16989_ ( .A(_10441_ ), .B(_10444_ ), .S(_08943_ ), .Z(_10454_ ) );
AOI21_X1 _16990_ ( .A(_10453_ ), .B1(_10454_ ), .B2(fanout_net_7 ), .ZN(_10455_ ) );
OAI21_X1 _16991_ ( .A(_10448_ ), .B1(_10455_ ), .B2(fanout_net_6 ), .ZN(_10456_ ) );
AOI221_X4 _16992_ ( .A(_10446_ ), .B1(_08938_ ), .B2(_10441_ ), .C1(_10456_ ), .C2(_08931_ ), .ZN(_10457_ ) );
OAI221_X1 _16993_ ( .A(_10445_ ), .B1(_08929_ ), .B2(_10442_ ), .C1(_10457_ ), .C2(\exu.bge.io_is ), .ZN(_10458_ ) );
AOI221_X4 _16994_ ( .A(_10443_ ), .B1(_09307_ ), .B2(_10441_ ), .C1(_10458_ ), .C2(_08812_ ), .ZN(_10459_ ) );
OAI221_X1 _16995_ ( .A(_10440_ ), .B1(_08790_ ), .B2(_10442_ ), .C1(_10459_ ), .C2(\exu.beq.io_is ), .ZN(_10460_ ) );
NAND2_X1 _16996_ ( .A1(_10460_ ), .A2(_08702_ ), .ZN(_10461_ ) );
NAND2_X1 _16997_ ( .A1(\exu.io_in_bits_jal ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_26_A_$_MUX__A_B ), .ZN(_10462_ ) );
MUX2_X1 _16998_ ( .A(_10462_ ), .B(_10439_ ), .S(_08700_ ), .Z(_10463_ ) );
NAND3_X1 _16999_ ( .A1(_10461_ ), .A2(_08989_ ), .A3(_10463_ ), .ZN(_10464_ ) );
NAND3_X1 _17000_ ( .A1(_09192_ ), .A2(fanout_net_8 ), .A3(\exu.csrrs.io_csr_rdata [5] ), .ZN(_10465_ ) );
NAND3_X1 _17001_ ( .A1(_10464_ ), .A2(_09042_ ), .A3(_10465_ ), .ZN(_10466_ ) );
AND3_X1 _17002_ ( .A1(_09064_ ), .A2(_09050_ ), .A3(_09066_ ), .ZN(_10467_ ) );
NOR2_X1 _17003_ ( .A1(_10467_ ), .A2(_09071_ ), .ZN(_10468_ ) );
XNOR2_X1 _17004_ ( .A(_10468_ ), .B(_09069_ ), .ZN(\exu.addi._io_rd_T_4 [5] ) );
NAND2_X1 _17005_ ( .A1(\exu.addi._io_rd_T_4 [5] ), .A2(_09174_ ), .ZN(_10469_ ) );
OAI211_X1 _17006_ ( .A(_10469_ ), .B(\exu.io_in_bits_jalr ), .C1(_09395_ ), .C2(\exu.addi._io_rd_T_4_$_NOT__Y_26_A_$_MUX__A_B ), .ZN(_10470_ ) );
AND3_X1 _17007_ ( .A1(_10466_ ), .A2(_09184_ ), .A3(_10470_ ), .ZN(_10471_ ) );
NOR2_X1 _17008_ ( .A1(_09184_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_12_A_$_MUX__Y_B ), .ZN(_10472_ ) );
OR3_X1 _17009_ ( .A1(_10471_ ), .A2(\ifu._start_T ), .A3(_10472_ ), .ZN(_10473_ ) );
OAI21_X1 _17010_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_12_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10474_ ) );
AND2_X1 _17011_ ( .A1(_10473_ ), .A2(_10474_ ), .ZN(_10475_ ) );
MUX2_X1 _17012_ ( .A(\icache.tag_reg_0 [0] ), .B(\icache.tag_reg_1 [0] ), .S(_09245_ ), .Z(_10476_ ) );
XNOR2_X1 _17013_ ( .A(_10475_ ), .B(_10476_ ), .ZN(_10477_ ) );
OR3_X1 _17014_ ( .A1(_10434_ ), .A2(_10433_ ), .A3(_10435_ ), .ZN(_10478_ ) );
NAND2_X1 _17015_ ( .A1(_08793_ ), .A2(_10421_ ), .ZN(_10479_ ) );
XNOR2_X1 _17016_ ( .A(_10479_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_24_A_$_MUX__A_B ), .ZN(_10480_ ) );
INV_X1 _17017_ ( .A(_10480_ ), .ZN(_10481_ ) );
NAND4_X1 _17018_ ( .A1(_08977_ ), .A2(_08922_ ), .A3(_08931_ ), .A4(\exu.blt.io_is ), .ZN(_10482_ ) );
AOI21_X1 _17019_ ( .A(_10481_ ), .B1(_08929_ ), .B2(_10482_ ), .ZN(_10483_ ) );
NOR2_X1 _17020_ ( .A1(\exu.auipc.io_rs1_data [6] ), .A2(\exu.addi.io_imm [6] ), .ZN(_10484_ ) );
NOR3_X1 _17021_ ( .A1(_10395_ ), .A2(_08604_ ), .A3(_10484_ ), .ZN(_10485_ ) );
NOR2_X1 _17022_ ( .A1(_10485_ ), .A2(_08604_ ), .ZN(_10486_ ) );
XNOR2_X1 _17023_ ( .A(_10486_ ), .B(_08599_ ), .ZN(_10487_ ) );
INV_X1 _17024_ ( .A(_10487_ ), .ZN(_10488_ ) );
AOI21_X1 _17025_ ( .A(_10483_ ), .B1(_08925_ ), .B2(_10488_ ), .ZN(_10489_ ) );
AND3_X1 _17026_ ( .A1(_10487_ ), .A2(_09428_ ), .A3(_08941_ ), .ZN(_10490_ ) );
AOI211_X1 _17027_ ( .A(_09254_ ), .B(_10490_ ), .C1(_09207_ ), .C2(_10481_ ), .ZN(_10491_ ) );
XNOR2_X1 _17028_ ( .A(_08952_ ), .B(\exu.csrrs.io_csr_rdata [7] ), .ZN(_10492_ ) );
NAND2_X1 _17029_ ( .A1(_10492_ ), .A2(_08972_ ), .ZN(_10493_ ) );
OAI211_X1 _17030_ ( .A(_10493_ ), .B(\exu.io_in_bits_mret ), .C1(\exu.addi._io_rd_T_4_$_NOT__Y_24_A_$_MUX__A_B ), .C2(_09414_ ), .ZN(_10494_ ) );
OAI21_X1 _17031_ ( .A(_09211_ ), .B1(_10480_ ), .B2(_09035_ ), .ZN(_10495_ ) );
AOI21_X1 _17032_ ( .A(fanout_net_7 ), .B1(_10494_ ), .B2(_10495_ ), .ZN(_10496_ ) );
OAI21_X1 _17033_ ( .A(_09222_ ), .B1(_10491_ ), .B2(_10496_ ), .ZN(_10497_ ) );
NAND3_X1 _17034_ ( .A1(_08920_ ), .A2(_08975_ ), .A3(_10488_ ), .ZN(_10498_ ) );
AOI21_X1 _17035_ ( .A(\exu.bgeu.io_is ), .B1(_10497_ ), .B2(_10498_ ), .ZN(_10499_ ) );
NAND2_X1 _17036_ ( .A1(_10488_ ), .A2(_08935_ ), .ZN(_10500_ ) );
OAI21_X1 _17037_ ( .A(_10500_ ), .B1(_09299_ ), .B2(_10481_ ), .ZN(_10501_ ) );
OAI21_X1 _17038_ ( .A(_09250_ ), .B1(_10499_ ), .B2(_10501_ ), .ZN(_10502_ ) );
AOI21_X1 _17039_ ( .A(\exu.bne.io_is ), .B1(_10489_ ), .B2(_10502_ ), .ZN(_10503_ ) );
OAI22_X1 _17040_ ( .A1(_10487_ ), .A2(_09202_ ), .B1(_09308_ ), .B2(_10481_ ), .ZN(_10504_ ) );
OAI21_X1 _17041_ ( .A(_08788_ ), .B1(_10503_ ), .B2(_10504_ ), .ZN(_10505_ ) );
AOI22_X1 _17042_ ( .A1(_10488_ ), .A2(_08784_ ), .B1(_09313_ ), .B2(_10480_ ), .ZN(_10506_ ) );
AOI21_X1 _17043_ ( .A(\exu.io_in_bits_jal ), .B1(_10505_ ), .B2(_10506_ ), .ZN(_10507_ ) );
AND2_X1 _17044_ ( .A1(\exu.io_in_bits_jal ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_24_A_$_MUX__A_B ), .ZN(_10508_ ) );
MUX2_X1 _17045_ ( .A(_10508_ ), .B(_10488_ ), .S(_08700_ ), .Z(_10509_ ) );
NOR3_X1 _17046_ ( .A1(_10507_ ), .A2(fanout_net_8 ), .A3(_10509_ ), .ZN(_10510_ ) );
AOI211_X1 _17047_ ( .A(\exu.io_in_bits_jalr ), .B(_10510_ ), .C1(\exu.csrrs.io_csr_rdata [7] ), .C2(_08990_ ), .ZN(_10511_ ) );
OAI21_X1 _17048_ ( .A(\exu.io_in_bits_jalr ), .B1(_09395_ ), .B2(\exu.addi._io_rd_T_4_$_NOT__Y_24_A_$_MUX__A_B ), .ZN(_10512_ ) );
NOR2_X1 _17049_ ( .A1(_09076_ ), .A2(_09074_ ), .ZN(_10513_ ) );
NOR2_X1 _17050_ ( .A1(_09077_ ), .A2(_09079_ ), .ZN(_10514_ ) );
XNOR2_X1 _17051_ ( .A(_10513_ ), .B(_10514_ ), .ZN(\exu.addi._io_rd_T_4 [7] ) );
AOI21_X1 _17052_ ( .A(_10512_ ), .B1(\exu.addi._io_rd_T_4 [7] ), .B2(_09174_ ), .ZN(_10515_ ) );
OR3_X1 _17053_ ( .A1(_10511_ ), .A2(_09039_ ), .A3(_10515_ ), .ZN(_10516_ ) );
OR2_X1 _17054_ ( .A1(_09184_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_10_A_$_MUX__Y_B ), .ZN(_10517_ ) );
NAND3_X1 _17055_ ( .A1(_10516_ ), .A2(_09181_ ), .A3(_10517_ ), .ZN(_10518_ ) );
OAI21_X1 _17056_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_10_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10519_ ) );
AND2_X1 _17057_ ( .A1(_10518_ ), .A2(_10519_ ), .ZN(_10520_ ) );
NAND2_X1 _17058_ ( .A1(_09245_ ), .A2(\icache.tag_reg_1 [2] ), .ZN(_10521_ ) );
NAND3_X1 _17059_ ( .A1(_09334_ ), .A2(\icache.tag_reg_0 [2] ), .A3(_09336_ ), .ZN(_10522_ ) );
AND2_X1 _17060_ ( .A1(_10521_ ), .A2(_10522_ ), .ZN(_10523_ ) );
XNOR2_X1 _17061_ ( .A(_10520_ ), .B(_10523_ ), .ZN(_10524_ ) );
XNOR2_X1 _17062_ ( .A(_08795_ ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_23_A_$_MUX__A_B ), .ZN(_10525_ ) );
AOI21_X1 _17063_ ( .A(_09222_ ), .B1(_08977_ ), .B2(_10525_ ), .ZN(_10526_ ) );
XNOR2_X1 _17064_ ( .A(_08615_ ), .B(_08617_ ), .ZN(_10527_ ) );
INV_X1 _17065_ ( .A(_10527_ ), .ZN(_10528_ ) );
OAI21_X1 _17066_ ( .A(_10526_ ), .B1(_09798_ ), .B2(_10528_ ), .ZN(_10529_ ) );
INV_X1 _17067_ ( .A(_10525_ ), .ZN(_10530_ ) );
AOI21_X1 _17068_ ( .A(_10530_ ), .B1(_09428_ ), .B2(_08941_ ), .ZN(_10531_ ) );
AND4_X1 _17069_ ( .A1(_09190_ ), .A2(_08866_ ), .A3(_08917_ ), .A4(_10527_ ), .ZN(_10532_ ) );
OAI21_X1 _17070_ ( .A(\exu.bltu.io_is ), .B1(_10531_ ), .B2(_10532_ ), .ZN(_10533_ ) );
XNOR2_X1 _17071_ ( .A(_08954_ ), .B(\ifu.io_out_bits_pc_$_NOT__Y_9_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ), .ZN(_10534_ ) );
AND2_X1 _17072_ ( .A1(_10525_ ), .A2(_09209_ ), .ZN(_10535_ ) );
AOI21_X1 _17073_ ( .A(_09211_ ), .B1(fanout_net_18 ), .B2(\exu.addi._io_rd_T_4_$_NOT__Y_23_A_$_MUX__A_B ), .ZN(_10536_ ) );
OAI221_X1 _17074_ ( .A(_09254_ ), .B1(_09271_ ), .B2(_10534_ ), .C1(_10535_ ), .C2(_10536_ ), .ZN(_10537_ ) );
NAND3_X1 _17075_ ( .A1(_10533_ ), .A2(_09222_ ), .A3(_10537_ ), .ZN(_10538_ ) );
NAND3_X1 _17076_ ( .A1(_10529_ ), .A2(_09412_ ), .A3(_10538_ ), .ZN(_10539_ ) );
OR3_X1 _17077_ ( .A1(_09428_ ), .A2(_08933_ ), .A3(_10527_ ), .ZN(_10540_ ) );
OAI211_X1 _17078_ ( .A(_10540_ ), .B(\exu.bgeu.io_is ), .C1(_09437_ ), .C2(_10525_ ), .ZN(_10541_ ) );
NAND3_X1 _17079_ ( .A1(_10539_ ), .A2(_09250_ ), .A3(_10541_ ), .ZN(_10542_ ) );
NAND3_X1 _17080_ ( .A1(_09944_ ), .A2(_08923_ ), .A3(_10527_ ), .ZN(_10543_ ) );
OAI211_X1 _17081_ ( .A(\exu.bge.io_is ), .B(_10543_ ), .C1(_08925_ ), .C2(_10530_ ), .ZN(_10544_ ) );
AOI21_X1 _17082_ ( .A(\exu.bne.io_is ), .B1(_10542_ ), .B2(_10544_ ), .ZN(_10545_ ) );
OAI22_X1 _17083_ ( .A1(_10527_ ), .A2(_09202_ ), .B1(_09309_ ), .B2(_10525_ ), .ZN(_10546_ ) );
OAI21_X1 _17084_ ( .A(_08788_ ), .B1(_10545_ ), .B2(_10546_ ), .ZN(_10547_ ) );
AOI22_X1 _17085_ ( .A1(_10528_ ), .A2(_08784_ ), .B1(_09313_ ), .B2(_10530_ ), .ZN(_10548_ ) );
AOI21_X1 _17086_ ( .A(\exu.io_in_bits_jal ), .B1(_10547_ ), .B2(_10548_ ), .ZN(_10549_ ) );
MUX2_X1 _17087_ ( .A(_10259_ ), .B(_10527_ ), .S(_08700_ ), .Z(_10550_ ) );
NOR2_X1 _17088_ ( .A1(_10550_ ), .A2(_08698_ ), .ZN(_10551_ ) );
NOR3_X1 _17089_ ( .A1(_10549_ ), .A2(fanout_net_8 ), .A3(_10551_ ), .ZN(_10552_ ) );
AOI211_X1 _17090_ ( .A(\exu.io_in_bits_jalr ), .B(_10552_ ), .C1(\exu.csrrs.io_csr_rdata [8] ), .C2(_08990_ ), .ZN(_10553_ ) );
NOR2_X1 _17091_ ( .A1(_09078_ ), .A2(_09079_ ), .ZN(_10554_ ) );
XNOR2_X1 _17092_ ( .A(_10554_ ), .B(_10286_ ), .ZN(\exu.addi._io_rd_T_4 [8] ) );
AND2_X1 _17093_ ( .A1(\exu.addi._io_rd_T_4 [8] ), .A2(_09174_ ), .ZN(_10555_ ) );
AOI211_X1 _17094_ ( .A(_09042_ ), .B(_10555_ ), .C1(fanout_net_19 ), .C2(_10259_ ), .ZN(_10556_ ) );
OR3_X1 _17095_ ( .A1(_10553_ ), .A2(_09039_ ), .A3(_10556_ ), .ZN(_10557_ ) );
OR2_X1 _17096_ ( .A1(_09184_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_9_A_$_MUX__Y_B ), .ZN(_10558_ ) );
NAND3_X1 _17097_ ( .A1(_10557_ ), .A2(_09181_ ), .A3(_10558_ ), .ZN(_10559_ ) );
OAI21_X1 _17098_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_9_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_10560_ ) );
AND2_X1 _17099_ ( .A1(_10559_ ), .A2(_10560_ ), .ZN(_10561_ ) );
NAND2_X1 _17100_ ( .A1(_09245_ ), .A2(\icache.tag_reg_1 [3] ), .ZN(_10562_ ) );
NAND3_X1 _17101_ ( .A1(_09334_ ), .A2(\icache.tag_reg_0 [3] ), .A3(_09336_ ), .ZN(_10563_ ) );
AND3_X1 _17102_ ( .A1(_10561_ ), .A2(_10562_ ), .A3(_10563_ ), .ZN(_10564_ ) );
AOI21_X1 _17103_ ( .A(_10561_ ), .B1(_10562_ ), .B2(_10563_ ), .ZN(_10565_ ) );
NOR3_X1 _17104_ ( .A1(_10524_ ), .A2(_10564_ ), .A3(_10565_ ), .ZN(_10566_ ) );
AND4_X1 _17105_ ( .A1(_10436_ ), .A2(_10477_ ), .A3(_10478_ ), .A4(_10566_ ), .ZN(_10567_ ) );
NAND4_X1 _17106_ ( .A1(_10301_ ), .A2(_10353_ ), .A3(_10392_ ), .A4(_10567_ ), .ZN(_10568_ ) );
NOR4_X2 _17107_ ( .A1(_09921_ ), .A2(_10109_ ), .A3(_10207_ ), .A4(_10568_ ), .ZN(_10569_ ) );
INV_X1 _17108_ ( .A(_10569_ ), .ZN(_10570_ ) );
NOR3_X1 _17109_ ( .A1(_09656_ ), .A2(_09823_ ), .A3(_10570_ ), .ZN(_10571_ ) );
AND4_X1 _17110_ ( .A1(\exu.io_in_valid ), .A2(_09013_ ), .A3(_09034_ ), .A4(\exu.io_in_bits_fencei ), .ZN(_10572_ ) );
NOR2_X1 _17111_ ( .A1(_09775_ ), .A2(_10572_ ), .ZN(_10573_ ) );
INV_X1 _17112_ ( .A(\idu.rs_reg ), .ZN(_10574_ ) );
NOR2_X1 _17113_ ( .A1(_10574_ ), .A2(\idu.io_in_valid ), .ZN(_10575_ ) );
BUF_X4 _17114_ ( .A(_10575_ ), .Z(_10576_ ) );
INV_X1 _17115_ ( .A(\idu.io_in_bits_inst [27] ), .ZN(_10577_ ) );
NOR2_X1 _17116_ ( .A1(_10576_ ), .A2(_10577_ ), .ZN(_10578_ ) );
INV_X1 _17117_ ( .A(\idu.io_in_bits_inst [26] ), .ZN(_10579_ ) );
NOR2_X1 _17118_ ( .A1(_10576_ ), .A2(_10579_ ), .ZN(_10580_ ) );
NOR2_X1 _17119_ ( .A1(_10578_ ), .A2(_10580_ ), .ZN(_10581_ ) );
INV_X1 _17120_ ( .A(\idu.io_in_bits_inst [25] ), .ZN(_10582_ ) );
NOR2_X1 _17121_ ( .A1(_10576_ ), .A2(_10582_ ), .ZN(\idu.funct7 [0] ) );
INV_X1 _17122_ ( .A(\idu.funct7 [0] ), .ZN(_10583_ ) );
AND2_X1 _17123_ ( .A1(_10581_ ), .A2(_10583_ ), .ZN(_10584_ ) );
BUF_X4 _17124_ ( .A(_10576_ ), .Z(_10585_ ) );
INV_X1 _17125_ ( .A(\idu.io_in_bits_inst [31] ), .ZN(_10586_ ) );
NOR2_X1 _17126_ ( .A1(_10585_ ), .A2(_10586_ ), .ZN(_10587_ ) );
INV_X1 _17127_ ( .A(_10587_ ), .ZN(_10588_ ) );
INV_X1 _17128_ ( .A(\idu.io_in_bits_inst [30] ), .ZN(_10589_ ) );
NOR2_X1 _17129_ ( .A1(_10585_ ), .A2(_10589_ ), .ZN(_10590_ ) );
INV_X1 _17130_ ( .A(_10590_ ), .ZN(_10591_ ) );
AND3_X1 _17131_ ( .A1(_10584_ ), .A2(_10588_ ), .A3(_10591_ ), .ZN(_10592_ ) );
INV_X1 _17132_ ( .A(\idu.io_in_bits_inst [16] ), .ZN(_10593_ ) );
NOR2_X1 _17133_ ( .A1(_10585_ ), .A2(_10593_ ), .ZN(_10594_ ) );
INV_X1 _17134_ ( .A(_10594_ ), .ZN(_10595_ ) );
INV_X1 _17135_ ( .A(\idu.io_in_bits_inst [17] ), .ZN(_10596_ ) );
NOR2_X1 _17136_ ( .A1(_10576_ ), .A2(_10596_ ), .ZN(_10597_ ) );
INV_X1 _17137_ ( .A(_10597_ ), .ZN(_10598_ ) );
INV_X1 _17138_ ( .A(\idu.io_in_bits_inst [18] ), .ZN(_10599_ ) );
NOR2_X1 _17139_ ( .A1(_10576_ ), .A2(_10599_ ), .ZN(_10600_ ) );
INV_X1 _17140_ ( .A(_10600_ ), .ZN(_10601_ ) );
NAND3_X1 _17141_ ( .A1(_10595_ ), .A2(_10598_ ), .A3(_10601_ ), .ZN(_10602_ ) );
BUF_X4 _17142_ ( .A(_10585_ ), .Z(_10603_ ) );
INV_X1 _17143_ ( .A(\idu.io_in_bits_inst [19] ), .ZN(_10604_ ) );
NOR2_X1 _17144_ ( .A1(_10603_ ), .A2(_10604_ ), .ZN(_10605_ ) );
NOR2_X1 _17145_ ( .A1(_10602_ ), .A2(_10605_ ), .ZN(_10606_ ) );
INV_X1 _17146_ ( .A(\idu.io_in_bits_inst [29] ), .ZN(_10607_ ) );
NOR2_X1 _17147_ ( .A1(_10603_ ), .A2(_10607_ ), .ZN(_10608_ ) );
INV_X1 _17148_ ( .A(\idu.io_in_bits_inst [28] ), .ZN(_10609_ ) );
NOR2_X1 _17149_ ( .A1(_10603_ ), .A2(_10609_ ), .ZN(_10610_ ) );
NOR2_X1 _17150_ ( .A1(_10608_ ), .A2(_10610_ ), .ZN(_10611_ ) );
NAND3_X1 _17151_ ( .A1(_10592_ ), .A2(_10606_ ), .A3(_10611_ ), .ZN(_10612_ ) );
INV_X1 _17152_ ( .A(\idu.io_in_bits_inst [22] ), .ZN(_10613_ ) );
NOR2_X1 _17153_ ( .A1(_10576_ ), .A2(_10613_ ), .ZN(\idu.immI [2] ) );
INV_X1 _17154_ ( .A(\idu.io_in_bits_inst [23] ), .ZN(_10614_ ) );
NOR2_X1 _17155_ ( .A1(_10576_ ), .A2(_10614_ ), .ZN(\idu.immI [3] ) );
NOR2_X1 _17156_ ( .A1(\idu.immI [2] ), .A2(\idu.immI [3] ), .ZN(_10615_ ) );
INV_X1 _17157_ ( .A(\idu.io_in_bits_inst [20] ), .ZN(_10616_ ) );
NOR2_X1 _17158_ ( .A1(_10576_ ), .A2(_10616_ ), .ZN(\idu.immI [0] ) );
INV_X1 _17159_ ( .A(\idu.io_in_bits_inst [21] ), .ZN(_10617_ ) );
NOR2_X1 _17160_ ( .A1(_10576_ ), .A2(_10617_ ), .ZN(\idu.immI [1] ) );
NOR2_X1 _17161_ ( .A1(\idu.immI [0] ), .A2(\idu.immI [1] ), .ZN(_10618_ ) );
INV_X1 _17162_ ( .A(\idu.io_in_bits_inst [24] ), .ZN(_10619_ ) );
NOR2_X1 _17163_ ( .A1(_10603_ ), .A2(_10619_ ), .ZN(_10620_ ) );
INV_X1 _17164_ ( .A(_10620_ ), .ZN(_10621_ ) );
NAND3_X1 _17165_ ( .A1(_10615_ ), .A2(_10618_ ), .A3(_10621_ ), .ZN(_10622_ ) );
NOR2_X1 _17166_ ( .A1(_10612_ ), .A2(_10622_ ), .ZN(_10623_ ) );
INV_X1 _17167_ ( .A(\idu.io_in_bits_inst [14] ), .ZN(_10624_ ) );
NOR2_X1 _17168_ ( .A1(_10585_ ), .A2(_10624_ ), .ZN(_10625_ ) );
INV_X1 _17169_ ( .A(_10625_ ), .ZN(_10626_ ) );
INV_X1 _17170_ ( .A(_10575_ ), .ZN(_10627_ ) );
AND2_X1 _17171_ ( .A1(_10627_ ), .A2(\idu.io_in_bits_inst [7] ), .ZN(\idu.immB [11] ) );
INV_X1 _17172_ ( .A(\idu.io_in_bits_inst [15] ), .ZN(_10628_ ) );
NOR2_X1 _17173_ ( .A1(_10585_ ), .A2(_10628_ ), .ZN(_10629_ ) );
NOR2_X1 _17174_ ( .A1(\idu.immB [11] ), .A2(_10629_ ), .ZN(_10630_ ) );
INV_X1 _17175_ ( .A(\idu.io_in_bits_inst [12] ), .ZN(_10631_ ) );
NOR2_X1 _17176_ ( .A1(_10585_ ), .A2(_10631_ ), .ZN(_10632_ ) );
INV_X1 _17177_ ( .A(\idu.io_in_bits_inst [13] ), .ZN(_10633_ ) );
AND2_X1 _17178_ ( .A1(_10632_ ), .A2(_10633_ ), .ZN(_10634_ ) );
INV_X1 _17179_ ( .A(\idu.io_in_bits_inst [5] ), .ZN(_10635_ ) );
INV_X1 _17180_ ( .A(\idu.io_in_bits_inst [6] ), .ZN(_10636_ ) );
NAND2_X1 _17181_ ( .A1(_10635_ ), .A2(_10636_ ), .ZN(_10637_ ) );
OAI21_X1 _17182_ ( .A(_10627_ ), .B1(\idu.io_in_bits_inst [4] ), .B2(_10637_ ), .ZN(_10638_ ) );
AND4_X1 _17183_ ( .A1(_10626_ ), .A2(_10630_ ), .A3(_10634_ ), .A4(_10638_ ), .ZN(_10639_ ) );
AND2_X1 _17184_ ( .A1(_10627_ ), .A2(\idu.io_in_bits_inst [8] ), .ZN(\idu.immB [1] ) );
INV_X1 _17185_ ( .A(\idu.io_in_bits_inst [9] ), .ZN(_10640_ ) );
NOR2_X1 _17186_ ( .A1(_10603_ ), .A2(_10640_ ), .ZN(\idu.immB [2] ) );
INV_X1 _17187_ ( .A(\idu.io_in_bits_inst [10] ), .ZN(_10641_ ) );
NOR2_X1 _17188_ ( .A1(_10585_ ), .A2(_10641_ ), .ZN(\idu.immB [3] ) );
OR3_X1 _17189_ ( .A1(\idu.immB [1] ), .A2(\idu.immB [2] ), .A3(\idu.immB [3] ), .ZN(_10642_ ) );
AND2_X1 _17190_ ( .A1(_10627_ ), .A2(\idu.io_in_bits_inst [11] ), .ZN(\idu.immB [4] ) );
NOR2_X1 _17191_ ( .A1(_10642_ ), .A2(\idu.immB [4] ), .ZN(_10643_ ) );
AND2_X1 _17192_ ( .A1(_10627_ ), .A2(\idu.io_in_bits_inst [0] ), .ZN(_10644_ ) );
AND2_X1 _17193_ ( .A1(_10644_ ), .A2(\idu.io_in_bits_inst [1] ), .ZN(_10645_ ) );
BUF_X4 _17194_ ( .A(_10627_ ), .Z(_10646_ ) );
AND3_X1 _17195_ ( .A1(_10645_ ), .A2(\idu.io_in_bits_inst [2] ), .A3(_10646_ ), .ZN(_10647_ ) );
AND4_X1 _17196_ ( .A1(\idu.io_in_bits_inst [3] ), .A2(_10639_ ), .A3(_10643_ ), .A4(_10647_ ), .ZN(_10648_ ) );
AND2_X1 _17197_ ( .A1(_10623_ ), .A2(_10648_ ), .ZN(\idu.io_out_bits_fencei ) );
INV_X1 _17198_ ( .A(\idu.io_out_bits_fencei ), .ZN(_10649_ ) );
AND2_X1 _17199_ ( .A1(\idu.immI [0] ), .A2(_10617_ ), .ZN(_10650_ ) );
AND2_X2 _17200_ ( .A1(_10650_ ), .A2(_10615_ ), .ZN(_10651_ ) );
AND2_X1 _17201_ ( .A1(_10651_ ), .A2(_10621_ ), .ZN(_10652_ ) );
CLKBUF_X2 _17202_ ( .A(_10611_ ), .Z(_10653_ ) );
CLKBUF_X2 _17203_ ( .A(_10592_ ), .Z(_10654_ ) );
AND4_X1 _17204_ ( .A1(_10606_ ), .A2(_10652_ ), .A3(_10653_ ), .A4(_10654_ ), .ZN(_10655_ ) );
NOR2_X1 _17205_ ( .A1(\idu.io_in_bits_inst [3] ), .A2(\idu.io_in_bits_inst [2] ), .ZN(_10656_ ) );
AND3_X1 _17206_ ( .A1(_10645_ ), .A2(\idu.io_in_bits_inst [6] ), .A3(_10656_ ), .ZN(_10657_ ) );
NOR2_X1 _17207_ ( .A1(_10585_ ), .A2(_10635_ ), .ZN(_10658_ ) );
AND2_X1 _17208_ ( .A1(_10658_ ), .A2(\idu.io_in_bits_inst [4] ), .ZN(_10659_ ) );
AND2_X1 _17209_ ( .A1(_10657_ ), .A2(_10659_ ), .ZN(_10660_ ) );
OAI21_X1 _17210_ ( .A(_10627_ ), .B1(\idu.io_in_bits_inst [13] ), .B2(\idu.io_in_bits_inst [12] ), .ZN(_10661_ ) );
AND2_X1 _17211_ ( .A1(_10661_ ), .A2(_10626_ ), .ZN(_10662_ ) );
AND3_X1 _17212_ ( .A1(_10662_ ), .A2(_10643_ ), .A3(_10630_ ), .ZN(_10663_ ) );
NAND3_X1 _17213_ ( .A1(_10655_ ), .A2(_10660_ ), .A3(_10663_ ), .ZN(_10664_ ) );
NAND3_X1 _17214_ ( .A1(_10649_ ), .A2(\ifu.ren_REG ), .A3(_10664_ ), .ZN(_10665_ ) );
INV_X1 _17215_ ( .A(\idu.io_in_bits_inst [4] ), .ZN(_10666_ ) );
AND2_X2 _17216_ ( .A1(_10658_ ), .A2(_10666_ ), .ZN(_10667_ ) );
NOR2_X1 _17217_ ( .A1(_10585_ ), .A2(_10633_ ), .ZN(_10668_ ) );
AND2_X1 _17218_ ( .A1(_10668_ ), .A2(_10631_ ), .ZN(_10669_ ) );
AND2_X1 _17219_ ( .A1(_10669_ ), .A2(\idu.io_in_bits_inst [14] ), .ZN(_10670_ ) );
AND2_X1 _17220_ ( .A1(_10661_ ), .A2(_10625_ ), .ZN(_10671_ ) );
OAI211_X1 _17221_ ( .A(_10657_ ), .B(_10667_ ), .C1(_10670_ ), .C2(_10671_ ), .ZN(_10672_ ) );
AND2_X2 _17222_ ( .A1(_10645_ ), .A2(_10656_ ), .ZN(_10673_ ) );
AND2_X1 _17223_ ( .A1(_10634_ ), .A2(\idu.io_in_bits_inst [14] ), .ZN(_10674_ ) );
NAND4_X1 _17224_ ( .A1(_10673_ ), .A2(\idu.io_in_bits_inst [6] ), .A3(_10667_ ), .A4(_10674_ ), .ZN(_10675_ ) );
AND2_X2 _17225_ ( .A1(_10667_ ), .A2(\idu.io_in_bits_inst [6] ), .ZN(_10676_ ) );
NAND4_X1 _17226_ ( .A1(_10676_ ), .A2(_10645_ ), .A3(_10656_ ), .A4(_10662_ ), .ZN(_10677_ ) );
AND3_X1 _17227_ ( .A1(_10672_ ), .A2(_10675_ ), .A3(_10677_ ), .ZN(_10678_ ) );
AND2_X1 _17228_ ( .A1(_10632_ ), .A2(\idu.io_in_bits_inst [13] ), .ZN(_10679_ ) );
AND2_X1 _17229_ ( .A1(_10679_ ), .A2(\idu.io_in_bits_inst [14] ), .ZN(_10680_ ) );
AND2_X1 _17230_ ( .A1(_10634_ ), .A2(_10624_ ), .ZN(_10681_ ) );
OAI211_X1 _17231_ ( .A(_10657_ ), .B(_10667_ ), .C1(_10680_ ), .C2(_10681_ ), .ZN(_10682_ ) );
AND2_X1 _17232_ ( .A1(_10678_ ), .A2(_10682_ ), .ZN(_10683_ ) );
AND2_X1 _17233_ ( .A1(_10663_ ), .A2(_10660_ ), .ZN(_10684_ ) );
AND2_X2 _17234_ ( .A1(\idu.immI [1] ), .A2(_10616_ ), .ZN(_10685_ ) );
AND2_X1 _17235_ ( .A1(_10685_ ), .A2(_10615_ ), .ZN(_10686_ ) );
AND2_X2 _17236_ ( .A1(_10686_ ), .A2(_10621_ ), .ZN(_10687_ ) );
INV_X1 _17237_ ( .A(_10687_ ), .ZN(_10688_ ) );
NAND4_X1 _17238_ ( .A1(_10592_ ), .A2(\idu.io_in_bits_inst [28] ), .A3(_10606_ ), .A4(_10608_ ), .ZN(_10689_ ) );
NOR2_X1 _17239_ ( .A1(_10688_ ), .A2(_10689_ ), .ZN(_10690_ ) );
OAI21_X1 _17240_ ( .A(_10684_ ), .B1(_10623_ ), .B2(_10690_ ), .ZN(_10691_ ) );
AND2_X1 _17241_ ( .A1(_10647_ ), .A2(\idu.io_in_bits_inst [3] ), .ZN(_10692_ ) );
AND2_X1 _17242_ ( .A1(_10692_ ), .A2(_10676_ ), .ZN(\idu.io_out_bits_jal ) );
NAND3_X1 _17243_ ( .A1(_10645_ ), .A2(\idu.io_in_bits_inst [2] ), .A3(_10646_ ), .ZN(_10693_ ) );
NOR2_X1 _17244_ ( .A1(_10693_ ), .A2(\idu.io_in_bits_inst [3] ), .ZN(_10694_ ) );
CLKBUF_X2 _17245_ ( .A(_10662_ ), .Z(_10695_ ) );
AND3_X1 _17246_ ( .A1(_10694_ ), .A2(_10695_ ), .A3(_10676_ ), .ZN(\idu.io_out_bits_jalr ) );
NOR2_X1 _17247_ ( .A1(\idu.io_out_bits_jal ), .A2(\idu.io_out_bits_jalr ), .ZN(_10696_ ) );
NAND3_X1 _17248_ ( .A1(_10683_ ), .A2(_10691_ ), .A3(_10696_ ), .ZN(\idu.io_out_bits_en_dnpc ) );
OAI21_X1 _17249_ ( .A(_10573_ ), .B1(_10665_ ), .B2(\idu.io_out_bits_en_dnpc ), .ZN(_10697_ ) );
BUF_X4 _17250_ ( .A(_09463_ ), .Z(_10698_ ) );
BUF_X2 _17251_ ( .A(_10698_ ), .Z(_10699_ ) );
NAND4_X1 _17252_ ( .A1(_10697_ ), .A2(_10699_ ), .A3(\ifu.state [0] ), .A4(_09466_ ), .ZN(_10700_ ) );
INV_X1 _17253_ ( .A(\ifu._start_T_2 [0] ), .ZN(_10701_ ) );
OAI211_X1 _17254_ ( .A(_10699_ ), .B(_10701_ ), .C1(fanout_net_14 ), .C2(fanout_net_15 ), .ZN(_10702_ ) );
AND2_X1 _17255_ ( .A1(_10700_ ), .A2(_10702_ ), .ZN(_10703_ ) );
INV_X1 _17256_ ( .A(_10703_ ), .ZN(_10704_ ) );
MUX2_X1 _17257_ ( .A(\icache.valid_reg_0 ), .B(\icache.valid_reg_1 ), .S(_09818_ ), .Z(_10705_ ) );
AND3_X2 _17258_ ( .A1(_10571_ ), .A2(_10704_ ), .A3(_10705_ ), .ZN(_10706_ ) );
AND2_X1 _17259_ ( .A1(_10706_ ), .A2(fanout_net_13 ), .ZN(_10707_ ) );
BUF_X2 _17260_ ( .A(_10707_ ), .Z(_10708_ ) );
AND2_X1 _17261_ ( .A1(fanout_net_2 ), .A2(io_master_rvalid ), .ZN(\icache.offset_buf_$_SDFFE_PP0P__Q_E ) );
AND2_X1 _17262_ ( .A1(\icache.offset_buf_$_SDFFE_PP0P__Q_E ), .A2(io_master_rlast ), .ZN(_10709_ ) );
NOR2_X4 _17263_ ( .A1(_10708_ ), .A2(_10709_ ), .ZN(_10710_ ) );
INV_X1 _17264_ ( .A(_10710_ ), .ZN(_10711_ ) );
NOR2_X1 _17265_ ( .A1(_10711_ ), .A2(\ifu.state [2] ), .ZN(_10712_ ) );
XNOR2_X1 _17266_ ( .A(\idu.io_in_bits_pc [22] ), .B(\lsu.io_in_bits_pc [22] ), .ZN(_10713_ ) );
XNOR2_X1 _17267_ ( .A(\idu.io_in_bits_pc [23] ), .B(\lsu.io_in_bits_pc [23] ), .ZN(_10714_ ) );
XNOR2_X1 _17268_ ( .A(\idu.io_in_bits_pc [18] ), .B(\lsu.io_in_bits_pc [18] ), .ZN(_10715_ ) );
XNOR2_X1 _17269_ ( .A(\idu.io_in_bits_pc [19] ), .B(\lsu.io_in_bits_pc [19] ), .ZN(_10716_ ) );
AND4_X1 _17270_ ( .A1(_10713_ ), .A2(_10714_ ), .A3(_10715_ ), .A4(_10716_ ), .ZN(_10717_ ) );
XNOR2_X1 _17271_ ( .A(\idu.io_in_bits_pc [25] ), .B(\lsu.io_in_bits_pc [25] ), .ZN(_10718_ ) );
XNOR2_X1 _17272_ ( .A(\idu.io_in_bits_pc [29] ), .B(\lsu.io_in_bits_pc [29] ), .ZN(_10719_ ) );
XNOR2_X1 _17273_ ( .A(\idu.io_in_bits_pc [28] ), .B(\lsu.io_in_bits_pc [28] ), .ZN(_10720_ ) );
XNOR2_X1 _17274_ ( .A(\idu.io_in_bits_pc [24] ), .B(\lsu.io_in_bits_pc [24] ), .ZN(_10721_ ) );
AND4_X1 _17275_ ( .A1(_10718_ ), .A2(_10719_ ), .A3(_10720_ ), .A4(_10721_ ), .ZN(_10722_ ) );
XNOR2_X1 _17276_ ( .A(\idu.io_in_bits_pc [4] ), .B(\lsu.io_in_bits_pc [4] ), .ZN(_10723_ ) );
XNOR2_X1 _17277_ ( .A(\idu.io_in_bits_pc [5] ), .B(\lsu.io_in_bits_pc [5] ), .ZN(_10724_ ) );
XNOR2_X1 _17278_ ( .A(\idu.io_in_bits_pc [1] ), .B(\lsu.io_in_bits_pc [1] ), .ZN(_10725_ ) );
XNOR2_X1 _17279_ ( .A(\idu.io_in_bits_pc [0] ), .B(\lsu.io_in_bits_pc [0] ), .ZN(_10726_ ) );
AND4_X1 _17280_ ( .A1(_10723_ ), .A2(_10724_ ), .A3(_10725_ ), .A4(_10726_ ), .ZN(_10727_ ) );
XNOR2_X1 _17281_ ( .A(\idu.io_in_bits_pc [15] ), .B(\lsu.io_in_bits_pc [15] ), .ZN(_10728_ ) );
XNOR2_X1 _17282_ ( .A(\idu.io_in_bits_pc [14] ), .B(\lsu.io_in_bits_pc [14] ), .ZN(_10729_ ) );
XNOR2_X1 _17283_ ( .A(\idu.io_in_bits_pc [11] ), .B(\lsu.io_in_bits_pc [11] ), .ZN(_10730_ ) );
XNOR2_X1 _17284_ ( .A(\idu.io_in_bits_pc [10] ), .B(\lsu.io_in_bits_pc [10] ), .ZN(_10731_ ) );
AND4_X1 _17285_ ( .A1(_10728_ ), .A2(_10729_ ), .A3(_10730_ ), .A4(_10731_ ), .ZN(_10732_ ) );
AND4_X1 _17286_ ( .A1(_10717_ ), .A2(_10722_ ), .A3(_10727_ ), .A4(_10732_ ), .ZN(_10733_ ) );
XNOR2_X1 _17287_ ( .A(\idu.io_in_bits_pc [17] ), .B(\lsu.io_in_bits_pc [17] ), .ZN(_10734_ ) );
XNOR2_X1 _17288_ ( .A(\idu.io_in_bits_pc [21] ), .B(\lsu.io_in_bits_pc [21] ), .ZN(_10735_ ) );
XNOR2_X1 _17289_ ( .A(\idu.io_in_bits_pc [20] ), .B(\lsu.io_in_bits_pc [20] ), .ZN(_10736_ ) );
XNOR2_X1 _17290_ ( .A(\idu.io_in_bits_pc [16] ), .B(\lsu.io_in_bits_pc [16] ), .ZN(_10737_ ) );
AND4_X1 _17291_ ( .A1(_10734_ ), .A2(_10735_ ), .A3(_10736_ ), .A4(_10737_ ), .ZN(_10738_ ) );
XNOR2_X1 _17292_ ( .A(\idu.io_in_bits_pc [27] ), .B(\lsu.io_in_bits_pc [27] ), .ZN(_10739_ ) );
XNOR2_X1 _17293_ ( .A(\idu.io_in_bits_pc [26] ), .B(\lsu.io_in_bits_pc [26] ), .ZN(_10740_ ) );
XNOR2_X1 _17294_ ( .A(\idu.io_in_bits_pc [31] ), .B(\lsu.io_in_bits_pc [31] ), .ZN(_10741_ ) );
XNOR2_X1 _17295_ ( .A(\idu.io_in_bits_pc [30] ), .B(\lsu.io_in_bits_pc [30] ), .ZN(_10742_ ) );
AND4_X1 _17296_ ( .A1(_10739_ ), .A2(_10740_ ), .A3(_10741_ ), .A4(_10742_ ), .ZN(_10743_ ) );
XNOR2_X1 _17297_ ( .A(\idu.io_in_bits_pc [2] ), .B(\lsu.io_in_bits_pc [2] ), .ZN(_10744_ ) );
XNOR2_X1 _17298_ ( .A(\idu.io_in_bits_pc [3] ), .B(\lsu.io_in_bits_pc [3] ), .ZN(_10745_ ) );
XNOR2_X1 _17299_ ( .A(\idu.io_in_bits_pc [7] ), .B(\lsu.io_in_bits_pc [7] ), .ZN(_10746_ ) );
XNOR2_X1 _17300_ ( .A(\idu.io_in_bits_pc [6] ), .B(\lsu.io_in_bits_pc [6] ), .ZN(_10747_ ) );
AND4_X1 _17301_ ( .A1(_10744_ ), .A2(_10745_ ), .A3(_10746_ ), .A4(_10747_ ), .ZN(_10748_ ) );
XNOR2_X1 _17302_ ( .A(\idu.io_in_bits_pc [8] ), .B(\lsu.io_in_bits_pc [8] ), .ZN(_10749_ ) );
XNOR2_X1 _17303_ ( .A(\idu.io_in_bits_pc [13] ), .B(\lsu.io_in_bits_pc [13] ), .ZN(_10750_ ) );
XNOR2_X1 _17304_ ( .A(\idu.io_in_bits_pc [12] ), .B(\lsu.io_in_bits_pc [12] ), .ZN(_10751_ ) );
XNOR2_X1 _17305_ ( .A(\idu.io_in_bits_pc [9] ), .B(\lsu.io_in_bits_pc [9] ), .ZN(_10752_ ) );
AND4_X1 _17306_ ( .A1(_10749_ ), .A2(_10750_ ), .A3(_10751_ ), .A4(_10752_ ), .ZN(_10753_ ) );
AND4_X1 _17307_ ( .A1(_10738_ ), .A2(_10743_ ), .A3(_10748_ ), .A4(_10753_ ), .ZN(_10754_ ) );
NAND2_X1 _17308_ ( .A1(_10733_ ), .A2(_10754_ ), .ZN(_10755_ ) );
BUF_X4 _17309_ ( .A(_10629_ ), .Z(_10756_ ) );
XNOR2_X1 _17310_ ( .A(_10756_ ), .B(\lsu.io_in_bits_rd [0] ), .ZN(_10757_ ) );
INV_X1 _17311_ ( .A(\lsu.io_in_bits_rd [1] ), .ZN(_10758_ ) );
NAND3_X1 _17312_ ( .A1(_10646_ ), .A2(\idu.io_in_bits_inst [16] ), .A3(_10758_ ), .ZN(_10759_ ) );
BUF_X4 _17313_ ( .A(_10603_ ), .Z(_10760_ ) );
OAI21_X1 _17314_ ( .A(\lsu.io_in_bits_rd [1] ), .B1(_10760_ ), .B2(_10593_ ), .ZN(_10761_ ) );
NAND3_X1 _17315_ ( .A1(_10757_ ), .A2(_10759_ ), .A3(_10761_ ), .ZN(_10762_ ) );
XNOR2_X1 _17316_ ( .A(_10600_ ), .B(\lsu.io_in_bits_rd [3] ), .ZN(_10763_ ) );
XNOR2_X1 _17317_ ( .A(_10597_ ), .B(\lsu.io_in_bits_rd [2] ), .ZN(_10764_ ) );
NAND2_X1 _17318_ ( .A1(_10763_ ), .A2(_10764_ ), .ZN(_10765_ ) );
CLKBUF_X2 _17319_ ( .A(_10605_ ), .Z(_10766_ ) );
BUF_X2 _17320_ ( .A(_10766_ ), .Z(_10767_ ) );
INV_X1 _17321_ ( .A(\lsu.io_in_bits_rd [4] ), .ZN(_10768_ ) );
XNOR2_X1 _17322_ ( .A(_10767_ ), .B(_10768_ ), .ZN(_10769_ ) );
NOR3_X1 _17323_ ( .A1(_10762_ ), .A2(_10765_ ), .A3(_10769_ ), .ZN(_10770_ ) );
NOR4_X1 _17324_ ( .A1(\lsu.io_in_bits_rd [0] ), .A2(\lsu.io_in_bits_rd [1] ), .A3(\lsu.io_in_bits_rd [3] ), .A4(\lsu.io_in_bits_rd [2] ), .ZN(_10771_ ) );
NAND2_X1 _17325_ ( .A1(_10771_ ), .A2(_10768_ ), .ZN(_10772_ ) );
AND2_X1 _17326_ ( .A1(_10770_ ), .A2(_10772_ ), .ZN(_10773_ ) );
XNOR2_X1 _17327_ ( .A(\idu.immI [0] ), .B(\lsu.io_in_bits_rd [0] ), .ZN(_10774_ ) );
OAI21_X1 _17328_ ( .A(\lsu.io_in_bits_rd [1] ), .B1(_10760_ ), .B2(_10617_ ), .ZN(_10775_ ) );
NAND3_X1 _17329_ ( .A1(_10646_ ), .A2(\idu.io_in_bits_inst [21] ), .A3(_10758_ ), .ZN(_10776_ ) );
NAND3_X1 _17330_ ( .A1(_10774_ ), .A2(_10775_ ), .A3(_10776_ ), .ZN(_10777_ ) );
OR3_X1 _17331_ ( .A1(_10603_ ), .A2(_10613_ ), .A3(\lsu.io_in_bits_rd [2] ), .ZN(_10778_ ) );
OR3_X1 _17332_ ( .A1(_10603_ ), .A2(_10614_ ), .A3(\lsu.io_in_bits_rd [3] ), .ZN(_10779_ ) );
OAI21_X1 _17333_ ( .A(\lsu.io_in_bits_rd [2] ), .B1(_10760_ ), .B2(_10613_ ), .ZN(_10780_ ) );
OAI21_X1 _17334_ ( .A(\lsu.io_in_bits_rd [3] ), .B1(_10760_ ), .B2(_10614_ ), .ZN(_10781_ ) );
NAND4_X1 _17335_ ( .A1(_10778_ ), .A2(_10779_ ), .A3(_10780_ ), .A4(_10781_ ), .ZN(_10782_ ) );
CLKBUF_X2 _17336_ ( .A(_10620_ ), .Z(_10783_ ) );
XNOR2_X1 _17337_ ( .A(_10783_ ), .B(_10768_ ), .ZN(_10784_ ) );
NOR3_X1 _17338_ ( .A1(_10777_ ), .A2(_10782_ ), .A3(_10784_ ), .ZN(_10785_ ) );
AND2_X1 _17339_ ( .A1(_10785_ ), .A2(_10772_ ), .ZN(_10786_ ) );
OAI211_X1 _17340_ ( .A(\lsu.io_in_valid ), .B(_10755_ ), .C1(_10773_ ), .C2(_10786_ ), .ZN(_10787_ ) );
OR3_X1 _17341_ ( .A1(_wbu_io_in_bits_T ), .A2(\idu.io_raw_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B ), .A3(_10787_ ), .ZN(_10788_ ) );
OAI21_X1 _17342_ ( .A(\exu.io_in_bits_rd [0] ), .B1(_10603_ ), .B2(_10628_ ), .ZN(_10789_ ) );
OAI21_X1 _17343_ ( .A(_10789_ ), .B1(_10598_ ), .B2(\exu.io_in_bits_rd [2] ), .ZN(_10790_ ) );
INV_X1 _17344_ ( .A(\exu.io_in_bits_rd [1] ), .ZN(_10791_ ) );
BUF_X4 _17345_ ( .A(_10594_ ), .Z(_10792_ ) );
AOI221_X4 _17346_ ( .A(_10790_ ), .B1(_10791_ ), .B2(_10792_ ), .C1(\exu.io_in_bits_rd [2] ), .C2(_10598_ ), .ZN(_10793_ ) );
INV_X1 _17347_ ( .A(\exu.io_in_bits_rd [4] ), .ZN(_10794_ ) );
AOI21_X1 _17348_ ( .A(_10794_ ), .B1(_10646_ ), .B2(\idu.io_in_bits_inst [19] ), .ZN(_10795_ ) );
NOR3_X1 _17349_ ( .A1(_10760_ ), .A2(\exu.io_in_bits_rd [4] ), .A3(_10604_ ), .ZN(_10796_ ) );
NOR3_X1 _17350_ ( .A1(_10760_ ), .A2(\exu.io_in_bits_rd [0] ), .A3(_10628_ ), .ZN(_10797_ ) );
NOR3_X1 _17351_ ( .A1(_10795_ ), .A2(_10796_ ), .A3(_10797_ ), .ZN(_10798_ ) );
OAI22_X1 _17352_ ( .A1(_10601_ ), .A2(\exu.io_in_bits_rd [3] ), .B1(_10791_ ), .B2(_10792_ ), .ZN(_10799_ ) );
INV_X1 _17353_ ( .A(\exu.io_in_bits_rd [3] ), .ZN(_10800_ ) );
AOI21_X1 _17354_ ( .A(_10800_ ), .B1(_10646_ ), .B2(\idu.io_in_bits_inst [18] ), .ZN(_10801_ ) );
NOR4_X1 _17355_ ( .A1(\exu.io_in_bits_rd [0] ), .A2(\exu.io_in_bits_rd [1] ), .A3(\exu.io_in_bits_rd [3] ), .A4(\exu.io_in_bits_rd [2] ), .ZN(_10802_ ) );
AND2_X1 _17356_ ( .A1(_10802_ ), .A2(_10794_ ), .ZN(_10803_ ) );
NOR3_X1 _17357_ ( .A1(_10799_ ), .A2(_10801_ ), .A3(_10803_ ), .ZN(_10804_ ) );
AND3_X1 _17358_ ( .A1(_10793_ ), .A2(_10798_ ), .A3(_10804_ ), .ZN(_10805_ ) );
INV_X1 _17359_ ( .A(_10805_ ), .ZN(_10806_ ) );
XNOR2_X1 _17360_ ( .A(\idu.immI [0] ), .B(\exu.io_in_bits_rd [0] ), .ZN(_10807_ ) );
XNOR2_X1 _17361_ ( .A(\idu.immI [3] ), .B(\exu.io_in_bits_rd [3] ), .ZN(_10808_ ) );
XNOR2_X1 _17362_ ( .A(\idu.immI [1] ), .B(\exu.io_in_bits_rd [1] ), .ZN(_10809_ ) );
XNOR2_X1 _17363_ ( .A(\idu.immI [2] ), .B(\exu.io_in_bits_rd [2] ), .ZN(_10810_ ) );
NAND4_X1 _17364_ ( .A1(_10807_ ), .A2(_10808_ ), .A3(_10809_ ), .A4(_10810_ ), .ZN(_10811_ ) );
CLKBUF_X2 _17365_ ( .A(_10783_ ), .Z(_10812_ ) );
XNOR2_X1 _17366_ ( .A(_10812_ ), .B(_10794_ ), .ZN(_10813_ ) );
OR3_X1 _17367_ ( .A1(_10811_ ), .A2(_10803_ ), .A3(_10813_ ), .ZN(_10814_ ) );
AOI21_X1 _17368_ ( .A(exu_io_in_valid_REG_$_NOT__A_Y ), .B1(_10806_ ), .B2(_10814_ ), .ZN(_10815_ ) );
AND2_X1 _17369_ ( .A1(_09013_ ), .A2(_09034_ ), .ZN(_10816_ ) );
INV_X1 _17370_ ( .A(_10816_ ), .ZN(_10817_ ) );
NOR3_X1 _17371_ ( .A1(\exu.io_in_bits_lb ), .A2(\exu.io_in_bits_lw ), .A3(\exu.io_in_bits_lbu ), .ZN(_10818_ ) );
NOR2_X1 _17372_ ( .A1(\exu.io_in_bits_lhu ), .A2(\exu.io_in_bits_lh ), .ZN(_10819_ ) );
AND2_X1 _17373_ ( .A1(_10818_ ), .A2(_10819_ ), .ZN(_10820_ ) );
INV_X1 _17374_ ( .A(_10820_ ), .ZN(_10821_ ) );
BUF_X2 _17375_ ( .A(_10821_ ), .Z(\exu.io_out_bits_ren ) );
NAND3_X1 _17376_ ( .A1(_10815_ ), .A2(_10817_ ), .A3(\exu.io_out_bits_ren ), .ZN(_10822_ ) );
AND2_X1 _17377_ ( .A1(\lsu.io_in_valid ), .A2(\lsu.io_in_bits_ren ), .ZN(_10823_ ) );
AND2_X1 _17378_ ( .A1(\lsu.io_in_valid ), .A2(\lsu.io_in_bits_wen ), .ZN(_10824_ ) );
NOR2_X1 _17379_ ( .A1(_10823_ ), .A2(_10824_ ), .ZN(_10825_ ) );
AND2_X1 _17380_ ( .A1(_10825_ ), .A2(\lsu._io_in_ready_T ), .ZN(_10826_ ) );
INV_X1 _17381_ ( .A(\exu.state ), .ZN(_10827_ ) );
AND2_X1 _17382_ ( .A1(_10826_ ), .A2(_10827_ ), .ZN(_10828_ ) );
AND3_X1 _17383_ ( .A1(_10788_ ), .A2(_10822_ ), .A3(_10828_ ), .ZN(_10829_ ) );
INV_X1 _17384_ ( .A(\idu.state ), .ZN(_10830_ ) );
AND2_X2 _17385_ ( .A1(_10829_ ), .A2(_10830_ ), .ZN(_10831_ ) );
INV_X1 _17386_ ( .A(_10831_ ), .ZN(_10832_ ) );
NOR2_X4 _17387_ ( .A1(_10712_ ), .A2(_10832_ ), .ZN(_10833_ ) );
BUF_X2 _17388_ ( .A(_10833_ ), .Z(_idu_io_in_bits_T ) );
BUF_X2 _17389_ ( .A(_09870_ ), .Z(_10834_ ) );
BUF_X2 _17390_ ( .A(_10834_ ), .Z(_10835_ ) );
BUF_X2 _17391_ ( .A(_10835_ ), .Z(_10836_ ) );
CLKBUF_X2 _17392_ ( .A(_10836_ ), .Z(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__A_Y ) );
BUF_X2 _17393_ ( .A(_09818_ ), .Z(_10837_ ) );
BUF_X2 _17394_ ( .A(_10837_ ), .Z(_10838_ ) );
BUF_X2 _17395_ ( .A(_10838_ ), .Z(_10839_ ) );
BUF_X2 _17396_ ( .A(_10839_ ), .Z(_10840_ ) );
CLKBUF_X2 _17397_ ( .A(_10840_ ), .Z(_10841_ ) );
CLKBUF_X2 _17398_ ( .A(_10841_ ), .Z(\arbiter.io_ifu_araddr [4] ) );
BUF_X2 _17399_ ( .A(_10699_ ), .Z(_10842_ ) );
CLKBUF_X2 _17400_ ( .A(_10842_ ), .Z(_10843_ ) );
BUF_X2 _17401_ ( .A(_10843_ ), .Z(_10844_ ) );
BUF_X4 _17402_ ( .A(_10844_ ), .Z(_10845_ ) );
BUF_X4 _17403_ ( .A(_10845_ ), .Z(_10846_ ) );
CLKBUF_X2 _17404_ ( .A(_10846_ ), .Z(_10847_ ) );
AND2_X4 _17405_ ( .A1(\arbiter.clink.mtime [1] ), .A2(\arbiter.clink.mtime [0] ), .ZN(_10848_ ) );
AND2_X4 _17406_ ( .A1(_10848_ ), .A2(\arbiter.clink.mtime [2] ), .ZN(_10849_ ) );
AND2_X4 _17407_ ( .A1(_10849_ ), .A2(\arbiter.clink.mtime [3] ), .ZN(_10850_ ) );
AND2_X4 _17408_ ( .A1(_10850_ ), .A2(\arbiter.clink.mtime [4] ), .ZN(_10851_ ) );
AND2_X4 _17409_ ( .A1(_10851_ ), .A2(\arbiter.clink.mtime [5] ), .ZN(_10852_ ) );
AND2_X4 _17410_ ( .A1(_10852_ ), .A2(\arbiter.clink.mtime [6] ), .ZN(_10853_ ) );
AND2_X4 _17411_ ( .A1(_10853_ ), .A2(\arbiter.clink.mtime [7] ), .ZN(_10854_ ) );
AND2_X4 _17412_ ( .A1(_10854_ ), .A2(\arbiter.clink.mtime [8] ), .ZN(_10855_ ) );
AND2_X4 _17413_ ( .A1(_10855_ ), .A2(\arbiter.clink.mtime [9] ), .ZN(_10856_ ) );
AND2_X4 _17414_ ( .A1(_10856_ ), .A2(\arbiter.clink.mtime [10] ), .ZN(_10857_ ) );
AND2_X4 _17415_ ( .A1(_10857_ ), .A2(\arbiter.clink.mtime [11] ), .ZN(_10858_ ) );
AND2_X4 _17416_ ( .A1(_10858_ ), .A2(\arbiter.clink.mtime [12] ), .ZN(_10859_ ) );
AND2_X4 _17417_ ( .A1(_10859_ ), .A2(\arbiter.clink.mtime [13] ), .ZN(_10860_ ) );
AND2_X4 _17418_ ( .A1(_10860_ ), .A2(\arbiter.clink.mtime [14] ), .ZN(_10861_ ) );
AND2_X4 _17419_ ( .A1(_10861_ ), .A2(\arbiter.clink.mtime [15] ), .ZN(_10862_ ) );
AND2_X4 _17420_ ( .A1(_10862_ ), .A2(\arbiter.clink.mtime [16] ), .ZN(_10863_ ) );
AND2_X4 _17421_ ( .A1(_10863_ ), .A2(\arbiter.clink.mtime [17] ), .ZN(_10864_ ) );
AND2_X4 _17422_ ( .A1(_10864_ ), .A2(\arbiter.clink.mtime [18] ), .ZN(_10865_ ) );
AND2_X4 _17423_ ( .A1(_10865_ ), .A2(\arbiter.clink.mtime [19] ), .ZN(_10866_ ) );
AND2_X4 _17424_ ( .A1(_10866_ ), .A2(\arbiter.clink.mtime [20] ), .ZN(_10867_ ) );
AND2_X4 _17425_ ( .A1(_10867_ ), .A2(\arbiter.clink.mtime [21] ), .ZN(_10868_ ) );
AND2_X4 _17426_ ( .A1(_10868_ ), .A2(\arbiter.clink.mtime [22] ), .ZN(_10869_ ) );
AND2_X4 _17427_ ( .A1(_10869_ ), .A2(\arbiter.clink.mtime [23] ), .ZN(_10870_ ) );
AND2_X4 _17428_ ( .A1(_10870_ ), .A2(\arbiter.clink.mtime [24] ), .ZN(_10871_ ) );
AND2_X4 _17429_ ( .A1(_10871_ ), .A2(\arbiter.clink.mtime [25] ), .ZN(_10872_ ) );
AND2_X4 _17430_ ( .A1(_10872_ ), .A2(\arbiter.clink.mtime [26] ), .ZN(_10873_ ) );
AND2_X4 _17431_ ( .A1(_10873_ ), .A2(\arbiter.clink.mtime [27] ), .ZN(_10874_ ) );
AND2_X4 _17432_ ( .A1(_10874_ ), .A2(\arbiter.clink.mtime [28] ), .ZN(_10875_ ) );
AND2_X4 _17433_ ( .A1(_10875_ ), .A2(\arbiter.clink.mtime [29] ), .ZN(_10876_ ) );
AND2_X4 _17434_ ( .A1(_10876_ ), .A2(\arbiter.clink.mtime [30] ), .ZN(_10877_ ) );
AND2_X4 _17435_ ( .A1(_10877_ ), .A2(\arbiter.clink.mtime [31] ), .ZN(_10878_ ) );
AND2_X4 _17436_ ( .A1(_10878_ ), .A2(\arbiter.clink.mtime [32] ), .ZN(_10879_ ) );
AND2_X4 _17437_ ( .A1(_10879_ ), .A2(\arbiter.clink.mtime [33] ), .ZN(_10880_ ) );
AND2_X4 _17438_ ( .A1(_10880_ ), .A2(\arbiter.clink.mtime [34] ), .ZN(_10881_ ) );
AND2_X4 _17439_ ( .A1(_10881_ ), .A2(\arbiter.clink.mtime [35] ), .ZN(_10882_ ) );
AND2_X4 _17440_ ( .A1(_10882_ ), .A2(\arbiter.clink.mtime [36] ), .ZN(_10883_ ) );
AND2_X4 _17441_ ( .A1(_10883_ ), .A2(\arbiter.clink.mtime [37] ), .ZN(_10884_ ) );
AND2_X4 _17442_ ( .A1(_10884_ ), .A2(\arbiter.clink.mtime [38] ), .ZN(_10885_ ) );
AND2_X4 _17443_ ( .A1(_10885_ ), .A2(\arbiter.clink.mtime [39] ), .ZN(_10886_ ) );
AND2_X4 _17444_ ( .A1(_10886_ ), .A2(\arbiter.clink.mtime [40] ), .ZN(_10887_ ) );
AND2_X4 _17445_ ( .A1(_10887_ ), .A2(\arbiter.clink.mtime [41] ), .ZN(_10888_ ) );
AND2_X4 _17446_ ( .A1(_10888_ ), .A2(\arbiter.clink.mtime [42] ), .ZN(_10889_ ) );
AND2_X4 _17447_ ( .A1(_10889_ ), .A2(\arbiter.clink.mtime [43] ), .ZN(_10890_ ) );
AND2_X4 _17448_ ( .A1(_10890_ ), .A2(\arbiter.clink.mtime [44] ), .ZN(_10891_ ) );
AND2_X4 _17449_ ( .A1(_10891_ ), .A2(\arbiter.clink.mtime [45] ), .ZN(_10892_ ) );
AND2_X4 _17450_ ( .A1(_10892_ ), .A2(\arbiter.clink.mtime [46] ), .ZN(_10893_ ) );
AND2_X4 _17451_ ( .A1(_10893_ ), .A2(\arbiter.clink.mtime [47] ), .ZN(_10894_ ) );
AND2_X4 _17452_ ( .A1(_10894_ ), .A2(\arbiter.clink.mtime [48] ), .ZN(_10895_ ) );
AND2_X4 _17453_ ( .A1(_10895_ ), .A2(\arbiter.clink.mtime [49] ), .ZN(_10896_ ) );
AND2_X4 _17454_ ( .A1(_10896_ ), .A2(\arbiter.clink.mtime [50] ), .ZN(_10897_ ) );
AND2_X4 _17455_ ( .A1(_10897_ ), .A2(\arbiter.clink.mtime [51] ), .ZN(_10898_ ) );
AND2_X4 _17456_ ( .A1(_10898_ ), .A2(\arbiter.clink.mtime [52] ), .ZN(_10899_ ) );
AND2_X4 _17457_ ( .A1(_10899_ ), .A2(\arbiter.clink.mtime [53] ), .ZN(_10900_ ) );
AND2_X4 _17458_ ( .A1(_10900_ ), .A2(\arbiter.clink.mtime [54] ), .ZN(_10901_ ) );
AND2_X4 _17459_ ( .A1(_10901_ ), .A2(\arbiter.clink.mtime [55] ), .ZN(_10902_ ) );
AND2_X4 _17460_ ( .A1(_10902_ ), .A2(\arbiter.clink.mtime [56] ), .ZN(_10903_ ) );
NAND2_X4 _17461_ ( .A1(_10903_ ), .A2(\arbiter.clink.mtime [57] ), .ZN(_10904_ ) );
INV_X1 _17462_ ( .A(\arbiter.clink.mtime [58] ), .ZN(_10905_ ) );
NOR2_X4 _17463_ ( .A1(_10904_ ), .A2(_10905_ ), .ZN(_10906_ ) );
NAND2_X4 _17464_ ( .A1(_10906_ ), .A2(\arbiter.clink.mtime [59] ), .ZN(_10907_ ) );
INV_X1 _17465_ ( .A(\arbiter.clink.mtime [60] ), .ZN(_10908_ ) );
NOR2_X4 _17466_ ( .A1(_10907_ ), .A2(_10908_ ), .ZN(_10909_ ) );
NAND2_X4 _17467_ ( .A1(_10909_ ), .A2(\arbiter.clink.mtime [61] ), .ZN(_10910_ ) );
INV_X1 _17468_ ( .A(\arbiter.clink.mtime [62] ), .ZN(_10911_ ) );
NOR2_X2 _17469_ ( .A1(_10910_ ), .A2(_10911_ ), .ZN(_10912_ ) );
OAI21_X1 _17470_ ( .A(_10847_ ), .B1(_10912_ ), .B2(\arbiter.clink.mtime [63] ), .ZN(_10913_ ) );
INV_X2 _17471_ ( .A(_10910_ ), .ZN(_10914_ ) );
AND3_X2 _17472_ ( .A1(_10914_ ), .A2(\arbiter.clink.mtime [63] ), .A3(\arbiter.clink.mtime [62] ), .ZN(_10915_ ) );
NOR2_X1 _17473_ ( .A1(_10913_ ), .A2(_10915_ ), .ZN(_00034_ ) );
OAI21_X1 _17474_ ( .A(_10847_ ), .B1(_10914_ ), .B2(\arbiter.clink.mtime [62] ), .ZN(_10916_ ) );
NOR2_X1 _17475_ ( .A1(_10916_ ), .A2(_10912_ ), .ZN(_00035_ ) );
BUF_X2 _17476_ ( .A(_10846_ ), .Z(_10917_ ) );
OAI21_X1 _17477_ ( .A(_10917_ ), .B1(_10899_ ), .B2(\arbiter.clink.mtime [53] ), .ZN(_10918_ ) );
NOR2_X1 _17478_ ( .A1(_10900_ ), .A2(_10918_ ), .ZN(_00036_ ) );
OAI21_X1 _17479_ ( .A(_10917_ ), .B1(_10898_ ), .B2(\arbiter.clink.mtime [52] ), .ZN(_10919_ ) );
NOR2_X1 _17480_ ( .A1(_10899_ ), .A2(_10919_ ), .ZN(_00037_ ) );
OAI21_X1 _17481_ ( .A(_10917_ ), .B1(_10897_ ), .B2(\arbiter.clink.mtime [51] ), .ZN(_10920_ ) );
NOR2_X1 _17482_ ( .A1(_10898_ ), .A2(_10920_ ), .ZN(_00038_ ) );
OAI21_X1 _17483_ ( .A(_10917_ ), .B1(_10896_ ), .B2(\arbiter.clink.mtime [50] ), .ZN(_10921_ ) );
NOR2_X1 _17484_ ( .A1(_10897_ ), .A2(_10921_ ), .ZN(_00039_ ) );
BUF_X4 _17485_ ( .A(_10845_ ), .Z(_10922_ ) );
BUF_X4 _17486_ ( .A(_10922_ ), .Z(_10923_ ) );
OAI21_X1 _17487_ ( .A(_10923_ ), .B1(_10895_ ), .B2(\arbiter.clink.mtime [49] ), .ZN(_10924_ ) );
NOR2_X1 _17488_ ( .A1(_10896_ ), .A2(_10924_ ), .ZN(_00040_ ) );
OAI21_X1 _17489_ ( .A(_10923_ ), .B1(_10894_ ), .B2(\arbiter.clink.mtime [48] ), .ZN(_10925_ ) );
NOR2_X1 _17490_ ( .A1(_10895_ ), .A2(_10925_ ), .ZN(_00041_ ) );
AOI21_X1 _17491_ ( .A(\arbiter.clink.mtime [47] ), .B1(_10892_ ), .B2(\arbiter.clink.mtime [46] ), .ZN(_10926_ ) );
NOR3_X1 _17492_ ( .A1(_10894_ ), .A2(fanout_net_19 ), .A3(_10926_ ), .ZN(_00042_ ) );
OAI21_X1 _17493_ ( .A(_10923_ ), .B1(_10892_ ), .B2(\arbiter.clink.mtime [46] ), .ZN(_10927_ ) );
NOR2_X1 _17494_ ( .A1(_10893_ ), .A2(_10927_ ), .ZN(_00043_ ) );
AOI21_X1 _17495_ ( .A(\arbiter.clink.mtime [45] ), .B1(_10890_ ), .B2(\arbiter.clink.mtime [44] ), .ZN(_10928_ ) );
NOR3_X1 _17496_ ( .A1(_10892_ ), .A2(fanout_net_19 ), .A3(_10928_ ), .ZN(_00044_ ) );
OAI21_X1 _17497_ ( .A(_10923_ ), .B1(_10890_ ), .B2(\arbiter.clink.mtime [44] ), .ZN(_10929_ ) );
NOR2_X1 _17498_ ( .A1(_10891_ ), .A2(_10929_ ), .ZN(_00045_ ) );
OAI21_X1 _17499_ ( .A(_10923_ ), .B1(_10909_ ), .B2(\arbiter.clink.mtime [61] ), .ZN(_10930_ ) );
NOR2_X1 _17500_ ( .A1(_10914_ ), .A2(_10930_ ), .ZN(_00046_ ) );
OAI21_X1 _17501_ ( .A(_10923_ ), .B1(_10889_ ), .B2(\arbiter.clink.mtime [43] ), .ZN(_10931_ ) );
NOR2_X1 _17502_ ( .A1(_10890_ ), .A2(_10931_ ), .ZN(_00047_ ) );
OAI21_X1 _17503_ ( .A(_10923_ ), .B1(_10888_ ), .B2(\arbiter.clink.mtime [42] ), .ZN(_10932_ ) );
NOR2_X1 _17504_ ( .A1(_10889_ ), .A2(_10932_ ), .ZN(_00048_ ) );
OAI21_X1 _17505_ ( .A(_10923_ ), .B1(_10887_ ), .B2(\arbiter.clink.mtime [41] ), .ZN(_10933_ ) );
NOR2_X1 _17506_ ( .A1(_10888_ ), .A2(_10933_ ), .ZN(_00049_ ) );
OAI21_X1 _17507_ ( .A(_10923_ ), .B1(_10886_ ), .B2(\arbiter.clink.mtime [40] ), .ZN(_10934_ ) );
NOR2_X1 _17508_ ( .A1(_10887_ ), .A2(_10934_ ), .ZN(_00050_ ) );
AOI21_X1 _17509_ ( .A(\arbiter.clink.mtime [39] ), .B1(_10884_ ), .B2(\arbiter.clink.mtime [38] ), .ZN(_10935_ ) );
NOR3_X1 _17510_ ( .A1(_10886_ ), .A2(fanout_net_19 ), .A3(_10935_ ), .ZN(_00051_ ) );
OAI21_X1 _17511_ ( .A(_10923_ ), .B1(_10884_ ), .B2(\arbiter.clink.mtime [38] ), .ZN(_10936_ ) );
NOR2_X1 _17512_ ( .A1(_10885_ ), .A2(_10936_ ), .ZN(_00052_ ) );
BUF_X4 _17513_ ( .A(_10922_ ), .Z(_10937_ ) );
OAI21_X1 _17514_ ( .A(_10937_ ), .B1(_10883_ ), .B2(\arbiter.clink.mtime [37] ), .ZN(_10938_ ) );
NOR2_X1 _17515_ ( .A1(_10884_ ), .A2(_10938_ ), .ZN(_00053_ ) );
OAI21_X1 _17516_ ( .A(_10937_ ), .B1(_10882_ ), .B2(\arbiter.clink.mtime [36] ), .ZN(_10939_ ) );
NOR2_X1 _17517_ ( .A1(_10883_ ), .A2(_10939_ ), .ZN(_00054_ ) );
OAI21_X1 _17518_ ( .A(_10937_ ), .B1(_10881_ ), .B2(\arbiter.clink.mtime [35] ), .ZN(_10940_ ) );
NOR2_X1 _17519_ ( .A1(_10882_ ), .A2(_10940_ ), .ZN(_00055_ ) );
OAI21_X1 _17520_ ( .A(_10937_ ), .B1(_10880_ ), .B2(\arbiter.clink.mtime [34] ), .ZN(_10941_ ) );
NOR2_X1 _17521_ ( .A1(_10881_ ), .A2(_10941_ ), .ZN(_00056_ ) );
INV_X1 _17522_ ( .A(_10907_ ), .ZN(_10942_ ) );
OAI21_X1 _17523_ ( .A(_10847_ ), .B1(_10942_ ), .B2(\arbiter.clink.mtime [60] ), .ZN(_10943_ ) );
NOR2_X1 _17524_ ( .A1(_10943_ ), .A2(_10909_ ), .ZN(_00057_ ) );
OAI21_X1 _17525_ ( .A(_10937_ ), .B1(_10879_ ), .B2(\arbiter.clink.mtime [33] ), .ZN(_10944_ ) );
NOR2_X1 _17526_ ( .A1(_10880_ ), .A2(_10944_ ), .ZN(_00058_ ) );
OAI21_X1 _17527_ ( .A(_10937_ ), .B1(_10878_ ), .B2(\arbiter.clink.mtime [32] ), .ZN(_10945_ ) );
NOR2_X1 _17528_ ( .A1(_10879_ ), .A2(_10945_ ), .ZN(_00059_ ) );
AOI21_X1 _17529_ ( .A(\arbiter.clink.mtime [31] ), .B1(_10876_ ), .B2(\arbiter.clink.mtime [30] ), .ZN(_10946_ ) );
NOR3_X1 _17530_ ( .A1(_10878_ ), .A2(fanout_net_19 ), .A3(_10946_ ), .ZN(_00060_ ) );
OAI21_X1 _17531_ ( .A(_10937_ ), .B1(_10876_ ), .B2(\arbiter.clink.mtime [30] ), .ZN(_10947_ ) );
NOR2_X1 _17532_ ( .A1(_10877_ ), .A2(_10947_ ), .ZN(_00061_ ) );
AOI21_X1 _17533_ ( .A(\arbiter.clink.mtime [29] ), .B1(_10874_ ), .B2(\arbiter.clink.mtime [28] ), .ZN(_10948_ ) );
NOR3_X1 _17534_ ( .A1(_10876_ ), .A2(fanout_net_19 ), .A3(_10948_ ), .ZN(_00062_ ) );
OAI21_X1 _17535_ ( .A(_10937_ ), .B1(_10874_ ), .B2(\arbiter.clink.mtime [28] ), .ZN(_10949_ ) );
NOR2_X1 _17536_ ( .A1(_10875_ ), .A2(_10949_ ), .ZN(_00063_ ) );
OAI21_X1 _17537_ ( .A(_10937_ ), .B1(_10873_ ), .B2(\arbiter.clink.mtime [27] ), .ZN(_10950_ ) );
NOR2_X1 _17538_ ( .A1(_10874_ ), .A2(_10950_ ), .ZN(_00064_ ) );
OAI21_X1 _17539_ ( .A(_10937_ ), .B1(_10872_ ), .B2(\arbiter.clink.mtime [26] ), .ZN(_10951_ ) );
NOR2_X1 _17540_ ( .A1(_10873_ ), .A2(_10951_ ), .ZN(_00065_ ) );
BUF_X4 _17541_ ( .A(_10922_ ), .Z(_10952_ ) );
OAI21_X1 _17542_ ( .A(_10952_ ), .B1(_10871_ ), .B2(\arbiter.clink.mtime [25] ), .ZN(_10953_ ) );
NOR2_X1 _17543_ ( .A1(_10872_ ), .A2(_10953_ ), .ZN(_00066_ ) );
OAI21_X1 _17544_ ( .A(_10952_ ), .B1(_10870_ ), .B2(\arbiter.clink.mtime [24] ), .ZN(_10954_ ) );
NOR2_X1 _17545_ ( .A1(_10871_ ), .A2(_10954_ ), .ZN(_00067_ ) );
OAI21_X1 _17546_ ( .A(_10952_ ), .B1(_10906_ ), .B2(\arbiter.clink.mtime [59] ), .ZN(_10955_ ) );
NOR2_X1 _17547_ ( .A1(_10942_ ), .A2(_10955_ ), .ZN(_00068_ ) );
AOI21_X1 _17548_ ( .A(\arbiter.clink.mtime [23] ), .B1(_10868_ ), .B2(\arbiter.clink.mtime [22] ), .ZN(_10956_ ) );
NOR3_X1 _17549_ ( .A1(_10870_ ), .A2(fanout_net_19 ), .A3(_10956_ ), .ZN(_00069_ ) );
OAI21_X1 _17550_ ( .A(_10952_ ), .B1(_10868_ ), .B2(\arbiter.clink.mtime [22] ), .ZN(_10957_ ) );
NOR2_X1 _17551_ ( .A1(_10869_ ), .A2(_10957_ ), .ZN(_00070_ ) );
OAI21_X1 _17552_ ( .A(_10952_ ), .B1(_10867_ ), .B2(\arbiter.clink.mtime [21] ), .ZN(_10958_ ) );
NOR2_X1 _17553_ ( .A1(_10868_ ), .A2(_10958_ ), .ZN(_00071_ ) );
OAI21_X1 _17554_ ( .A(_10952_ ), .B1(_10866_ ), .B2(\arbiter.clink.mtime [20] ), .ZN(_10959_ ) );
NOR2_X1 _17555_ ( .A1(_10867_ ), .A2(_10959_ ), .ZN(_00072_ ) );
OAI21_X1 _17556_ ( .A(_10952_ ), .B1(_10865_ ), .B2(\arbiter.clink.mtime [19] ), .ZN(_10960_ ) );
NOR2_X1 _17557_ ( .A1(_10866_ ), .A2(_10960_ ), .ZN(_00073_ ) );
OAI21_X1 _17558_ ( .A(_10952_ ), .B1(_10864_ ), .B2(\arbiter.clink.mtime [18] ), .ZN(_10961_ ) );
NOR2_X1 _17559_ ( .A1(_10865_ ), .A2(_10961_ ), .ZN(_00074_ ) );
OAI21_X1 _17560_ ( .A(_10952_ ), .B1(_10863_ ), .B2(\arbiter.clink.mtime [17] ), .ZN(_10962_ ) );
NOR2_X1 _17561_ ( .A1(_10864_ ), .A2(_10962_ ), .ZN(_00075_ ) );
OAI21_X1 _17562_ ( .A(_10952_ ), .B1(_10862_ ), .B2(\arbiter.clink.mtime [16] ), .ZN(_10963_ ) );
NOR2_X1 _17563_ ( .A1(_10863_ ), .A2(_10963_ ), .ZN(_00076_ ) );
AOI21_X1 _17564_ ( .A(\arbiter.clink.mtime [15] ), .B1(_10860_ ), .B2(\arbiter.clink.mtime [14] ), .ZN(_10964_ ) );
NOR3_X1 _17565_ ( .A1(_10862_ ), .A2(fanout_net_19 ), .A3(_10964_ ), .ZN(_00077_ ) );
BUF_X4 _17566_ ( .A(_10922_ ), .Z(_10965_ ) );
OAI21_X1 _17567_ ( .A(_10965_ ), .B1(_10860_ ), .B2(\arbiter.clink.mtime [14] ), .ZN(_10966_ ) );
NOR2_X1 _17568_ ( .A1(_10861_ ), .A2(_10966_ ), .ZN(_00078_ ) );
INV_X1 _17569_ ( .A(_10904_ ), .ZN(_10967_ ) );
OAI21_X1 _17570_ ( .A(_10847_ ), .B1(_10967_ ), .B2(\arbiter.clink.mtime [58] ), .ZN(_10968_ ) );
NOR2_X1 _17571_ ( .A1(_10968_ ), .A2(_10906_ ), .ZN(_00079_ ) );
AOI21_X1 _17572_ ( .A(\arbiter.clink.mtime [13] ), .B1(_10858_ ), .B2(\arbiter.clink.mtime [12] ), .ZN(_10969_ ) );
NOR3_X1 _17573_ ( .A1(_10860_ ), .A2(fanout_net_19 ), .A3(_10969_ ), .ZN(_00080_ ) );
OAI21_X1 _17574_ ( .A(_10965_ ), .B1(_10858_ ), .B2(\arbiter.clink.mtime [12] ), .ZN(_10970_ ) );
NOR2_X1 _17575_ ( .A1(_10859_ ), .A2(_10970_ ), .ZN(_00081_ ) );
OAI21_X1 _17576_ ( .A(_10965_ ), .B1(_10857_ ), .B2(\arbiter.clink.mtime [11] ), .ZN(_10971_ ) );
NOR2_X1 _17577_ ( .A1(_10858_ ), .A2(_10971_ ), .ZN(_00082_ ) );
OAI21_X1 _17578_ ( .A(_10965_ ), .B1(_10856_ ), .B2(\arbiter.clink.mtime [10] ), .ZN(_10972_ ) );
NOR2_X1 _17579_ ( .A1(_10857_ ), .A2(_10972_ ), .ZN(_00083_ ) );
OAI21_X1 _17580_ ( .A(_10965_ ), .B1(_10855_ ), .B2(\arbiter.clink.mtime [9] ), .ZN(_10973_ ) );
NOR2_X1 _17581_ ( .A1(_10856_ ), .A2(_10973_ ), .ZN(_00084_ ) );
OAI21_X1 _17582_ ( .A(_10965_ ), .B1(_10854_ ), .B2(\arbiter.clink.mtime [8] ), .ZN(_10974_ ) );
NOR2_X1 _17583_ ( .A1(_10855_ ), .A2(_10974_ ), .ZN(_00085_ ) );
OAI21_X1 _17584_ ( .A(_10965_ ), .B1(_10853_ ), .B2(\arbiter.clink.mtime [7] ), .ZN(_10975_ ) );
NOR2_X1 _17585_ ( .A1(_10854_ ), .A2(_10975_ ), .ZN(_00086_ ) );
OAI21_X1 _17586_ ( .A(_10965_ ), .B1(_10852_ ), .B2(\arbiter.clink.mtime [6] ), .ZN(_10976_ ) );
NOR2_X1 _17587_ ( .A1(_10853_ ), .A2(_10976_ ), .ZN(_00087_ ) );
OAI21_X1 _17588_ ( .A(_10965_ ), .B1(_10851_ ), .B2(\arbiter.clink.mtime [5] ), .ZN(_10977_ ) );
NOR2_X1 _17589_ ( .A1(_10852_ ), .A2(_10977_ ), .ZN(_00088_ ) );
OAI21_X1 _17590_ ( .A(_10965_ ), .B1(_10850_ ), .B2(\arbiter.clink.mtime [4] ), .ZN(_10978_ ) );
NOR2_X1 _17591_ ( .A1(_10851_ ), .A2(_10978_ ), .ZN(_00089_ ) );
BUF_X4 _17592_ ( .A(_10846_ ), .Z(_10979_ ) );
OAI21_X1 _17593_ ( .A(_10979_ ), .B1(_10903_ ), .B2(\arbiter.clink.mtime [57] ), .ZN(_10980_ ) );
NOR2_X1 _17594_ ( .A1(_10967_ ), .A2(_10980_ ), .ZN(_00090_ ) );
OAI21_X1 _17595_ ( .A(_10979_ ), .B1(_10849_ ), .B2(\arbiter.clink.mtime [3] ), .ZN(_10981_ ) );
NOR2_X1 _17596_ ( .A1(_10850_ ), .A2(_10981_ ), .ZN(_00091_ ) );
OAI21_X1 _17597_ ( .A(_10979_ ), .B1(_10848_ ), .B2(\arbiter.clink.mtime [2] ), .ZN(_10982_ ) );
NOR2_X1 _17598_ ( .A1(_10849_ ), .A2(_10982_ ), .ZN(_00092_ ) );
NOR2_X1 _17599_ ( .A1(\arbiter.clink.mtime [1] ), .A2(\arbiter.clink.mtime [0] ), .ZN(_10983_ ) );
NOR3_X1 _17600_ ( .A1(_10848_ ), .A2(_10983_ ), .A3(fanout_net_19 ), .ZN(_00093_ ) );
CLKBUF_X2 _17601_ ( .A(_10846_ ), .Z(\ifu.ren_REG_$_DFF_P__Q_D_$_NAND__Y_B ) );
AND2_X1 _17602_ ( .A1(\ifu.ren_REG_$_DFF_P__Q_D_$_NAND__Y_B ), .A2(\arbiter.clink._mtime_T_1 [0] ), .ZN(_00094_ ) );
OAI21_X1 _17603_ ( .A(_10979_ ), .B1(_10902_ ), .B2(\arbiter.clink.mtime [56] ), .ZN(_10984_ ) );
NOR2_X1 _17604_ ( .A1(_10903_ ), .A2(_10984_ ), .ZN(_00095_ ) );
OAI21_X1 _17605_ ( .A(_10979_ ), .B1(_10901_ ), .B2(\arbiter.clink.mtime [55] ), .ZN(_10985_ ) );
NOR2_X1 _17606_ ( .A1(_10902_ ), .A2(_10985_ ), .ZN(_00096_ ) );
OAI21_X1 _17607_ ( .A(_10979_ ), .B1(_10900_ ), .B2(\arbiter.clink.mtime [54] ), .ZN(_10986_ ) );
NOR2_X1 _17608_ ( .A1(_10901_ ), .A2(_10986_ ), .ZN(_00097_ ) );
CLKBUF_X2 _17609_ ( .A(_10846_ ), .Z(_10987_ ) );
AND3_X1 _17610_ ( .A1(_10987_ ), .A2(io_master_rlast ), .A3(io_master_rvalid ), .ZN(_00098_ ) );
INV_X1 _17611_ ( .A(fanout_net_1 ), .ZN(_10988_ ) );
BUF_X2 _17612_ ( .A(_10988_ ), .Z(_10989_ ) );
BUF_X2 _17613_ ( .A(_10989_ ), .Z(_10990_ ) );
AOI211_X1 _17614_ ( .A(fanout_net_19 ), .B(_10990_ ), .C1(_08564_ ), .C2(_08565_ ), .ZN(_00099_ ) );
INV_X1 _17615_ ( .A(_10826_ ), .ZN(_10991_ ) );
CLKBUF_X2 _17616_ ( .A(_10846_ ), .Z(_10992_ ) );
OAI211_X1 _17617_ ( .A(_10991_ ), .B(_10992_ ), .C1(\exu.io_in_valid ), .C2(\exu.state ), .ZN(_10993_ ) );
INV_X1 _17618_ ( .A(_10993_ ), .ZN(_00100_ ) );
NOR3_X1 _17619_ ( .A1(_10603_ ), .A2(_10637_ ), .A3(_10666_ ), .ZN(_10994_ ) );
AND2_X2 _17620_ ( .A1(_10673_ ), .A2(_10994_ ), .ZN(_10995_ ) );
AND2_X1 _17621_ ( .A1(_10995_ ), .A2(_10671_ ), .ZN(\idu.io_out_bits_xori ) );
AND2_X1 _17622_ ( .A1(_10669_ ), .A2(_10624_ ), .ZN(_10996_ ) );
AND2_X1 _17623_ ( .A1(_10995_ ), .A2(_10996_ ), .ZN(\idu.io_out_bits_slti ) );
OR2_X1 _17624_ ( .A1(\idu.io_out_bits_xori ), .A2(\idu.io_out_bits_slti ), .ZN(_10997_ ) );
AND2_X1 _17625_ ( .A1(_10673_ ), .A2(_10638_ ), .ZN(_10998_ ) );
AND2_X1 _17626_ ( .A1(_10998_ ), .A2(_10996_ ), .ZN(\idu.io_out_bits_lw ) );
AND3_X1 _17627_ ( .A1(_10668_ ), .A2(\idu.io_in_bits_inst [12] ), .A3(_10624_ ), .ZN(_10999_ ) );
AND2_X1 _17628_ ( .A1(_10995_ ), .A2(_10999_ ), .ZN(\idu.io_out_bits_sltiu ) );
NOR3_X1 _17629_ ( .A1(_10997_ ), .A2(\idu.io_out_bits_lw ), .A3(\idu.io_out_bits_sltiu ), .ZN(_11000_ ) );
CLKBUF_X2 _17630_ ( .A(_10673_ ), .Z(_11001_ ) );
OAI211_X1 _17631_ ( .A(_11001_ ), .B(_10638_ ), .C1(_10695_ ), .C2(_10634_ ), .ZN(_11002_ ) );
AOI22_X1 _17632_ ( .A1(_10671_ ), .A2(_10998_ ), .B1(_10995_ ), .B2(_10680_ ), .ZN(_11003_ ) );
INV_X1 _17633_ ( .A(\idu.io_out_bits_jalr ), .ZN(_11004_ ) );
OAI21_X1 _17634_ ( .A(_10995_ ), .B1(_10695_ ), .B2(_10670_ ), .ZN(_11005_ ) );
AND2_X1 _17635_ ( .A1(_11004_ ), .A2(_11005_ ), .ZN(_11006_ ) );
NAND4_X1 _17636_ ( .A1(_11000_ ), .A2(_11002_ ), .A3(_11003_ ), .A4(_11006_ ), .ZN(_11007_ ) );
NAND3_X1 _17637_ ( .A1(_10673_ ), .A2(_10611_ ), .A3(_10994_ ), .ZN(_11008_ ) );
INV_X1 _17638_ ( .A(_10581_ ), .ZN(_11009_ ) );
INV_X1 _17639_ ( .A(_10674_ ), .ZN(_11010_ ) );
NAND2_X1 _17640_ ( .A1(_10590_ ), .A2(_10586_ ), .ZN(_11011_ ) );
NOR4_X1 _17641_ ( .A1(_11008_ ), .A2(_11009_ ), .A3(_11010_ ), .A4(_11011_ ), .ZN(\idu.io_out_bits_srai ) );
AND3_X1 _17642_ ( .A1(_10657_ ), .A2(_10659_ ), .A3(_10681_ ), .ZN(\idu.io_out_bits_csrrw ) );
AND3_X1 _17643_ ( .A1(_10657_ ), .A2(_10659_ ), .A3(_10996_ ), .ZN(\idu.io_out_bits_csrrs ) );
NOR3_X1 _17644_ ( .A1(\idu.io_out_bits_srai ), .A2(\idu.io_out_bits_csrrw ), .A3(\idu.io_out_bits_csrrs ), .ZN(_11012_ ) );
AND4_X1 _17645_ ( .A1(_10653_ ), .A2(_10995_ ), .A3(_10654_ ), .A4(_10674_ ), .ZN(\idu.io_out_bits_srli ) );
INV_X1 _17646_ ( .A(\idu.io_out_bits_srli ), .ZN(_11013_ ) );
NAND2_X1 _17647_ ( .A1(_11012_ ), .A2(_11013_ ), .ZN(_11014_ ) );
NOR2_X1 _17648_ ( .A1(_11007_ ), .A2(_11014_ ), .ZN(_11015_ ) );
INV_X1 _17649_ ( .A(\idu.io_out_bits_jal ), .ZN(_11016_ ) );
AND2_X1 _17650_ ( .A1(_11015_ ), .A2(_11016_ ), .ZN(_11017_ ) );
AND4_X1 _17651_ ( .A1(_10636_ ), .A2(_10673_ ), .A3(_10667_ ), .A4(_10996_ ), .ZN(\idu.io_out_bits_sw ) );
AND4_X1 _17652_ ( .A1(_10636_ ), .A2(_10673_ ), .A3(_10667_ ), .A4(_10681_ ), .ZN(\idu.io_out_bits_sh ) );
OR2_X1 _17653_ ( .A1(\idu.io_out_bits_sw ), .A2(\idu.io_out_bits_sh ), .ZN(_11018_ ) );
AND4_X1 _17654_ ( .A1(_10636_ ), .A2(_10673_ ), .A3(_10695_ ), .A4(_10667_ ), .ZN(\idu.io_out_bits_sb ) );
NOR2_X1 _17655_ ( .A1(_11018_ ), .A2(\idu.io_out_bits_sb ), .ZN(_11019_ ) );
AND2_X1 _17656_ ( .A1(_11019_ ), .A2(_10683_ ), .ZN(_11020_ ) );
AND2_X2 _17657_ ( .A1(_11017_ ), .A2(_11020_ ), .ZN(_11021_ ) );
NOR2_X1 _17658_ ( .A1(_11015_ ), .A2(_10588_ ), .ZN(_11022_ ) );
NOR2_X1 _17659_ ( .A1(_11019_ ), .A2(_10588_ ), .ZN(_11023_ ) );
INV_X1 _17660_ ( .A(_11023_ ), .ZN(_11024_ ) );
AND3_X1 _17661_ ( .A1(_11001_ ), .A2(_10676_ ), .A3(_10680_ ), .ZN(\idu.io_out_bits_bgeu ) );
AND3_X1 _17662_ ( .A1(_11001_ ), .A2(_10695_ ), .A3(_10676_ ), .ZN(\idu.io_out_bits_beq ) );
AND3_X1 _17663_ ( .A1(_10673_ ), .A2(_10676_ ), .A3(_10674_ ), .ZN(\idu.io_out_bits_bge ) );
AND3_X1 _17664_ ( .A1(_10673_ ), .A2(_10676_ ), .A3(_10681_ ), .ZN(\idu.io_out_bits_bne ) );
OR4_X1 _17665_ ( .A1(\idu.io_out_bits_bgeu ), .A2(\idu.io_out_bits_beq ), .A3(\idu.io_out_bits_bge ), .A4(\idu.io_out_bits_bne ), .ZN(_11025_ ) );
AND3_X1 _17666_ ( .A1(_11001_ ), .A2(_10676_ ), .A3(_10670_ ), .ZN(\idu.io_out_bits_bltu ) );
AND3_X1 _17667_ ( .A1(_11001_ ), .A2(_10676_ ), .A3(_10671_ ), .ZN(\idu.io_out_bits_blt ) );
OR2_X1 _17668_ ( .A1(\idu.io_out_bits_bltu ), .A2(\idu.io_out_bits_blt ), .ZN(_11026_ ) );
OAI21_X1 _17669_ ( .A(\idu.immB [11] ), .B1(_11025_ ), .B2(_11026_ ), .ZN(_11027_ ) );
INV_X1 _17670_ ( .A(\idu.immI [0] ), .ZN(_11028_ ) );
OAI211_X1 _17671_ ( .A(_11024_ ), .B(_11027_ ), .C1(_11028_ ), .C2(_11016_ ), .ZN(_11029_ ) );
OR2_X1 _17672_ ( .A1(_11022_ ), .A2(_11029_ ), .ZN(\idu.io_out_bits_imm [11] ) );
BUF_X4 _17673_ ( .A(_10646_ ), .Z(_11030_ ) );
NAND3_X1 _17674_ ( .A1(_11030_ ), .A2(\idu.io_in_bits_inst [28] ), .A3(\idu.io_in_bits_inst [29] ), .ZN(_11031_ ) );
NOR4_X1 _17675_ ( .A1(_11021_ ), .A2(\idu.io_out_bits_imm [11] ), .A3(_10590_ ), .A4(_11031_ ), .ZN(_11032_ ) );
INV_X1 _17676_ ( .A(_11022_ ), .ZN(_11033_ ) );
OAI21_X1 _17677_ ( .A(_10587_ ), .B1(_11025_ ), .B2(_11026_ ), .ZN(_11034_ ) );
AND2_X2 _17678_ ( .A1(_11024_ ), .A2(_11034_ ), .ZN(_11035_ ) );
AND3_X1 _17679_ ( .A1(_10658_ ), .A2(\idu.io_in_bits_inst [4] ), .A3(_10636_ ), .ZN(_11036_ ) );
AND2_X2 _17680_ ( .A1(_10694_ ), .A2(_11036_ ), .ZN(\idu.io_out_bits_lui ) );
AND2_X2 _17681_ ( .A1(_10694_ ), .A2(_10994_ ), .ZN(\idu.io_out_bits_auipc ) );
NOR2_X1 _17682_ ( .A1(\idu.io_out_bits_lui ), .A2(\idu.io_out_bits_auipc ), .ZN(_11037_ ) );
AND2_X1 _17683_ ( .A1(_11016_ ), .A2(_11037_ ), .ZN(_11038_ ) );
INV_X1 _17684_ ( .A(_11038_ ), .ZN(_11039_ ) );
NAND3_X1 _17685_ ( .A1(_11039_ ), .A2(\idu.io_in_bits_inst [15] ), .A3(_11030_ ), .ZN(_11040_ ) );
NAND3_X1 _17686_ ( .A1(_11033_ ), .A2(_11035_ ), .A3(_11040_ ), .ZN(\idu.io_out_bits_imm [15] ) );
INV_X1 _17687_ ( .A(_10668_ ), .ZN(_11041_ ) );
OR2_X1 _17688_ ( .A1(_11038_ ), .A2(_11041_ ), .ZN(_11042_ ) );
NAND3_X1 _17689_ ( .A1(_11033_ ), .A2(_11035_ ), .A3(_11042_ ), .ZN(\idu.io_out_bits_imm [13] ) );
NAND2_X1 _17690_ ( .A1(_11039_ ), .A2(_10632_ ), .ZN(_11043_ ) );
OR2_X1 _17691_ ( .A1(_11038_ ), .A2(_10626_ ), .ZN(_11044_ ) );
NAND3_X1 _17692_ ( .A1(_11024_ ), .A2(_11043_ ), .A3(_11044_ ), .ZN(_11045_ ) );
NOR3_X1 _17693_ ( .A1(\idu.io_out_bits_imm [15] ), .A2(\idu.io_out_bits_imm [13] ), .A3(_11045_ ), .ZN(_11046_ ) );
AND2_X2 _17694_ ( .A1(_11032_ ), .A2(_11046_ ), .ZN(_11047_ ) );
AOI21_X1 _17695_ ( .A(_11021_ ), .B1(_10581_ ), .B2(_10583_ ), .ZN(_11048_ ) );
CLKBUF_X2 _17696_ ( .A(_10621_ ), .Z(_11049_ ) );
BUF_X2 _17697_ ( .A(_11049_ ), .Z(_11050_ ) );
CLKBUF_X2 _17698_ ( .A(_11050_ ), .Z(_11051_ ) );
BUF_X2 _17699_ ( .A(_11051_ ), .Z(_11052_ ) );
AOI21_X1 _17700_ ( .A(_11052_ ), .B1(_11015_ ), .B2(_11016_ ), .ZN(_11053_ ) );
INV_X1 _17701_ ( .A(_11020_ ), .ZN(_11054_ ) );
AND2_X1 _17702_ ( .A1(_11054_ ), .A2(\idu.immB [4] ), .ZN(_11055_ ) );
OR2_X1 _17703_ ( .A1(_11053_ ), .A2(_11055_ ), .ZN(\idu.io_out_bits_imm [4] ) );
NOR2_X1 _17704_ ( .A1(_11048_ ), .A2(\idu.io_out_bits_imm [4] ), .ZN(_11056_ ) );
AND2_X2 _17705_ ( .A1(_10684_ ), .A2(_10623_ ), .ZN(_11057_ ) );
NOR2_X1 _17706_ ( .A1(\idu.io_out_bits_csrrw ), .A2(\idu.io_out_bits_csrrs ), .ZN(_11058_ ) );
INV_X1 _17707_ ( .A(_11058_ ), .ZN(_11059_ ) );
NOR2_X1 _17708_ ( .A1(_11057_ ), .A2(_11059_ ), .ZN(_11060_ ) );
INV_X1 _17709_ ( .A(_11060_ ), .ZN(\idu.io_out_bits_wen_csr ) );
INV_X1 _17710_ ( .A(\idu.immB [3] ), .ZN(_11061_ ) );
INV_X1 _17711_ ( .A(\idu.immI [3] ), .ZN(_11062_ ) );
OAI221_X1 _17712_ ( .A(\idu.io_out_bits_wen_csr ), .B1(_11061_ ), .B2(_11020_ ), .C1(_11017_ ), .C2(_11062_ ), .ZN(_11063_ ) );
AOI211_X1 _17713_ ( .A(_10640_ ), .B(_10760_ ), .C1(_11019_ ), .C2(_10683_ ), .ZN(_11064_ ) );
INV_X1 _17714_ ( .A(_11017_ ), .ZN(_11065_ ) );
AOI21_X1 _17715_ ( .A(_11064_ ), .B1(_11065_ ), .B2(\idu.immI [2] ), .ZN(_11066_ ) );
INV_X1 _17716_ ( .A(\idu.immI [1] ), .ZN(_11067_ ) );
NOR2_X1 _17717_ ( .A1(_11015_ ), .A2(_11067_ ), .ZN(_11068_ ) );
OR2_X1 _17718_ ( .A1(\idu.io_out_bits_beq ), .A2(\idu.io_out_bits_bne ), .ZN(_11069_ ) );
OR4_X1 _17719_ ( .A1(\idu.io_out_bits_blt ), .A2(_11069_ ), .A3(\idu.io_out_bits_bgeu ), .A4(\idu.io_out_bits_bge ), .ZN(_11070_ ) );
OAI21_X1 _17720_ ( .A(\idu.immB [1] ), .B1(_11070_ ), .B2(\idu.io_out_bits_bltu ), .ZN(_11071_ ) );
OAI21_X1 _17721_ ( .A(\idu.immB [1] ), .B1(_11018_ ), .B2(\idu.io_out_bits_sb ), .ZN(_11072_ ) );
OAI211_X1 _17722_ ( .A(_11071_ ), .B(_11072_ ), .C1(_11067_ ), .C2(_11016_ ), .ZN(_11073_ ) );
NOR2_X1 _17723_ ( .A1(_11068_ ), .A2(_11073_ ), .ZN(_11074_ ) );
INV_X1 _17724_ ( .A(_11074_ ), .ZN(\idu.io_out_bits_imm [1] ) );
OAI21_X1 _17725_ ( .A(\idu.immI [0] ), .B1(_11007_ ), .B2(_11014_ ), .ZN(_11075_ ) );
OAI21_X1 _17726_ ( .A(\idu.immB [11] ), .B1(_11018_ ), .B2(\idu.io_out_bits_sb ), .ZN(_11076_ ) );
AND2_X1 _17727_ ( .A1(_11075_ ), .A2(_11076_ ), .ZN(_11077_ ) );
NOR4_X1 _17728_ ( .A1(_11063_ ), .A2(_11066_ ), .A3(\idu.io_out_bits_imm [1] ), .A4(_11077_ ), .ZN(_11078_ ) );
AND3_X1 _17729_ ( .A1(_11047_ ), .A2(_11056_ ), .A3(_11078_ ), .ZN(_11079_ ) );
NOR2_X1 _17730_ ( .A1(_11079_ ), .A2(_11057_ ), .ZN(_11080_ ) );
NOR2_X1 _17731_ ( .A1(_11021_ ), .A2(_10591_ ), .ZN(\idu.io_out_bits_imm [10] ) );
AND3_X1 _17732_ ( .A1(\idu.io_out_bits_imm [10] ), .A2(\idu.io_out_bits_imm [11] ), .A3(\idu.io_out_bits_imm [4] ), .ZN(_11081_ ) );
BUF_X4 _17733_ ( .A(_10760_ ), .Z(_11082_ ) );
NOR3_X1 _17734_ ( .A1(_11021_ ), .A2(_10609_ ), .A3(_11082_ ), .ZN(\idu.io_out_bits_imm [8] ) );
AOI211_X1 _17735_ ( .A(_10607_ ), .B(_11082_ ), .C1(_11017_ ), .C2(_11020_ ), .ZN(\idu.io_out_bits_imm [9] ) );
NAND3_X1 _17736_ ( .A1(_11081_ ), .A2(\idu.io_out_bits_imm [8] ), .A3(\idu.io_out_bits_imm [9] ), .ZN(_11083_ ) );
NOR2_X1 _17737_ ( .A1(_11083_ ), .A2(_11048_ ), .ZN(_11084_ ) );
AOI21_X1 _17738_ ( .A(_11061_ ), .B1(_11019_ ), .B2(_10683_ ), .ZN(_11085_ ) );
AOI21_X1 _17739_ ( .A(_11085_ ), .B1(_11065_ ), .B2(\idu.immI [3] ), .ZN(_11086_ ) );
AND2_X1 _17740_ ( .A1(_11066_ ), .A2(_11086_ ), .ZN(_11087_ ) );
AND4_X1 _17741_ ( .A1(\idu.io_out_bits_imm [1] ), .A2(_11087_ ), .A3(_11077_ ), .A4(\idu.io_out_bits_wen_csr ), .ZN(_11088_ ) );
OAI21_X1 _17742_ ( .A(_10608_ ), .B1(\idu.io_out_bits_lui ), .B2(\idu.io_out_bits_auipc ), .ZN(_11089_ ) );
AND2_X1 _17743_ ( .A1(\idu.io_out_bits_jal ), .A2(_10587_ ), .ZN(_11090_ ) );
INV_X1 _17744_ ( .A(_11090_ ), .ZN(_11091_ ) );
AND3_X1 _17745_ ( .A1(_11034_ ), .A2(_11089_ ), .A3(_11091_ ), .ZN(_11092_ ) );
AND3_X1 _17746_ ( .A1(_11033_ ), .A2(_11024_ ), .A3(_11092_ ), .ZN(_11093_ ) );
NOR3_X1 _17747_ ( .A1(_11068_ ), .A2(_11073_ ), .A3(_11060_ ), .ZN(_11094_ ) );
INV_X1 _17748_ ( .A(_11035_ ), .ZN(_11095_ ) );
INV_X1 _17749_ ( .A(_10605_ ), .ZN(_11096_ ) );
CLKBUF_X2 _17750_ ( .A(_11096_ ), .Z(_11097_ ) );
BUF_X2 _17751_ ( .A(_11097_ ), .Z(_11098_ ) );
BUF_X2 _17752_ ( .A(_11098_ ), .Z(_11099_ ) );
BUF_X2 _17753_ ( .A(_11099_ ), .Z(_11100_ ) );
BUF_X2 _17754_ ( .A(_11100_ ), .Z(_11101_ ) );
AOI21_X1 _17755_ ( .A(_11101_ ), .B1(_11016_ ), .B2(_11037_ ), .ZN(_11102_ ) );
NOR3_X1 _17756_ ( .A1(_11022_ ), .A2(_11095_ ), .A3(_11102_ ), .ZN(_11103_ ) );
AND3_X1 _17757_ ( .A1(_11093_ ), .A2(_11094_ ), .A3(_11103_ ), .ZN(_11104_ ) );
OAI21_X1 _17758_ ( .A(_11035_ ), .B1(_10595_ ), .B2(_11038_ ), .ZN(_11105_ ) );
INV_X1 _17759_ ( .A(_11105_ ), .ZN(_11106_ ) );
BUF_X2 _17760_ ( .A(_11024_ ), .Z(_11107_ ) );
OAI21_X1 _17761_ ( .A(_10580_ ), .B1(\idu.io_out_bits_lui ), .B2(\idu.io_out_bits_auipc ), .ZN(_11108_ ) );
OAI21_X1 _17762_ ( .A(_10610_ ), .B1(\idu.io_out_bits_lui ), .B2(\idu.io_out_bits_auipc ), .ZN(_11109_ ) );
OAI21_X1 _17763_ ( .A(\idu.funct7 [0] ), .B1(\idu.io_out_bits_lui ), .B2(\idu.io_out_bits_auipc ), .ZN(_11110_ ) );
AND3_X1 _17764_ ( .A1(_11024_ ), .A2(_11109_ ), .A3(_11110_ ), .ZN(_11111_ ) );
AND4_X1 _17765_ ( .A1(_11107_ ), .A2(_11077_ ), .A3(_11108_ ), .A4(_11111_ ), .ZN(_11112_ ) );
AND4_X2 _17766_ ( .A1(_11104_ ), .A2(_11087_ ), .A3(_11106_ ), .A4(_11112_ ), .ZN(_11113_ ) );
AND3_X1 _17767_ ( .A1(_11056_ ), .A2(_11046_ ), .A3(_11032_ ), .ZN(_11114_ ) );
AOI22_X1 _17768_ ( .A1(_11084_ ), .A2(_11088_ ), .B1(_11113_ ), .B2(_11114_ ), .ZN(_11115_ ) );
AND2_X2 _17769_ ( .A1(_11080_ ), .A2(_11115_ ), .ZN(_11116_ ) );
BUF_X4 _17770_ ( .A(_11116_ ), .Z(_11117_ ) );
BUF_X4 _17771_ ( .A(_11117_ ), .Z(_11118_ ) );
NOR3_X1 _17772_ ( .A1(_11031_ ), .A2(_10587_ ), .A3(_10590_ ), .ZN(_11119_ ) );
NAND3_X1 _17773_ ( .A1(_10606_ ), .A2(_10584_ ), .A3(_11119_ ), .ZN(_11120_ ) );
CLKBUF_X2 _17774_ ( .A(_10620_ ), .Z(_11121_ ) );
BUF_X2 _17775_ ( .A(_11121_ ), .Z(_11122_ ) );
BUF_X2 _17776_ ( .A(_11122_ ), .Z(_11123_ ) );
BUF_X2 _17777_ ( .A(_11123_ ), .Z(_11124_ ) );
BUF_X2 _17778_ ( .A(_11124_ ), .Z(_11125_ ) );
INV_X1 _17779_ ( .A(_10686_ ), .ZN(_11126_ ) );
CLKBUF_X2 _17780_ ( .A(_11126_ ), .Z(_11127_ ) );
NOR3_X1 _17781_ ( .A1(_11120_ ), .A2(_11125_ ), .A3(_11127_ ), .ZN(_11128_ ) );
AND3_X2 _17782_ ( .A1(_10663_ ), .A2(_11128_ ), .A3(_10660_ ), .ZN(_11129_ ) );
BUF_X2 _17783_ ( .A(_11129_ ), .Z(\idu._io_csr_raddr_T_15 [1] ) );
INV_X1 _17784_ ( .A(_11079_ ), .ZN(_11130_ ) );
INV_X1 _17785_ ( .A(_10578_ ), .ZN(_11131_ ) );
NAND3_X1 _17786_ ( .A1(\idu.io_out_bits_wen_csr ), .A2(_10582_ ), .A3(_11131_ ), .ZN(_11132_ ) );
OR3_X1 _17787_ ( .A1(_11053_ ), .A2(_11055_ ), .A3(_11132_ ), .ZN(_11133_ ) );
INV_X1 _17788_ ( .A(_10580_ ), .ZN(_11134_ ) );
NOR3_X1 _17789_ ( .A1(_11133_ ), .A2(_11134_ ), .A3(_11021_ ), .ZN(_11135_ ) );
NOR3_X1 _17790_ ( .A1(_11077_ ), .A2(_11073_ ), .A3(_11068_ ), .ZN(_11136_ ) );
AND3_X1 _17791_ ( .A1(_11087_ ), .A2(_11135_ ), .A3(_11136_ ), .ZN(_11137_ ) );
NAND2_X1 _17792_ ( .A1(_11137_ ), .A2(_11047_ ), .ZN(_11138_ ) );
INV_X1 _17793_ ( .A(_11057_ ), .ZN(_11139_ ) );
NAND3_X1 _17794_ ( .A1(_11130_ ), .A2(_11138_ ), .A3(_11139_ ), .ZN(_11140_ ) );
BUF_X2 _17795_ ( .A(_11140_ ), .Z(\idu._io_out_bits_csr_waddr_T_16 [1] ) );
OAI211_X1 _17796_ ( .A(_11118_ ), .B(\wbu.csr_2 [30] ), .C1(\idu._io_csr_raddr_T_15 [1] ), .C2(\idu._io_out_bits_csr_waddr_T_16 [1] ), .ZN(_11141_ ) );
BUF_X4 _17797_ ( .A(_11084_ ), .Z(_11142_ ) );
AND3_X2 _17798_ ( .A1(_11087_ ), .A2(_11136_ ), .A3(\idu.io_out_bits_wen_csr ), .ZN(_11143_ ) );
BUF_X4 _17799_ ( .A(_11143_ ), .Z(_11144_ ) );
NAND3_X1 _17800_ ( .A1(_11056_ ), .A2(_11046_ ), .A3(_11032_ ), .ZN(_11145_ ) );
NAND4_X1 _17801_ ( .A1(_11104_ ), .A2(_11087_ ), .A3(_11106_ ), .A4(_11112_ ), .ZN(_11146_ ) );
NOR2_X1 _17802_ ( .A1(_11145_ ), .A2(_11146_ ), .ZN(_11147_ ) );
BUF_X4 _17803_ ( .A(_11147_ ), .Z(_11148_ ) );
AOI22_X1 _17804_ ( .A1(_11142_ ), .A2(_11144_ ), .B1(_11148_ ), .B2(\wbu._GEN_135 [30] ), .ZN(_11149_ ) );
BUF_X4 _17805_ ( .A(_11079_ ), .Z(_11150_ ) );
BUF_X4 _17806_ ( .A(_11150_ ), .Z(_11151_ ) );
BUF_X4 _17807_ ( .A(_11057_ ), .Z(_11152_ ) );
BUF_X4 _17808_ ( .A(_11152_ ), .Z(_11153_ ) );
OAI21_X1 _17809_ ( .A(\wbu.csr_3 [30] ), .B1(_11151_ ), .B2(_11153_ ), .ZN(_11154_ ) );
AND2_X1 _17810_ ( .A1(_11149_ ), .A2(_11154_ ), .ZN(_11155_ ) );
NAND2_X1 _17811_ ( .A1(_11141_ ), .A2(_11155_ ), .ZN(_00101_ ) );
OAI211_X1 _17812_ ( .A(_11118_ ), .B(\wbu.csr_2 [28] ), .C1(\idu._io_csr_raddr_T_15 [1] ), .C2(\idu._io_out_bits_csr_waddr_T_16 [1] ), .ZN(_11156_ ) );
BUF_X4 _17813_ ( .A(_11084_ ), .Z(_11157_ ) );
AOI22_X1 _17814_ ( .A1(_11157_ ), .A2(_11144_ ), .B1(_11148_ ), .B2(\wbu._GEN_135 [28] ), .ZN(_11158_ ) );
OAI21_X1 _17815_ ( .A(\wbu.csr_3 [28] ), .B1(_11150_ ), .B2(_11152_ ), .ZN(_11159_ ) );
AND2_X1 _17816_ ( .A1(_11158_ ), .A2(_11159_ ), .ZN(_11160_ ) );
NAND2_X1 _17817_ ( .A1(_11156_ ), .A2(_11160_ ), .ZN(_00102_ ) );
BUF_X4 _17818_ ( .A(_11116_ ), .Z(_11161_ ) );
BUF_X4 _17819_ ( .A(_11129_ ), .Z(_11162_ ) );
BUF_X4 _17820_ ( .A(_11140_ ), .Z(_11163_ ) );
OAI211_X1 _17821_ ( .A(_11161_ ), .B(\wbu.csr_2 [12] ), .C1(_11162_ ), .C2(_11163_ ), .ZN(_11164_ ) );
BUF_X2 _17822_ ( .A(_11150_ ), .Z(_11165_ ) );
BUF_X2 _17823_ ( .A(_11152_ ), .Z(\idu._io_csr_raddr_T_14 [0] ) );
OAI21_X1 _17824_ ( .A(\wbu.csr_3 [12] ), .B1(_11165_ ), .B2(\idu._io_csr_raddr_T_14 [0] ), .ZN(_11166_ ) );
BUF_X2 _17825_ ( .A(_11148_ ), .Z(_11167_ ) );
AOI22_X1 _17826_ ( .A1(_11142_ ), .A2(_11144_ ), .B1(_11167_ ), .B2(\wbu._GEN_135 [12] ), .ZN(_11168_ ) );
NAND3_X1 _17827_ ( .A1(_11164_ ), .A2(_11166_ ), .A3(_11168_ ), .ZN(_00103_ ) );
OAI211_X1 _17828_ ( .A(_11118_ ), .B(\wbu.csr_2 [11] ), .C1(\idu._io_csr_raddr_T_15 [1] ), .C2(\idu._io_out_bits_csr_waddr_T_16 [1] ), .ZN(_11169_ ) );
AOI22_X1 _17829_ ( .A1(_11157_ ), .A2(_11144_ ), .B1(_11148_ ), .B2(\wbu._GEN_135 [11] ), .ZN(_11170_ ) );
OAI21_X1 _17830_ ( .A(\wbu.csr_3 [11] ), .B1(_11150_ ), .B2(_11152_ ), .ZN(_11171_ ) );
AND2_X1 _17831_ ( .A1(_11170_ ), .A2(_11171_ ), .ZN(_11172_ ) );
NAND2_X1 _17832_ ( .A1(_11169_ ), .A2(_11172_ ), .ZN(_00104_ ) );
OAI211_X1 _17833_ ( .A(_11117_ ), .B(\wbu.csr_2 [8] ), .C1(_11162_ ), .C2(_11163_ ), .ZN(_11173_ ) );
OAI21_X1 _17834_ ( .A(\wbu.csr_3 [8] ), .B1(_11165_ ), .B2(\idu._io_csr_raddr_T_14 [0] ), .ZN(_11174_ ) );
AOI22_X1 _17835_ ( .A1(_11142_ ), .A2(_11144_ ), .B1(_11167_ ), .B2(\wbu._GEN_135 [8] ), .ZN(_11175_ ) );
NAND3_X1 _17836_ ( .A1(_11173_ ), .A2(_11174_ ), .A3(_11175_ ), .ZN(_00105_ ) );
OAI211_X1 _17837_ ( .A(_11118_ ), .B(\wbu.csr_2 [6] ), .C1(\idu._io_csr_raddr_T_15 [1] ), .C2(\idu._io_out_bits_csr_waddr_T_16 [1] ), .ZN(_11176_ ) );
AOI22_X1 _17838_ ( .A1(_11157_ ), .A2(_11144_ ), .B1(_11148_ ), .B2(\wbu._GEN_135 [6] ), .ZN(_11177_ ) );
OAI21_X1 _17839_ ( .A(\wbu.csr_3 [6] ), .B1(_11150_ ), .B2(_11152_ ), .ZN(_11178_ ) );
AND2_X1 _17840_ ( .A1(_11177_ ), .A2(_11178_ ), .ZN(_11179_ ) );
NAND2_X1 _17841_ ( .A1(_11176_ ), .A2(_11179_ ), .ZN(_00106_ ) );
OAI211_X1 _17842_ ( .A(_11117_ ), .B(\wbu.csr_2 [4] ), .C1(_11162_ ), .C2(_11163_ ), .ZN(_11180_ ) );
OAI21_X1 _17843_ ( .A(\wbu.csr_3 [4] ), .B1(_11165_ ), .B2(\idu._io_csr_raddr_T_14 [0] ), .ZN(_11181_ ) );
AOI22_X1 _17844_ ( .A1(_11142_ ), .A2(_11144_ ), .B1(_11167_ ), .B2(\wbu._GEN_135 [4] ), .ZN(_11182_ ) );
NAND3_X1 _17845_ ( .A1(_11180_ ), .A2(_11181_ ), .A3(_11182_ ), .ZN(_00107_ ) );
NAND2_X1 _17846_ ( .A1(_11084_ ), .A2(_11088_ ), .ZN(_11183_ ) );
INV_X1 _17847_ ( .A(_11183_ ), .ZN(_11184_ ) );
AND2_X1 _17848_ ( .A1(_11137_ ), .A2(_11047_ ), .ZN(_11185_ ) );
NOR4_X1 _17849_ ( .A1(_11079_ ), .A2(_11185_ ), .A3(_11057_ ), .A4(_11129_ ), .ZN(_11186_ ) );
INV_X1 _17850_ ( .A(_11186_ ), .ZN(_11187_ ) );
AND2_X1 _17851_ ( .A1(_11187_ ), .A2(_11116_ ), .ZN(_11188_ ) );
INV_X1 _17852_ ( .A(_11147_ ), .ZN(_11189_ ) );
NAND2_X1 _17853_ ( .A1(_11189_ ), .A2(\wbu.csr_0 [0] ), .ZN(_11190_ ) );
BUF_X4 _17854_ ( .A(_11113_ ), .Z(_11191_ ) );
BUF_X4 _17855_ ( .A(_11047_ ), .Z(_11192_ ) );
BUF_X4 _17856_ ( .A(_11056_ ), .Z(_11193_ ) );
NAND4_X1 _17857_ ( .A1(_11191_ ), .A2(\wbu._GEN_135 [3] ), .A3(_11192_ ), .A4(_11193_ ), .ZN(_11194_ ) );
AOI21_X1 _17858_ ( .A(_11188_ ), .B1(_11190_ ), .B2(_11194_ ), .ZN(_11195_ ) );
AND4_X1 _17859_ ( .A1(\wbu.csr_2 [3] ), .A2(_11187_ ), .A3(_11080_ ), .A4(_11115_ ), .ZN(_11196_ ) );
OAI21_X1 _17860_ ( .A(_11080_ ), .B1(_11195_ ), .B2(_11196_ ), .ZN(_11197_ ) );
AND2_X1 _17861_ ( .A1(_11157_ ), .A2(_11143_ ), .ZN(_11198_ ) );
INV_X1 _17862_ ( .A(_11080_ ), .ZN(_11199_ ) );
AOI21_X1 _17863_ ( .A(_11198_ ), .B1(_11199_ ), .B2(\wbu.csr_3 [3] ), .ZN(_11200_ ) );
AOI21_X1 _17864_ ( .A(_11184_ ), .B1(_11197_ ), .B2(_11200_ ), .ZN(_00108_ ) );
NAND4_X1 _17865_ ( .A1(_11113_ ), .A2(\wbu._GEN_135 [29] ), .A3(_11047_ ), .A4(_11056_ ), .ZN(_11201_ ) );
INV_X1 _17866_ ( .A(_11157_ ), .ZN(_11202_ ) );
INV_X1 _17867_ ( .A(_11143_ ), .ZN(_11203_ ) );
OAI211_X1 _17868_ ( .A(_11183_ ), .B(_11201_ ), .C1(_11202_ ), .C2(_11203_ ), .ZN(_11204_ ) );
AOI21_X1 _17869_ ( .A(_11204_ ), .B1(\wbu.csr_3 [29] ), .B2(_11199_ ), .ZN(_11205_ ) );
BUF_X4 _17870_ ( .A(_11129_ ), .Z(_11206_ ) );
BUF_X4 _17871_ ( .A(_11140_ ), .Z(_11207_ ) );
OAI211_X1 _17872_ ( .A(_11161_ ), .B(\wbu.csr_2 [29] ), .C1(_11206_ ), .C2(_11207_ ), .ZN(_11208_ ) );
NAND2_X1 _17873_ ( .A1(_11205_ ), .A2(_11208_ ), .ZN(_00109_ ) );
OAI211_X1 _17874_ ( .A(_11117_ ), .B(\wbu.csr_2 [26] ), .C1(_11162_ ), .C2(_11163_ ), .ZN(_11209_ ) );
OAI21_X1 _17875_ ( .A(\wbu.csr_3 [26] ), .B1(_11165_ ), .B2(\idu._io_csr_raddr_T_14 [0] ), .ZN(_11210_ ) );
AOI22_X1 _17876_ ( .A1(_11142_ ), .A2(_11088_ ), .B1(_11167_ ), .B2(\wbu._GEN_135 [26] ), .ZN(_11211_ ) );
NAND3_X1 _17877_ ( .A1(_11209_ ), .A2(_11210_ ), .A3(_11211_ ), .ZN(_00110_ ) );
NAND4_X1 _17878_ ( .A1(_11113_ ), .A2(\wbu._GEN_135 [24] ), .A3(_11047_ ), .A4(_11056_ ), .ZN(_11212_ ) );
OAI211_X1 _17879_ ( .A(_11183_ ), .B(_11212_ ), .C1(_11202_ ), .C2(_11203_ ), .ZN(_11213_ ) );
AOI21_X1 _17880_ ( .A(_11213_ ), .B1(\wbu.csr_3 [24] ), .B2(_11199_ ), .ZN(_11214_ ) );
OAI211_X1 _17881_ ( .A(_11161_ ), .B(\wbu.csr_2 [24] ), .C1(_11206_ ), .C2(_11207_ ), .ZN(_11215_ ) );
NAND2_X1 _17882_ ( .A1(_11214_ ), .A2(_11215_ ), .ZN(_00111_ ) );
OAI211_X1 _17883_ ( .A(_11117_ ), .B(\wbu.csr_2 [19] ), .C1(_11162_ ), .C2(_11163_ ), .ZN(_11216_ ) );
OAI21_X1 _17884_ ( .A(\wbu.csr_3 [19] ), .B1(_11165_ ), .B2(\idu._io_csr_raddr_T_14 [0] ), .ZN(_11217_ ) );
AOI22_X1 _17885_ ( .A1(_11142_ ), .A2(_11088_ ), .B1(_11167_ ), .B2(\wbu._GEN_135 [19] ), .ZN(_11218_ ) );
NAND3_X1 _17886_ ( .A1(_11216_ ), .A2(_11217_ ), .A3(_11218_ ), .ZN(_00112_ ) );
OAI211_X1 _17887_ ( .A(_11117_ ), .B(\wbu.csr_2 [27] ), .C1(_11162_ ), .C2(_11163_ ), .ZN(_11219_ ) );
OAI21_X1 _17888_ ( .A(\wbu.csr_3 [27] ), .B1(_11165_ ), .B2(\idu._io_csr_raddr_T_14 [0] ), .ZN(_11220_ ) );
AOI22_X1 _17889_ ( .A1(_11142_ ), .A2(_11144_ ), .B1(_11167_ ), .B2(\wbu._GEN_135 [27] ), .ZN(_11221_ ) );
NAND3_X1 _17890_ ( .A1(_11219_ ), .A2(_11220_ ), .A3(_11221_ ), .ZN(_00113_ ) );
OAI211_X1 _17891_ ( .A(_11117_ ), .B(\wbu.csr_2 [9] ), .C1(_11162_ ), .C2(_11163_ ), .ZN(_11222_ ) );
OAI21_X1 _17892_ ( .A(\wbu.csr_3 [9] ), .B1(_11165_ ), .B2(\idu._io_csr_raddr_T_14 [0] ), .ZN(_11223_ ) );
AOI22_X1 _17893_ ( .A1(_11142_ ), .A2(_11088_ ), .B1(_11167_ ), .B2(\wbu._GEN_135 [9] ), .ZN(_11224_ ) );
NAND3_X1 _17894_ ( .A1(_11222_ ), .A2(_11223_ ), .A3(_11224_ ), .ZN(_00114_ ) );
OAI211_X1 _17895_ ( .A(_11117_ ), .B(\wbu.csr_2 [5] ), .C1(_11162_ ), .C2(_11163_ ), .ZN(_11225_ ) );
OAI21_X1 _17896_ ( .A(\wbu.csr_3 [5] ), .B1(_11165_ ), .B2(\idu._io_csr_raddr_T_14 [0] ), .ZN(_11226_ ) );
AND3_X1 _17897_ ( .A1(_11114_ ), .A2(\wbu._GEN_135 [5] ), .A3(_11113_ ), .ZN(_11227_ ) );
NOR3_X1 _17898_ ( .A1(_11184_ ), .A2(_11198_ ), .A3(_11227_ ), .ZN(_11228_ ) );
NAND3_X1 _17899_ ( .A1(_11225_ ), .A2(_11226_ ), .A3(_11228_ ), .ZN(_00115_ ) );
INV_X1 _17900_ ( .A(\wbu.csr_3 [1] ), .ZN(_11229_ ) );
AOI21_X1 _17901_ ( .A(_11229_ ), .B1(_11130_ ), .B2(_11139_ ), .ZN(_11230_ ) );
NAND4_X1 _17902_ ( .A1(_11113_ ), .A2(\wbu._GEN_135 [1] ), .A3(_11047_ ), .A4(_11056_ ), .ZN(_11231_ ) );
NAND2_X1 _17903_ ( .A1(_11190_ ), .A2(_11231_ ), .ZN(_11232_ ) );
MUX2_X1 _17904_ ( .A(_11232_ ), .B(\wbu.csr_2 [1] ), .S(_11188_ ), .Z(_11233_ ) );
AOI21_X1 _17905_ ( .A(_11230_ ), .B1(_11233_ ), .B2(_11080_ ), .ZN(_11234_ ) );
OAI21_X1 _17906_ ( .A(_11183_ ), .B1(_11234_ ), .B2(_11198_ ), .ZN(_00116_ ) );
OAI211_X1 _17907_ ( .A(_11118_ ), .B(\wbu.csr_2 [31] ), .C1(\idu._io_csr_raddr_T_15 [1] ), .C2(\idu._io_out_bits_csr_waddr_T_16 [1] ), .ZN(_11235_ ) );
OAI21_X1 _17908_ ( .A(\wbu.csr_3 [31] ), .B1(_11151_ ), .B2(_11153_ ), .ZN(_11236_ ) );
NAND4_X1 _17909_ ( .A1(_11191_ ), .A2(\wbu._GEN_135 [31] ), .A3(_11192_ ), .A4(_11193_ ), .ZN(_11237_ ) );
AND2_X1 _17910_ ( .A1(_11236_ ), .A2(_11237_ ), .ZN(_11238_ ) );
NAND2_X1 _17911_ ( .A1(_11235_ ), .A2(_11238_ ), .ZN(_00117_ ) );
OAI211_X1 _17912_ ( .A(_11118_ ), .B(\wbu.csr_2 [25] ), .C1(\idu._io_csr_raddr_T_15 [1] ), .C2(\idu._io_out_bits_csr_waddr_T_16 [1] ), .ZN(_11239_ ) );
OAI21_X1 _17913_ ( .A(\wbu.csr_3 [25] ), .B1(_11151_ ), .B2(_11153_ ), .ZN(_11240_ ) );
NAND4_X1 _17914_ ( .A1(_11191_ ), .A2(\wbu._GEN_135 [25] ), .A3(_11192_ ), .A4(_11193_ ), .ZN(_11241_ ) );
AND2_X1 _17915_ ( .A1(_11240_ ), .A2(_11241_ ), .ZN(_11242_ ) );
NAND2_X1 _17916_ ( .A1(_11239_ ), .A2(_11242_ ), .ZN(_00118_ ) );
OAI211_X1 _17917_ ( .A(_11118_ ), .B(\wbu.csr_2 [23] ), .C1(\idu._io_csr_raddr_T_15 [1] ), .C2(\idu._io_out_bits_csr_waddr_T_16 [1] ), .ZN(_11243_ ) );
OAI21_X1 _17918_ ( .A(\wbu.csr_3 [23] ), .B1(_11151_ ), .B2(_11153_ ), .ZN(_11244_ ) );
NAND4_X1 _17919_ ( .A1(_11191_ ), .A2(\wbu._GEN_135 [23] ), .A3(_11192_ ), .A4(_11193_ ), .ZN(_11245_ ) );
AND2_X1 _17920_ ( .A1(_11244_ ), .A2(_11245_ ), .ZN(_11246_ ) );
NAND2_X1 _17921_ ( .A1(_11243_ ), .A2(_11246_ ), .ZN(_00119_ ) );
OAI211_X1 _17922_ ( .A(_11118_ ), .B(\wbu.csr_2 [18] ), .C1(\idu._io_csr_raddr_T_15 [1] ), .C2(\idu._io_out_bits_csr_waddr_T_16 [1] ), .ZN(_11247_ ) );
OAI21_X1 _17923_ ( .A(\wbu.csr_3 [18] ), .B1(_11151_ ), .B2(_11153_ ), .ZN(_11248_ ) );
NAND4_X1 _17924_ ( .A1(_11191_ ), .A2(\wbu._GEN_135 [18] ), .A3(_11192_ ), .A4(_11193_ ), .ZN(_11249_ ) );
AND2_X1 _17925_ ( .A1(_11248_ ), .A2(_11249_ ), .ZN(_11250_ ) );
NAND2_X1 _17926_ ( .A1(_11247_ ), .A2(_11250_ ), .ZN(_00120_ ) );
OAI211_X1 _17927_ ( .A(_11118_ ), .B(\wbu.csr_2 [15] ), .C1(\idu._io_csr_raddr_T_15 [1] ), .C2(\idu._io_out_bits_csr_waddr_T_16 [1] ), .ZN(_11251_ ) );
OAI21_X1 _17928_ ( .A(\wbu.csr_3 [15] ), .B1(_11151_ ), .B2(_11153_ ), .ZN(_11252_ ) );
NAND4_X1 _17929_ ( .A1(_11191_ ), .A2(\wbu._GEN_135 [15] ), .A3(_11192_ ), .A4(_11193_ ), .ZN(_11253_ ) );
AND2_X1 _17930_ ( .A1(_11252_ ), .A2(_11253_ ), .ZN(_11254_ ) );
NAND2_X1 _17931_ ( .A1(_11251_ ), .A2(_11254_ ), .ZN(_00121_ ) );
OAI211_X1 _17932_ ( .A(_11118_ ), .B(\wbu.csr_2 [10] ), .C1(_11206_ ), .C2(_11207_ ), .ZN(_11255_ ) );
OAI21_X1 _17933_ ( .A(\wbu.csr_3 [10] ), .B1(_11151_ ), .B2(_11153_ ), .ZN(_11256_ ) );
NAND4_X1 _17934_ ( .A1(_11191_ ), .A2(\wbu._GEN_135 [10] ), .A3(_11192_ ), .A4(_11193_ ), .ZN(_11257_ ) );
AND2_X1 _17935_ ( .A1(_11256_ ), .A2(_11257_ ), .ZN(_11258_ ) );
NAND2_X1 _17936_ ( .A1(_11255_ ), .A2(_11258_ ), .ZN(_00122_ ) );
OAI211_X1 _17937_ ( .A(_11161_ ), .B(\wbu.csr_2 [7] ), .C1(_11206_ ), .C2(_11207_ ), .ZN(_11259_ ) );
OAI21_X1 _17938_ ( .A(\wbu.csr_3 [7] ), .B1(_11151_ ), .B2(_11153_ ), .ZN(_11260_ ) );
NAND4_X1 _17939_ ( .A1(_11191_ ), .A2(\wbu._GEN_135 [7] ), .A3(_11192_ ), .A4(_11193_ ), .ZN(_11261_ ) );
AND2_X1 _17940_ ( .A1(_11260_ ), .A2(_11261_ ), .ZN(_11262_ ) );
NAND2_X1 _17941_ ( .A1(_11259_ ), .A2(_11262_ ), .ZN(_00123_ ) );
OAI211_X1 _17942_ ( .A(_11161_ ), .B(\wbu.csr_2 [22] ), .C1(_11206_ ), .C2(_11207_ ), .ZN(_11263_ ) );
AOI22_X1 _17943_ ( .A1(_11157_ ), .A2(_11143_ ), .B1(_11148_ ), .B2(\wbu._GEN_135 [22] ), .ZN(_11264_ ) );
OAI21_X1 _17944_ ( .A(\wbu.csr_3 [22] ), .B1(_11150_ ), .B2(_11152_ ), .ZN(_11265_ ) );
AND2_X1 _17945_ ( .A1(_11264_ ), .A2(_11265_ ), .ZN(_11266_ ) );
NAND2_X1 _17946_ ( .A1(_11263_ ), .A2(_11266_ ), .ZN(_00124_ ) );
OAI211_X1 _17947_ ( .A(_11161_ ), .B(\wbu.csr_2 [2] ), .C1(_11206_ ), .C2(_11207_ ), .ZN(_11267_ ) );
OAI21_X1 _17948_ ( .A(\wbu.csr_3 [2] ), .B1(_11151_ ), .B2(_11153_ ), .ZN(_11268_ ) );
NAND4_X1 _17949_ ( .A1(_11191_ ), .A2(\wbu._GEN_135 [2] ), .A3(_11192_ ), .A4(_11193_ ), .ZN(_11269_ ) );
AND2_X1 _17950_ ( .A1(_11268_ ), .A2(_11269_ ), .ZN(_11270_ ) );
NAND2_X1 _17951_ ( .A1(_11267_ ), .A2(_11270_ ), .ZN(_00125_ ) );
OAI221_X1 _17952_ ( .A(_11183_ ), .B1(_11202_ ), .B2(_11203_ ), .C1(_11080_ ), .C2(\wbu.csr_3 [0] ), .ZN(_11271_ ) );
INV_X1 _17953_ ( .A(_11116_ ), .ZN(_11272_ ) );
OR3_X1 _17954_ ( .A1(_11272_ ), .A2(_11186_ ), .A3(\wbu.csr_2 [0] ), .ZN(_11273_ ) );
NAND4_X1 _17955_ ( .A1(_11191_ ), .A2(\wbu._GEN_135 [0] ), .A3(_11192_ ), .A4(_11193_ ), .ZN(_11274_ ) );
NAND2_X1 _17956_ ( .A1(_11190_ ), .A2(_11274_ ), .ZN(_11275_ ) );
OAI21_X1 _17957_ ( .A(_11273_ ), .B1(_11188_ ), .B2(_11275_ ), .ZN(_11276_ ) );
AOI21_X1 _17958_ ( .A(_11271_ ), .B1(_11276_ ), .B2(_11080_ ), .ZN(_00126_ ) );
OAI211_X1 _17959_ ( .A(_11161_ ), .B(\wbu.csr_2 [21] ), .C1(_11206_ ), .C2(_11207_ ), .ZN(_11277_ ) );
AOI22_X1 _17960_ ( .A1(_11157_ ), .A2(_11143_ ), .B1(_11148_ ), .B2(\wbu._GEN_135 [21] ), .ZN(_11278_ ) );
OAI21_X1 _17961_ ( .A(\wbu.csr_3 [21] ), .B1(_11150_ ), .B2(_11152_ ), .ZN(_11279_ ) );
AND2_X1 _17962_ ( .A1(_11278_ ), .A2(_11279_ ), .ZN(_11280_ ) );
NAND2_X1 _17963_ ( .A1(_11277_ ), .A2(_11280_ ), .ZN(_00127_ ) );
OAI211_X1 _17964_ ( .A(_11161_ ), .B(\wbu.csr_2 [20] ), .C1(_11206_ ), .C2(_11207_ ), .ZN(_11281_ ) );
AOI22_X1 _17965_ ( .A1(_11157_ ), .A2(_11143_ ), .B1(_11148_ ), .B2(\wbu._GEN_135 [20] ), .ZN(_11282_ ) );
OAI21_X1 _17966_ ( .A(\wbu.csr_3 [20] ), .B1(_11150_ ), .B2(_11152_ ), .ZN(_11283_ ) );
AND2_X1 _17967_ ( .A1(_11282_ ), .A2(_11283_ ), .ZN(_11284_ ) );
NAND2_X1 _17968_ ( .A1(_11281_ ), .A2(_11284_ ), .ZN(_00128_ ) );
OAI211_X1 _17969_ ( .A(_11161_ ), .B(\wbu.csr_2 [17] ), .C1(_11206_ ), .C2(_11207_ ), .ZN(_11285_ ) );
AOI22_X1 _17970_ ( .A1(_11157_ ), .A2(_11143_ ), .B1(_11148_ ), .B2(\wbu._GEN_135 [17] ), .ZN(_11286_ ) );
OAI21_X1 _17971_ ( .A(\wbu.csr_3 [17] ), .B1(_11150_ ), .B2(_11152_ ), .ZN(_11287_ ) );
AND2_X1 _17972_ ( .A1(_11286_ ), .A2(_11287_ ), .ZN(_11288_ ) );
NAND2_X1 _17973_ ( .A1(_11285_ ), .A2(_11288_ ), .ZN(_00129_ ) );
OAI211_X1 _17974_ ( .A(_11117_ ), .B(\wbu.csr_2 [16] ), .C1(_11162_ ), .C2(_11163_ ), .ZN(_11289_ ) );
OAI21_X1 _17975_ ( .A(\wbu.csr_3 [16] ), .B1(_11165_ ), .B2(\idu._io_csr_raddr_T_14 [0] ), .ZN(_11290_ ) );
AOI22_X1 _17976_ ( .A1(_11142_ ), .A2(_11144_ ), .B1(_11167_ ), .B2(\wbu._GEN_135 [16] ), .ZN(_11291_ ) );
NAND3_X1 _17977_ ( .A1(_11289_ ), .A2(_11290_ ), .A3(_11291_ ), .ZN(_00130_ ) );
OAI211_X1 _17978_ ( .A(_11161_ ), .B(\wbu.csr_2 [14] ), .C1(_11206_ ), .C2(_11207_ ), .ZN(_11292_ ) );
AOI22_X1 _17979_ ( .A1(_11157_ ), .A2(_11143_ ), .B1(_11148_ ), .B2(\wbu._GEN_135 [14] ), .ZN(_11293_ ) );
OAI21_X1 _17980_ ( .A(\wbu.csr_3 [14] ), .B1(_11150_ ), .B2(_11152_ ), .ZN(_11294_ ) );
AND2_X1 _17981_ ( .A1(_11293_ ), .A2(_11294_ ), .ZN(_11295_ ) );
NAND2_X1 _17982_ ( .A1(_11292_ ), .A2(_11295_ ), .ZN(_00131_ ) );
OAI211_X1 _17983_ ( .A(_11117_ ), .B(\wbu.csr_2 [13] ), .C1(_11162_ ), .C2(_11163_ ), .ZN(_11296_ ) );
OAI21_X1 _17984_ ( .A(\wbu.csr_3 [13] ), .B1(_11151_ ), .B2(_11153_ ), .ZN(_11297_ ) );
AOI22_X1 _17985_ ( .A1(_11142_ ), .A2(_11144_ ), .B1(_11167_ ), .B2(\wbu._GEN_135 [13] ), .ZN(_11298_ ) );
NAND3_X1 _17986_ ( .A1(_11296_ ), .A2(_11297_ ), .A3(_11298_ ), .ZN(_00132_ ) );
AND3_X1 _17987_ ( .A1(fanout_net_2 ), .A2(\icache._icache_reg_T ), .A3(io_master_rvalid ), .ZN(_11299_ ) );
INV_X1 _17988_ ( .A(_11299_ ), .ZN(_11300_ ) );
BUF_X4 _17989_ ( .A(_11300_ ), .Z(_11301_ ) );
AND3_X1 _17990_ ( .A1(_09399_ ), .A2(_09466_ ), .A3(_09403_ ), .ZN(_11302_ ) );
INV_X1 _17991_ ( .A(_09650_ ), .ZN(_11303_ ) );
AND2_X1 _17992_ ( .A1(_09330_ ), .A2(_09331_ ), .ZN(_11304_ ) );
AND2_X1 _17993_ ( .A1(_09468_ ), .A2(_09469_ ), .ZN(_11305_ ) );
AND3_X1 _17994_ ( .A1(_09404_ ), .A2(_11305_ ), .A3(_09405_ ), .ZN(_11306_ ) );
NAND3_X1 _17995_ ( .A1(_09189_ ), .A2(_11304_ ), .A3(_11306_ ), .ZN(_11307_ ) );
INV_X1 _17996_ ( .A(_09523_ ), .ZN(_11308_ ) );
AOI21_X1 _17997_ ( .A(_09611_ ), .B1(_09561_ ), .B2(_09562_ ), .ZN(_11309_ ) );
AOI211_X1 _17998_ ( .A(_11303_ ), .B(_11307_ ), .C1(_11308_ ), .C2(_11309_ ), .ZN(_11310_ ) );
AOI211_X1 _17999_ ( .A(_11302_ ), .B(_11310_ ), .C1(\ifu.pc [28] ), .C2(\ifu._start_T ), .ZN(_11311_ ) );
AND2_X1 _18000_ ( .A1(_09816_ ), .A2(_09817_ ), .ZN(_11312_ ) );
AND3_X1 _18001_ ( .A1(_09715_ ), .A2(_09716_ ), .A3(_11312_ ), .ZN(_11313_ ) );
AND3_X1 _18002_ ( .A1(_11308_ ), .A2(_09650_ ), .A3(_11309_ ), .ZN(_11314_ ) );
AND3_X1 _18003_ ( .A1(_09189_ ), .A2(_11304_ ), .A3(_11306_ ), .ZN(_11315_ ) );
AND2_X1 _18004_ ( .A1(_09869_ ), .A2(_09918_ ), .ZN(_11316_ ) );
NAND3_X1 _18005_ ( .A1(_11316_ ), .A2(_10153_ ), .A3(_10202_ ), .ZN(_11317_ ) );
AOI22_X1 _18006_ ( .A1(_10102_ ), .A2(_10103_ ), .B1(_10010_ ), .B2(_10012_ ), .ZN(_11318_ ) );
NAND3_X1 _18007_ ( .A1(_09969_ ), .A2(_10057_ ), .A3(_11318_ ), .ZN(_11319_ ) );
OAI211_X1 _18008_ ( .A(_11314_ ), .B(_11315_ ), .C1(_11317_ ), .C2(_11319_ ), .ZN(_11320_ ) );
NAND4_X1 _18009_ ( .A1(_11311_ ), .A2(_09772_ ), .A3(_11313_ ), .A4(_11320_ ), .ZN(_11321_ ) );
AND4_X1 _18010_ ( .A1(_09772_ ), .A2(_11313_ ), .A3(_10834_ ), .A4(_11315_ ), .ZN(_11322_ ) );
AND4_X1 _18011_ ( .A1(_09969_ ), .A2(_11314_ ), .A3(_10057_ ), .A4(_11318_ ), .ZN(_11323_ ) );
NAND4_X1 _18012_ ( .A1(_11316_ ), .A2(_10153_ ), .A3(_10199_ ), .A4(_10201_ ), .ZN(_11324_ ) );
AOI21_X1 _18013_ ( .A(_10433_ ), .B1(_10473_ ), .B2(_10474_ ), .ZN(_11325_ ) );
INV_X1 _18014_ ( .A(_10561_ ), .ZN(_11326_ ) );
INV_X1 _18015_ ( .A(_10520_ ), .ZN(_11327_ ) );
AND3_X1 _18016_ ( .A1(_11325_ ), .A2(_11326_ ), .A3(_11327_ ), .ZN(_11328_ ) );
AOI21_X1 _18017_ ( .A(_08788_ ), .B1(_08786_ ), .B2(_08591_ ), .ZN(_11329_ ) );
XOR2_X1 _18018_ ( .A(_08587_ ), .B(_08588_ ), .Z(_11330_ ) );
INV_X1 _18019_ ( .A(_11330_ ), .ZN(_11331_ ) );
NAND3_X1 _18020_ ( .A1(_08781_ ), .A2(_08783_ ), .A3(_11331_ ), .ZN(_11332_ ) );
INV_X1 _18021_ ( .A(_08781_ ), .ZN(_11333_ ) );
NAND3_X1 _18022_ ( .A1(_11333_ ), .A2(_08813_ ), .A3(_11330_ ), .ZN(_11334_ ) );
AND3_X1 _18023_ ( .A1(_09944_ ), .A2(_08923_ ), .A3(_11330_ ), .ZN(_11335_ ) );
AND2_X1 _18024_ ( .A1(fanout_net_19 ), .A2(\exu.auipc.io_rs1_data [1] ), .ZN(_11336_ ) );
INV_X1 _18025_ ( .A(_11336_ ), .ZN(_11337_ ) );
NAND2_X1 _18026_ ( .A1(_09190_ ), .A2(\exu.csrrs.io_csr_rdata [1] ), .ZN(_11338_ ) );
AOI21_X1 _18027_ ( .A(_09211_ ), .B1(_11337_ ), .B2(_11338_ ), .ZN(_11339_ ) );
NOR3_X1 _18028_ ( .A1(_08591_ ), .A2(\exu.io_in_bits_mret ), .A3(\exu.io_in_bits_en_dnpc ), .ZN(_11340_ ) );
OAI21_X1 _18029_ ( .A(_09254_ ), .B1(_11339_ ), .B2(_11340_ ), .ZN(_11341_ ) );
MUX2_X1 _18030_ ( .A(_08591_ ), .B(_11331_ ), .S(_08945_ ), .Z(_11342_ ) );
OAI211_X1 _18031_ ( .A(_09222_ ), .B(_11341_ ), .C1(_11342_ ), .C2(_09255_ ), .ZN(_11343_ ) );
AOI22_X1 _18032_ ( .A1(_08977_ ), .A2(_08591_ ), .B1(_08979_ ), .B2(_11331_ ), .ZN(_11344_ ) );
OAI211_X1 _18033_ ( .A(_09412_ ), .B(_11343_ ), .C1(_11344_ ), .C2(_09252_ ), .ZN(_11345_ ) );
MUX2_X1 _18034_ ( .A(_08591_ ), .B(_11331_ ), .S(_08935_ ), .Z(_11346_ ) );
OAI21_X1 _18035_ ( .A(_11345_ ), .B1(_09413_ ), .B2(_11346_ ), .ZN(_11347_ ) );
AOI221_X4 _18036_ ( .A(_11335_ ), .B1(\exu.auipc.io_rs1_data [1] ), .B2(_08928_ ), .C1(_11347_ ), .C2(_09250_ ), .ZN(_11348_ ) );
OAI221_X1 _18037_ ( .A(_11334_ ), .B1(_08591_ ), .B2(_09309_ ), .C1(_11348_ ), .C2(\exu.bne.io_is ), .ZN(_11349_ ) );
AOI221_X4 _18038_ ( .A(\exu.io_in_bits_jal ), .B1(_11329_ ), .B2(_11332_ ), .C1(_11349_ ), .C2(_09249_ ), .ZN(_11350_ ) );
AOI211_X1 _18039_ ( .A(_08702_ ), .B(_11336_ ), .C1(_11330_ ), .C2(_09396_ ), .ZN(_11351_ ) );
OR3_X1 _18040_ ( .A1(_11350_ ), .A2(fanout_net_8 ), .A3(_11351_ ), .ZN(_11352_ ) );
NAND3_X1 _18041_ ( .A1(_09462_ ), .A2(fanout_net_8 ), .A3(\exu.csrrs.io_csr_rdata [1] ), .ZN(_11353_ ) );
NAND3_X1 _18042_ ( .A1(_11352_ ), .A2(_09321_ ), .A3(_11353_ ), .ZN(_11354_ ) );
INV_X1 _18043_ ( .A(_09055_ ), .ZN(_11355_ ) );
NAND3_X1 _18044_ ( .A1(_09052_ ), .A2(_09054_ ), .A3(_11355_ ), .ZN(_11356_ ) );
OAI21_X1 _18045_ ( .A(_09053_ ), .B1(_09051_ ), .B2(_09055_ ), .ZN(_11357_ ) );
NAND2_X1 _18046_ ( .A1(_11356_ ), .A2(_11357_ ), .ZN(_11358_ ) );
AOI21_X1 _18047_ ( .A(_11336_ ), .B1(_11358_ ), .B2(_09396_ ), .ZN(_11359_ ) );
AOI211_X1 _18048_ ( .A(exu_io_in_valid_REG_$_NOT__A_Y ), .B(_09401_ ), .C1(\exu.io_in_bits_jalr ), .C2(_11359_ ), .ZN(_11360_ ) );
NAND2_X1 _18049_ ( .A1(_11354_ ), .A2(_11360_ ), .ZN(_11361_ ) );
OAI21_X1 _18050_ ( .A(\ifu._pc_T_8 [1] ), .B1(_09401_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_11362_ ) );
NAND3_X1 _18051_ ( .A1(_11361_ ), .A2(_09182_ ), .A3(_11362_ ), .ZN(_11363_ ) );
OR2_X1 _18052_ ( .A1(_09182_ ), .A2(\ifu._pc_T_8 [1] ), .ZN(_11364_ ) );
NAND2_X1 _18053_ ( .A1(_11363_ ), .A2(_11364_ ), .ZN(_11365_ ) );
XOR2_X1 _18054_ ( .A(\exu.addi.io_imm [0] ), .B(\exu.auipc.io_rs1_data [0] ), .Z(_11366_ ) );
NOR3_X1 _18055_ ( .A1(_08781_ ), .A2(_08814_ ), .A3(_11366_ ), .ZN(_11367_ ) );
INV_X1 _18056_ ( .A(_11366_ ), .ZN(_11368_ ) );
AOI211_X1 _18057_ ( .A(_08933_ ), .B(_11368_ ), .C1(_08866_ ), .C2(_08917_ ), .ZN(_11369_ ) );
OAI21_X1 _18058_ ( .A(\exu.bgeu.io_is ), .B1(_09437_ ), .B2(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_11370_ ) );
AND3_X1 _18059_ ( .A1(_08920_ ), .A2(_08975_ ), .A3(_11366_ ), .ZN(_11371_ ) );
INV_X1 _18060_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_11372_ ) );
AOI211_X1 _18061_ ( .A(_09252_ ), .B(_11371_ ), .C1(_09432_ ), .C2(_11372_ ), .ZN(_11373_ ) );
AND2_X1 _18062_ ( .A1(_09191_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_11374_ ) );
AND2_X1 _18063_ ( .A1(fanout_net_19 ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_11375_ ) );
OR3_X1 _18064_ ( .A1(_11374_ ), .A2(_09288_ ), .A3(_11375_ ), .ZN(_11376_ ) );
INV_X1 _18065_ ( .A(\exu.auipc.io_rs1_data [0] ), .ZN(_11377_ ) );
OR3_X1 _18066_ ( .A1(_11377_ ), .A2(\exu.io_in_bits_mret ), .A3(\exu.io_in_bits_en_dnpc ), .ZN(_11378_ ) );
NAND3_X1 _18067_ ( .A1(_11376_ ), .A2(_09256_ ), .A3(_11378_ ), .ZN(_11379_ ) );
MUX2_X1 _18068_ ( .A(_11372_ ), .B(_11366_ ), .S(_08945_ ), .Z(_11380_ ) );
OAI21_X1 _18069_ ( .A(_11379_ ), .B1(_11380_ ), .B2(_09256_ ), .ZN(_11381_ ) );
AOI21_X1 _18070_ ( .A(_11373_ ), .B1(_09253_ ), .B2(_11381_ ), .ZN(_11382_ ) );
OAI221_X1 _18071_ ( .A(_09251_ ), .B1(_11369_ ), .B2(_11370_ ), .C1(_11382_ ), .C2(\exu.bgeu.io_is ), .ZN(_11383_ ) );
MUX2_X1 _18072_ ( .A(_11372_ ), .B(_11366_ ), .S(_09303_ ), .Z(_11384_ ) );
AOI21_X1 _18073_ ( .A(\exu.bne.io_is ), .B1(_11384_ ), .B2(\exu.bge.io_is ), .ZN(_11385_ ) );
AOI221_X4 _18074_ ( .A(_11367_ ), .B1(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_09444_ ), .C1(_11383_ ), .C2(_11385_ ), .ZN(_11386_ ) );
NOR2_X1 _18075_ ( .A1(_11386_ ), .A2(\exu.beq.io_is ), .ZN(_11387_ ) );
AND4_X1 _18076_ ( .A1(_09395_ ), .A2(_08781_ ), .A3(\exu.beq.io_is ), .A4(_11366_ ), .ZN(_11388_ ) );
AOI211_X1 _18077_ ( .A(_09249_ ), .B(_11388_ ), .C1(_11372_ ), .C2(_08786_ ), .ZN(_11389_ ) );
OAI21_X1 _18078_ ( .A(_09409_ ), .B1(_11387_ ), .B2(_11389_ ), .ZN(_11390_ ) );
OR2_X1 _18079_ ( .A1(_11366_ ), .A2(_09999_ ), .ZN(_11391_ ) );
NAND3_X1 _18080_ ( .A1(fanout_net_19 ), .A2(\exu.io_in_bits_jal ), .A3(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_11392_ ) );
NAND4_X1 _18081_ ( .A1(_11390_ ), .A2(_08989_ ), .A3(_11391_ ), .A4(_11392_ ), .ZN(_11393_ ) );
NAND3_X1 _18082_ ( .A1(_09462_ ), .A2(fanout_net_8 ), .A3(\exu.csrrs.io_csr_rdata [0] ), .ZN(_11394_ ) );
NAND3_X1 _18083_ ( .A1(_11393_ ), .A2(_09321_ ), .A3(_11394_ ), .ZN(_11395_ ) );
NOR2_X1 _18084_ ( .A1(\exu.addi.io_imm [0] ), .A2(\exu.add.io_rs1_data [0] ), .ZN(_11396_ ) );
NOR2_X2 _18085_ ( .A1(_09053_ ), .A2(_11396_ ), .ZN(_11397_ ) );
NOR2_X1 _18086_ ( .A1(_11397_ ), .A2(_09177_ ), .ZN(_11398_ ) );
AND3_X1 _18087_ ( .A1(fanout_net_19 ), .A2(\exu.io_in_bits_jalr ), .A3(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_11399_ ) );
NOR4_X1 _18088_ ( .A1(_09401_ ), .A2(exu_io_in_valid_REG_$_NOT__A_Y ), .A3(_11398_ ), .A4(_11399_ ), .ZN(_11400_ ) );
NAND2_X1 _18089_ ( .A1(_11395_ ), .A2(_11400_ ), .ZN(_11401_ ) );
OR2_X1 _18090_ ( .A1(_09185_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_B ), .ZN(_11402_ ) );
NAND3_X1 _18091_ ( .A1(_11401_ ), .A2(_09182_ ), .A3(_11402_ ), .ZN(_11403_ ) );
OAI21_X1 _18092_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_11404_ ) );
NAND2_X1 _18093_ ( .A1(_11403_ ), .A2(_11404_ ), .ZN(_11405_ ) );
NAND3_X1 _18094_ ( .A1(_09191_ ), .A2(fanout_net_8 ), .A3(\exu.csrrs.io_csr_rdata [2] ), .ZN(_11406_ ) );
MUX2_X1 _18095_ ( .A(\exu.csrrs.io_csr_rdata [2] ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_29_A_$_MUX__A_B ), .S(fanout_net_19 ), .Z(_11407_ ) );
NOR2_X1 _18096_ ( .A1(_11407_ ), .A2(_08949_ ), .ZN(_11408_ ) );
NOR3_X1 _18097_ ( .A1(\exu.io_in_bits_mret ), .A2(\exu.auipc.io_rs1_data [2] ), .A3(\exu.io_in_bits_en_dnpc ), .ZN(_11409_ ) );
NOR3_X1 _18098_ ( .A1(_11408_ ), .A2(\exu.bltu.io_is ), .A3(_11409_ ), .ZN(_11410_ ) );
XOR2_X1 _18099_ ( .A(_08592_ ), .B(_08593_ ), .Z(_11411_ ) );
INV_X1 _18100_ ( .A(_11411_ ), .ZN(_11412_ ) );
MUX2_X1 _18101_ ( .A(\exu.auipc.io_rs1_data [2] ), .B(_11412_ ), .S(_08943_ ), .Z(_11413_ ) );
AOI211_X1 _18102_ ( .A(\exu.blt.io_is ), .B(_11410_ ), .C1(_11413_ ), .C2(\exu.bltu.io_is ), .ZN(_11414_ ) );
OAI22_X1 _18103_ ( .A1(_09798_ ), .A2(_11412_ ), .B1(_08976_ ), .B2(\exu.auipc.io_rs1_data [2] ), .ZN(_11415_ ) );
AOI211_X1 _18104_ ( .A(\exu.bgeu.io_is ), .B(_11414_ ), .C1(\exu.blt.io_is ), .C2(_11415_ ), .ZN(_11416_ ) );
MUX2_X1 _18105_ ( .A(\exu.auipc.io_rs1_data [2] ), .B(_11412_ ), .S(_08934_ ), .Z(_11417_ ) );
AOI211_X1 _18106_ ( .A(\exu.bge.io_is ), .B(_11416_ ), .C1(\exu.bgeu.io_is ), .C2(_11417_ ), .ZN(_11418_ ) );
MUX2_X1 _18107_ ( .A(_09197_ ), .B(_11411_ ), .S(_08925_ ), .Z(_11419_ ) );
AOI211_X1 _18108_ ( .A(\exu.bne.io_is ), .B(_11418_ ), .C1(\exu.bge.io_is ), .C2(_11419_ ), .ZN(_11420_ ) );
NOR3_X1 _18109_ ( .A1(_08781_ ), .A2(_08814_ ), .A3(_11412_ ), .ZN(_11421_ ) );
AOI211_X1 _18110_ ( .A(_08812_ ), .B(_11421_ ), .C1(_09197_ ), .C2(_09202_ ), .ZN(_11422_ ) );
OAI21_X1 _18111_ ( .A(_08788_ ), .B1(_11420_ ), .B2(_11422_ ), .ZN(_11423_ ) );
NAND4_X1 _18112_ ( .A1(_08781_ ), .A2(_09190_ ), .A3(\exu.beq.io_is ), .A4(_11411_ ), .ZN(_11424_ ) );
OAI211_X1 _18113_ ( .A(\exu.beq.io_is ), .B(_11424_ ), .C1(_09231_ ), .C2(\exu.auipc.io_rs1_data [2] ), .ZN(_11425_ ) );
AOI21_X1 _18114_ ( .A(\exu.io_in_bits_jal ), .B1(_11423_ ), .B2(_11425_ ), .ZN(_11426_ ) );
NAND3_X1 _18115_ ( .A1(fanout_net_19 ), .A2(\exu.io_in_bits_jal ), .A3(\exu.addi._io_rd_T_4_$_NOT__Y_29_A_$_MUX__A_B ), .ZN(_11427_ ) );
OAI211_X1 _18116_ ( .A(_08989_ ), .B(_11427_ ), .C1(_11411_ ), .C2(_09902_ ), .ZN(_11428_ ) );
OAI211_X1 _18117_ ( .A(_09041_ ), .B(_11406_ ), .C1(_11426_ ), .C2(_11428_ ), .ZN(_11429_ ) );
XOR2_X1 _18118_ ( .A(_09056_ ), .B(_09059_ ), .Z(\exu.addi._io_rd_T_4 [2] ) );
NOR2_X1 _18119_ ( .A1(\exu.addi._io_rd_T_4 [2] ), .A2(_09176_ ), .ZN(_11430_ ) );
AND2_X1 _18120_ ( .A1(_09176_ ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_29_A_$_MUX__A_B ), .ZN(_11431_ ) );
OAI21_X1 _18121_ ( .A(\exu.io_in_bits_jalr ), .B1(_11430_ ), .B2(_11431_ ), .ZN(_11432_ ) );
NAND3_X1 _18122_ ( .A1(_11429_ ), .A2(_09184_ ), .A3(_11432_ ), .ZN(_11433_ ) );
OR2_X1 _18123_ ( .A1(_09038_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_15_A_$_MUX__Y_B ), .ZN(_11434_ ) );
NAND3_X1 _18124_ ( .A1(_11433_ ), .A2(_09181_ ), .A3(_11434_ ), .ZN(_11435_ ) );
OAI21_X1 _18125_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_15_A_$_MUX__Y_B ), .B1(fanout_net_14 ), .B2(fanout_net_15 ), .ZN(_11436_ ) );
AND2_X2 _18126_ ( .A1(_11435_ ), .A2(_11436_ ), .ZN(_11437_ ) );
NAND3_X1 _18127_ ( .A1(_09191_ ), .A2(fanout_net_8 ), .A3(\exu.csrrs.io_csr_rdata [3] ), .ZN(_11438_ ) );
NAND2_X1 _18128_ ( .A1(_08594_ ), .A2(_08595_ ), .ZN(_11439_ ) );
XNOR2_X1 _18129_ ( .A(\exu.auipc.io_rs1_data [3] ), .B(\exu.addi.io_imm [3] ), .ZN(_11440_ ) );
XNOR2_X1 _18130_ ( .A(_11439_ ), .B(_11440_ ), .ZN(_11441_ ) );
OR3_X1 _18131_ ( .A1(_09428_ ), .A2(_08933_ ), .A3(_11441_ ), .ZN(_11442_ ) );
XOR2_X1 _18132_ ( .A(\exu.auipc.io_rs1_data [3] ), .B(\exu.auipc.io_rs1_data [2] ), .Z(_11443_ ) );
OAI211_X1 _18133_ ( .A(_11442_ ), .B(\exu.bgeu.io_is ), .C1(_08935_ ), .C2(_11443_ ), .ZN(_11444_ ) );
NOR2_X1 _18134_ ( .A1(_10110_ ), .A2(_11441_ ), .ZN(_11445_ ) );
INV_X1 _18135_ ( .A(_11443_ ), .ZN(_11446_ ) );
OAI211_X1 _18136_ ( .A(\exu.blt.io_is ), .B(_11446_ ), .C1(_08921_ ), .C2(fanout_net_19 ), .ZN(_11447_ ) );
AOI211_X1 _18137_ ( .A(_08940_ ), .B(_11443_ ), .C1(_08918_ ), .C2(_09190_ ), .ZN(_11448_ ) );
OAI21_X1 _18138_ ( .A(_08949_ ), .B1(_11446_ ), .B2(_09035_ ), .ZN(_11449_ ) );
AND3_X1 _18139_ ( .A1(fanout_net_19 ), .A2(\exu.io_in_bits_mret ), .A3(\exu.addi._io_rd_T_4_$_NOT__Y_28_A_$_MUX__A_B ), .ZN(_11450_ ) );
XNOR2_X1 _18140_ ( .A(\exu.csrrs.io_csr_rdata [3] ), .B(\exu.csrrs.io_csr_rdata [2] ), .ZN(_11451_ ) );
AOI21_X1 _18141_ ( .A(_11450_ ), .B1(_11451_ ), .B2(_08972_ ), .ZN(_11452_ ) );
AOI21_X1 _18142_ ( .A(\exu.bltu.io_is ), .B1(_11449_ ), .B2(_11452_ ), .ZN(_11453_ ) );
OAI21_X1 _18143_ ( .A(_08947_ ), .B1(_11448_ ), .B2(_11453_ ), .ZN(_11454_ ) );
NAND3_X1 _18144_ ( .A1(_11447_ ), .A2(_08931_ ), .A3(_11454_ ), .ZN(_11455_ ) );
OAI211_X1 _18145_ ( .A(_08922_ ), .B(_11444_ ), .C1(_11445_ ), .C2(_11455_ ), .ZN(_11456_ ) );
MUX2_X1 _18146_ ( .A(_11443_ ), .B(_11441_ ), .S(_08925_ ), .Z(_11457_ ) );
OAI211_X1 _18147_ ( .A(_11456_ ), .B(_08812_ ), .C1(_08922_ ), .C2(_11457_ ), .ZN(_11458_ ) );
INV_X1 _18148_ ( .A(_11441_ ), .ZN(_11459_ ) );
NAND3_X1 _18149_ ( .A1(_11333_ ), .A2(_08813_ ), .A3(_11459_ ), .ZN(_11460_ ) );
OAI211_X1 _18150_ ( .A(_11460_ ), .B(\exu.bne.io_is ), .C1(_08815_ ), .C2(_11443_ ), .ZN(_11461_ ) );
NAND3_X1 _18151_ ( .A1(_11458_ ), .A2(_08788_ ), .A3(_11461_ ), .ZN(_11462_ ) );
NAND4_X1 _18152_ ( .A1(_08781_ ), .A2(_09190_ ), .A3(\exu.beq.io_is ), .A4(_11441_ ), .ZN(_11463_ ) );
OAI211_X1 _18153_ ( .A(\exu.beq.io_is ), .B(_11463_ ), .C1(_09231_ ), .C2(_11446_ ), .ZN(_11464_ ) );
AOI21_X1 _18154_ ( .A(\exu.io_in_bits_jal ), .B1(_11462_ ), .B2(_11464_ ), .ZN(_11465_ ) );
NAND3_X1 _18155_ ( .A1(fanout_net_19 ), .A2(\exu.io_in_bits_jal ), .A3(\exu.addi._io_rd_T_4_$_NOT__Y_28_A_$_MUX__A_B ), .ZN(_11466_ ) );
OAI211_X1 _18156_ ( .A(_08988_ ), .B(_11466_ ), .C1(_11441_ ), .C2(_09902_ ), .ZN(_11467_ ) );
OAI211_X1 _18157_ ( .A(_09041_ ), .B(_11438_ ), .C1(_11465_ ), .C2(_11467_ ), .ZN(_11468_ ) );
AND3_X1 _18158_ ( .A1(fanout_net_19 ), .A2(\exu.io_in_bits_jalr ), .A3(\exu.addi._io_rd_T_4_$_NOT__Y_28_A_$_MUX__A_B ), .ZN(_11469_ ) );
AND2_X1 _18159_ ( .A1(_09060_ ), .A2(_09063_ ), .ZN(_11470_ ) );
NOR2_X1 _18160_ ( .A1(_09061_ ), .A2(_09065_ ), .ZN(_11471_ ) );
INV_X1 _18161_ ( .A(_11471_ ), .ZN(_11472_ ) );
XNOR2_X1 _18162_ ( .A(_11470_ ), .B(_11472_ ), .ZN(_11473_ ) );
AOI21_X1 _18163_ ( .A(_11469_ ), .B1(_11473_ ), .B2(_09173_ ), .ZN(_11474_ ) );
NAND3_X1 _18164_ ( .A1(_11468_ ), .A2(_09184_ ), .A3(_11474_ ), .ZN(_11475_ ) );
OR2_X1 _18165_ ( .A1(_09184_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_14_A_$_MUX__Y_B ), .ZN(_11476_ ) );
NAND3_X1 _18166_ ( .A1(_11475_ ), .A2(_09181_ ), .A3(_11476_ ), .ZN(_11477_ ) );
OAI21_X1 _18167_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_14_A_$_MUX__Y_B ), .B1(\ifu.start [0] ), .B2(\ifu.start [1] ), .ZN(_11478_ ) );
AND2_X2 _18168_ ( .A1(_11477_ ), .A2(_11478_ ), .ZN(_11479_ ) );
NOR2_X1 _18169_ ( .A1(_11437_ ), .A2(_11479_ ), .ZN(_11480_ ) );
NAND4_X1 _18170_ ( .A1(_11328_ ), .A2(_11365_ ), .A3(_11405_ ), .A4(_11480_ ), .ZN(_11481_ ) );
INV_X1 _18171_ ( .A(_10299_ ), .ZN(_11482_ ) );
INV_X1 _18172_ ( .A(_10390_ ), .ZN(_11483_ ) );
INV_X1 _18173_ ( .A(_10250_ ), .ZN(_11484_ ) );
NAND4_X1 _18174_ ( .A1(_11482_ ), .A2(_11483_ ), .A3(_11484_ ), .A4(_10349_ ), .ZN(_11485_ ) );
NOR3_X1 _18175_ ( .A1(_11324_ ), .A2(_11481_ ), .A3(_11485_ ), .ZN(_11486_ ) );
NAND3_X1 _18176_ ( .A1(_11322_ ), .A2(_11323_ ), .A3(_11486_ ), .ZN(_11487_ ) );
NAND2_X1 _18177_ ( .A1(_11321_ ), .A2(_11487_ ), .ZN(_11488_ ) );
BUF_X4 _18178_ ( .A(_11488_ ), .Z(_11489_ ) );
AND3_X1 _18179_ ( .A1(_09715_ ), .A2(_09772_ ), .A3(_09716_ ), .ZN(_11490_ ) );
NAND4_X1 _18180_ ( .A1(_09189_ ), .A2(_11305_ ), .A3(_11304_ ), .A4(_09650_ ), .ZN(_11491_ ) );
NAND4_X1 _18181_ ( .A1(_11490_ ), .A2(_11312_ ), .A3(_09406_ ), .A4(_11491_ ), .ZN(_11492_ ) );
BUF_X4 _18182_ ( .A(_11492_ ), .Z(_11493_ ) );
AOI211_X1 _18183_ ( .A(\io_master_rdata [31] ), .B(_11301_ ), .C1(_11489_ ), .C2(_11493_ ), .ZN(_11494_ ) );
AND2_X2 _18184_ ( .A1(_11488_ ), .A2(_11492_ ), .ZN(_11495_ ) );
INV_X1 _18185_ ( .A(_11495_ ), .ZN(_11496_ ) );
BUF_X4 _18186_ ( .A(_11299_ ), .Z(_11497_ ) );
AND2_X1 _18187_ ( .A1(_11496_ ), .A2(_11497_ ), .ZN(_11498_ ) );
INV_X1 _18188_ ( .A(_11498_ ), .ZN(_11499_ ) );
BUF_X4 _18189_ ( .A(_11499_ ), .Z(_11500_ ) );
AND2_X1 _18190_ ( .A1(\icache.offset_buf [1] ), .A2(\icache.offset_buf [0] ), .ZN(_11501_ ) );
CLKBUF_X2 _18191_ ( .A(_11501_ ), .Z(_11502_ ) );
CLKBUF_X2 _18192_ ( .A(_11502_ ), .Z(_11503_ ) );
AND3_X1 _18193_ ( .A1(\arbiter.io_ifu_araddr [4] ), .A2(\icache.icache_reg_1_3 [31] ), .A3(_11503_ ), .ZN(_11504_ ) );
BUF_X2 _18194_ ( .A(_10838_ ), .Z(_11505_ ) );
INV_X1 _18195_ ( .A(_11501_ ), .ZN(_11506_ ) );
NOR3_X1 _18196_ ( .A1(_11505_ ), .A2(\icache.icache_reg_0_3 [31] ), .A3(_11506_ ), .ZN(_11507_ ) );
INV_X1 _18197_ ( .A(\icache.offset_buf [0] ), .ZN(_11508_ ) );
NOR2_X1 _18198_ ( .A1(_11508_ ), .A2(\icache.offset_buf [1] ), .ZN(_11509_ ) );
INV_X1 _18199_ ( .A(_11509_ ), .ZN(_11510_ ) );
NOR2_X1 _18200_ ( .A1(_09818_ ), .A2(_11510_ ), .ZN(_11511_ ) );
BUF_X4 _18201_ ( .A(_11511_ ), .Z(_11512_ ) );
BUF_X4 _18202_ ( .A(_11512_ ), .Z(_11513_ ) );
BUF_X4 _18203_ ( .A(_11513_ ), .Z(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_ANDNOT__B_Y ) );
INV_X1 _18204_ ( .A(\icache.icache_reg_0_1 [31] ), .ZN(_11514_ ) );
BUF_X2 _18205_ ( .A(_10834_ ), .Z(_11515_ ) );
INV_X1 _18206_ ( .A(\icache.offset_buf [1] ), .ZN(_11516_ ) );
NOR2_X1 _18207_ ( .A1(_11516_ ), .A2(\icache.offset_buf [0] ), .ZN(_11517_ ) );
BUF_X4 _18208_ ( .A(_11517_ ), .Z(_11518_ ) );
AOI22_X1 _18209_ ( .A1(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_ANDNOT__B_Y ), .A2(_11514_ ), .B1(_11515_ ), .B2(_11518_ ), .ZN(_11519_ ) );
OAI21_X1 _18210_ ( .A(_11519_ ), .B1(\icache.icache_reg_0_0 [31] ), .B2(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_ANDNOT__B_Y ), .ZN(_11520_ ) );
OAI211_X1 _18211_ ( .A(_10835_ ), .B(\icache.offset_buf [1] ), .C1(\icache.icache_reg_0_2 [31] ), .C2(\icache.offset_buf [0] ), .ZN(_11521_ ) );
AOI21_X1 _18212_ ( .A(_11507_ ), .B1(_11520_ ), .B2(_11521_ ), .ZN(_11522_ ) );
NOR2_X1 _18213_ ( .A1(\icache.offset_buf [1] ), .A2(\icache.offset_buf [0] ), .ZN(_11523_ ) );
AND2_X2 _18214_ ( .A1(_10837_ ), .A2(_11523_ ), .ZN(\icache.offset_buf_$_OR__A_Y_$_NOR__A_Y ) );
INV_X2 _18215_ ( .A(\icache.offset_buf_$_OR__A_Y_$_NOR__A_Y ), .ZN(_11524_ ) );
BUF_X4 _18216_ ( .A(_11524_ ), .Z(_11525_ ) );
MUX2_X1 _18217_ ( .A(\icache.icache_reg_1_0 [31] ), .B(_11522_ ), .S(_11525_ ), .Z(_11526_ ) );
AND2_X1 _18218_ ( .A1(_10837_ ), .A2(_11509_ ), .ZN(_11527_ ) );
INV_X1 _18219_ ( .A(_11527_ ), .ZN(_11528_ ) );
BUF_X4 _18220_ ( .A(_11528_ ), .Z(_11529_ ) );
BUF_X4 _18221_ ( .A(_11529_ ), .Z(_11530_ ) );
MUX2_X1 _18222_ ( .A(\icache.icache_reg_1_1 [31] ), .B(_11526_ ), .S(_11530_ ), .Z(_11531_ ) );
AND2_X1 _18223_ ( .A1(_10838_ ), .A2(_11517_ ), .ZN(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_NOR__A_Y ) );
INV_X1 _18224_ ( .A(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_NOR__A_Y ), .ZN(_11532_ ) );
BUF_X4 _18225_ ( .A(_11532_ ), .Z(_11533_ ) );
BUF_X4 _18226_ ( .A(_11533_ ), .Z(_11534_ ) );
BUF_X4 _18227_ ( .A(_11534_ ), .Z(_11535_ ) );
MUX2_X1 _18228_ ( .A(\icache.icache_reg_1_2 [31] ), .B(_11531_ ), .S(_11535_ ), .Z(_11536_ ) );
AND2_X1 _18229_ ( .A1(_10839_ ), .A2(_11501_ ), .ZN(_11537_ ) );
INV_X1 _18230_ ( .A(_11537_ ), .ZN(_11538_ ) );
BUF_X4 _18231_ ( .A(_11538_ ), .Z(_11539_ ) );
BUF_X4 _18232_ ( .A(_11539_ ), .Z(_11540_ ) );
AOI21_X1 _18233_ ( .A(_11504_ ), .B1(_11536_ ), .B2(_11540_ ), .ZN(_11541_ ) );
AOI211_X1 _18234_ ( .A(fanout_net_19 ), .B(_11494_ ), .C1(_11500_ ), .C2(_11541_ ), .ZN(_00133_ ) );
OR3_X1 _18235_ ( .A1(\idu.io_out_valid_REG ), .A2(\idu.io_in_valid ), .A3(\idu.state ), .ZN(_11542_ ) );
AND4_X1 _18236_ ( .A1(_10788_ ), .A2(_10822_ ), .A3(_10828_ ), .A4(_11542_ ), .ZN(_exu_io_in_bits_T ) );
NAND3_X1 _18237_ ( .A1(_10788_ ), .A2(_10822_ ), .A3(_11542_ ), .ZN(_11543_ ) );
NOR4_X1 _18238_ ( .A1(_11543_ ), .A2(fanout_net_19 ), .A3(\exu.state ), .A4(_10991_ ), .ZN(_00134_ ) );
AOI211_X1 _18239_ ( .A(\io_master_rdata [30] ), .B(_11301_ ), .C1(_11489_ ), .C2(_11493_ ), .ZN(_11544_ ) );
AND3_X1 _18240_ ( .A1(\arbiter.io_ifu_araddr [4] ), .A2(\icache.icache_reg_1_3 [30] ), .A3(_11503_ ), .ZN(_11545_ ) );
MUX2_X1 _18241_ ( .A(\icache.icache_reg_0_0 [30] ), .B(\icache.icache_reg_0_1 [30] ), .S(_11513_ ), .Z(_11546_ ) );
INV_X1 _18242_ ( .A(_11517_ ), .ZN(_11547_ ) );
NOR2_X1 _18243_ ( .A1(_09818_ ), .A2(_11547_ ), .ZN(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_ANDNOT__B_Y ) );
INV_X1 _18244_ ( .A(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_ANDNOT__B_Y ), .ZN(_11548_ ) );
BUF_X4 _18245_ ( .A(_11548_ ), .Z(_11549_ ) );
BUF_X4 _18246_ ( .A(_11549_ ), .Z(_11550_ ) );
MUX2_X1 _18247_ ( .A(\icache.icache_reg_0_2 [30] ), .B(_11546_ ), .S(_11550_ ), .Z(_11551_ ) );
NOR2_X1 _18248_ ( .A1(_09818_ ), .A2(_11506_ ), .ZN(\icache.offset_buf_$_NAND__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _18249_ ( .A(\icache.offset_buf_$_NAND__A_Y_$_ANDNOT__B_Y ), .ZN(_11552_ ) );
BUF_X4 _18250_ ( .A(_11552_ ), .Z(_11553_ ) );
BUF_X4 _18251_ ( .A(_11553_ ), .Z(_11554_ ) );
MUX2_X1 _18252_ ( .A(\icache.icache_reg_0_3 [30] ), .B(_11551_ ), .S(_11554_ ), .Z(_11555_ ) );
MUX2_X1 _18253_ ( .A(\icache.icache_reg_1_0 [30] ), .B(_11555_ ), .S(_11525_ ), .Z(_11556_ ) );
MUX2_X1 _18254_ ( .A(\icache.icache_reg_1_1 [30] ), .B(_11556_ ), .S(_11530_ ), .Z(_11557_ ) );
MUX2_X1 _18255_ ( .A(\icache.icache_reg_1_2 [30] ), .B(_11557_ ), .S(_11535_ ), .Z(_11558_ ) );
AOI21_X1 _18256_ ( .A(_11545_ ), .B1(_11558_ ), .B2(_11540_ ), .ZN(_11559_ ) );
AOI211_X1 _18257_ ( .A(fanout_net_19 ), .B(_11544_ ), .C1(_11500_ ), .C2(_11559_ ), .ZN(_00135_ ) );
BUF_X4 _18258_ ( .A(_11537_ ), .Z(_11560_ ) );
BUF_X2 _18259_ ( .A(_09335_ ), .Z(_11561_ ) );
BUF_X2 _18260_ ( .A(_09337_ ), .Z(_11562_ ) );
AOI211_X1 _18261_ ( .A(\icache.icache_reg_1_2 [21] ), .B(_11547_ ), .C1(_11561_ ), .C2(_11562_ ), .ZN(_11563_ ) );
AND4_X1 _18262_ ( .A1(\icache.icache_reg_0_3 [21] ), .A2(_09335_ ), .A3(_09337_ ), .A4(_11501_ ), .ZN(_11564_ ) );
MUX2_X1 _18263_ ( .A(\icache.icache_reg_0_0 [21] ), .B(\icache.icache_reg_0_1 [21] ), .S(_11513_ ), .Z(_11565_ ) );
MUX2_X1 _18264_ ( .A(\icache.icache_reg_0_2 [21] ), .B(_11565_ ), .S(_11550_ ), .Z(_11566_ ) );
BUF_X4 _18265_ ( .A(_11554_ ), .Z(_11567_ ) );
AOI211_X1 _18266_ ( .A(\icache.offset_buf_$_OR__A_Y_$_NOR__A_Y ), .B(_11564_ ), .C1(_11566_ ), .C2(_11567_ ), .ZN(_11568_ ) );
BUF_X2 _18267_ ( .A(_11527_ ), .Z(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_NOR__A_Y ) );
NOR4_X1 _18268_ ( .A1(_10836_ ), .A2(\icache.icache_reg_1_0 [21] ), .A3(\icache.offset_buf [1] ), .A4(\icache.offset_buf [0] ), .ZN(_11569_ ) );
OR3_X1 _18269_ ( .A1(_11568_ ), .A2(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_NOR__A_Y ), .A3(_11569_ ), .ZN(_11570_ ) );
BUF_X2 _18270_ ( .A(_10839_ ), .Z(_11571_ ) );
BUF_X2 _18271_ ( .A(_11571_ ), .Z(_11572_ ) );
AOI22_X1 _18272_ ( .A1(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_NOR__A_Y ), .A2(\icache.icache_reg_1_1 [21] ), .B1(_11572_ ), .B2(_11518_ ), .ZN(_11573_ ) );
AOI211_X1 _18273_ ( .A(_11560_ ), .B(_11563_ ), .C1(_11570_ ), .C2(_11573_ ), .ZN(_11574_ ) );
BUF_X4 _18274_ ( .A(_11560_ ), .Z(_11575_ ) );
BUF_X4 _18275_ ( .A(_11496_ ), .Z(_11576_ ) );
BUF_X4 _18276_ ( .A(_11576_ ), .Z(_11577_ ) );
BUF_X4 _18277_ ( .A(_11497_ ), .Z(_11578_ ) );
AOI221_X4 _18278_ ( .A(_11574_ ), .B1(\icache.icache_reg_1_3 [21] ), .B2(_11575_ ), .C1(_11577_ ), .C2(_11578_ ), .ZN(_11579_ ) );
BUF_X4 _18279_ ( .A(_11300_ ), .Z(_11580_ ) );
BUF_X4 _18280_ ( .A(_11488_ ), .Z(_11581_ ) );
BUF_X4 _18281_ ( .A(_11581_ ), .Z(_11582_ ) );
BUF_X4 _18282_ ( .A(_11492_ ), .Z(_11583_ ) );
BUF_X4 _18283_ ( .A(_11583_ ), .Z(_11584_ ) );
AOI211_X1 _18284_ ( .A(\io_master_rdata [21] ), .B(_11580_ ), .C1(_11582_ ), .C2(_11584_ ), .ZN(_11585_ ) );
NOR3_X1 _18285_ ( .A1(_11579_ ), .A2(fanout_net_19 ), .A3(_11585_ ), .ZN(_00136_ ) );
AND3_X1 _18286_ ( .A1(_10841_ ), .A2(\icache.icache_reg_1_3 [20] ), .A3(_11502_ ), .ZN(_11586_ ) );
MUX2_X1 _18287_ ( .A(\icache.icache_reg_0_0 [20] ), .B(\icache.icache_reg_0_1 [20] ), .S(_11511_ ), .Z(_11587_ ) );
MUX2_X1 _18288_ ( .A(\icache.icache_reg_0_2 [20] ), .B(_11587_ ), .S(_11548_ ), .Z(_11588_ ) );
MUX2_X1 _18289_ ( .A(\icache.icache_reg_0_3 [20] ), .B(_11588_ ), .S(_11553_ ), .Z(_11589_ ) );
MUX2_X1 _18290_ ( .A(\icache.icache_reg_1_0 [20] ), .B(_11589_ ), .S(_11524_ ), .Z(_11590_ ) );
MUX2_X1 _18291_ ( .A(\icache.icache_reg_1_1 [20] ), .B(_11590_ ), .S(_11528_ ), .Z(_11591_ ) );
MUX2_X1 _18292_ ( .A(\icache.icache_reg_1_2 [20] ), .B(_11591_ ), .S(_11533_ ), .Z(_11592_ ) );
AOI221_X4 _18293_ ( .A(_11586_ ), .B1(_11539_ ), .B2(_11592_ ), .C1(_11577_ ), .C2(_11578_ ), .ZN(_11593_ ) );
AOI211_X1 _18294_ ( .A(\io_master_rdata [20] ), .B(_11580_ ), .C1(_11582_ ), .C2(_11584_ ), .ZN(_11594_ ) );
NOR3_X1 _18295_ ( .A1(_11593_ ), .A2(fanout_net_19 ), .A3(_11594_ ), .ZN(_00137_ ) );
AND3_X1 _18296_ ( .A1(_10841_ ), .A2(\icache.icache_reg_1_3 [19] ), .A3(_11502_ ), .ZN(_11595_ ) );
NOR3_X1 _18297_ ( .A1(_10838_ ), .A2(\icache.icache_reg_0_3 [19] ), .A3(_11506_ ), .ZN(_11596_ ) );
NOR3_X1 _18298_ ( .A1(_10837_ ), .A2(\icache.icache_reg_0_1 [19] ), .A3(_11510_ ), .ZN(_11597_ ) );
NOR2_X1 _18299_ ( .A1(_11597_ ), .A2(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_ANDNOT__B_Y ), .ZN(_11598_ ) );
OAI21_X1 _18300_ ( .A(_11598_ ), .B1(\icache.icache_reg_0_0 [19] ), .B2(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_ANDNOT__B_Y ), .ZN(_11599_ ) );
OAI211_X1 _18301_ ( .A(_10834_ ), .B(\icache.offset_buf [1] ), .C1(\icache.icache_reg_0_2 [19] ), .C2(\icache.offset_buf [0] ), .ZN(_11600_ ) );
AOI21_X1 _18302_ ( .A(_11596_ ), .B1(_11599_ ), .B2(_11600_ ), .ZN(_11601_ ) );
MUX2_X1 _18303_ ( .A(\icache.icache_reg_1_0 [19] ), .B(_11601_ ), .S(_11524_ ), .Z(_11602_ ) );
MUX2_X1 _18304_ ( .A(\icache.icache_reg_1_1 [19] ), .B(_11602_ ), .S(_11528_ ), .Z(_11603_ ) );
MUX2_X1 _18305_ ( .A(\icache.icache_reg_1_2 [19] ), .B(_11603_ ), .S(_11533_ ), .Z(_11604_ ) );
AOI221_X4 _18306_ ( .A(_11595_ ), .B1(_11539_ ), .B2(_11604_ ), .C1(_11577_ ), .C2(_11578_ ), .ZN(_11605_ ) );
AOI211_X1 _18307_ ( .A(\io_master_rdata [19] ), .B(_11580_ ), .C1(_11582_ ), .C2(_11584_ ), .ZN(_11606_ ) );
NOR3_X1 _18308_ ( .A1(_11605_ ), .A2(fanout_net_19 ), .A3(_11606_ ), .ZN(_00138_ ) );
INV_X1 _18309_ ( .A(\icache.icache_reg_1_3 [18] ), .ZN(_11607_ ) );
NAND3_X1 _18310_ ( .A1(\arbiter.io_ifu_araddr [4] ), .A2(_11607_ ), .A3(_11503_ ), .ZN(_11608_ ) );
MUX2_X1 _18311_ ( .A(\icache.icache_reg_0_0 [18] ), .B(\icache.icache_reg_0_1 [18] ), .S(_11512_ ), .Z(_11609_ ) );
MUX2_X1 _18312_ ( .A(\icache.icache_reg_0_2 [18] ), .B(_11609_ ), .S(_11549_ ), .Z(_11610_ ) );
MUX2_X1 _18313_ ( .A(\icache.icache_reg_0_3 [18] ), .B(_11610_ ), .S(_11553_ ), .Z(_11611_ ) );
BUF_X4 _18314_ ( .A(_11524_ ), .Z(_11612_ ) );
MUX2_X1 _18315_ ( .A(\icache.icache_reg_1_0 [18] ), .B(_11611_ ), .S(_11612_ ), .Z(_11613_ ) );
MUX2_X1 _18316_ ( .A(\icache.icache_reg_1_1 [18] ), .B(_11613_ ), .S(_11529_ ), .Z(_11614_ ) );
MUX2_X1 _18317_ ( .A(\icache.icache_reg_1_2 [18] ), .B(_11614_ ), .S(_11534_ ), .Z(_11615_ ) );
OAI221_X1 _18318_ ( .A(_11608_ ), .B1(_11575_ ), .B2(_11615_ ), .C1(_11495_ ), .C2(_11580_ ), .ZN(_11616_ ) );
NAND3_X1 _18319_ ( .A1(_11577_ ), .A2(\io_master_rdata [18] ), .A3(_11578_ ), .ZN(_11617_ ) );
AOI21_X1 _18320_ ( .A(fanout_net_19 ), .B1(_11616_ ), .B2(_11617_ ), .ZN(_00139_ ) );
MUX2_X1 _18321_ ( .A(\icache.icache_reg_0_0 [17] ), .B(\icache.icache_reg_0_1 [17] ), .S(_11512_ ), .Z(_11618_ ) );
MUX2_X1 _18322_ ( .A(\icache.icache_reg_0_2 [17] ), .B(_11618_ ), .S(_11548_ ), .Z(_11619_ ) );
MUX2_X1 _18323_ ( .A(\icache.icache_reg_0_3 [17] ), .B(_11619_ ), .S(_11553_ ), .Z(_11620_ ) );
MUX2_X1 _18324_ ( .A(\icache.icache_reg_1_0 [17] ), .B(_11620_ ), .S(_11524_ ), .Z(_11621_ ) );
MUX2_X1 _18325_ ( .A(\icache.icache_reg_1_1 [17] ), .B(_11621_ ), .S(_11529_ ), .Z(_11622_ ) );
NAND2_X1 _18326_ ( .A1(_11622_ ), .A2(_11533_ ), .ZN(_11623_ ) );
NAND3_X1 _18327_ ( .A1(_11572_ ), .A2(\icache.icache_reg_1_2 [17] ), .A3(_11518_ ), .ZN(_11624_ ) );
AOI21_X1 _18328_ ( .A(_11560_ ), .B1(_11623_ ), .B2(_11624_ ), .ZN(_11625_ ) );
AOI221_X4 _18329_ ( .A(_11625_ ), .B1(\icache.icache_reg_1_3 [17] ), .B2(_11560_ ), .C1(_11576_ ), .C2(_11497_ ), .ZN(_11626_ ) );
INV_X1 _18330_ ( .A(\io_master_rdata [17] ), .ZN(_11627_ ) );
AOI211_X1 _18331_ ( .A(fanout_net_19 ), .B(_11626_ ), .C1(_11627_ ), .C2(_11498_ ), .ZN(_00140_ ) );
AND3_X1 _18332_ ( .A1(_11572_ ), .A2(\icache.icache_reg_1_3 [16] ), .A3(_11502_ ), .ZN(_11628_ ) );
MUX2_X1 _18333_ ( .A(\icache.icache_reg_0_0 [16] ), .B(\icache.icache_reg_0_1 [16] ), .S(_11511_ ), .Z(_11629_ ) );
MUX2_X1 _18334_ ( .A(\icache.icache_reg_0_2 [16] ), .B(_11629_ ), .S(_11548_ ), .Z(_11630_ ) );
MUX2_X1 _18335_ ( .A(\icache.icache_reg_0_3 [16] ), .B(_11630_ ), .S(_11552_ ), .Z(_11631_ ) );
MUX2_X1 _18336_ ( .A(\icache.icache_reg_1_0 [16] ), .B(_11631_ ), .S(_11524_ ), .Z(_11632_ ) );
MUX2_X1 _18337_ ( .A(\icache.icache_reg_1_1 [16] ), .B(_11632_ ), .S(_11528_ ), .Z(_11633_ ) );
MUX2_X1 _18338_ ( .A(\icache.icache_reg_1_2 [16] ), .B(_11633_ ), .S(_11533_ ), .Z(_11634_ ) );
AOI221_X4 _18339_ ( .A(_11628_ ), .B1(_11539_ ), .B2(_11634_ ), .C1(_11576_ ), .C2(_11497_ ), .ZN(_11635_ ) );
INV_X1 _18340_ ( .A(\io_master_rdata [16] ), .ZN(_11636_ ) );
AOI211_X1 _18341_ ( .A(fanout_net_19 ), .B(_11635_ ), .C1(_11636_ ), .C2(_11498_ ), .ZN(_00141_ ) );
MUX2_X1 _18342_ ( .A(\icache.icache_reg_0_0 [15] ), .B(\icache.icache_reg_0_1 [15] ), .S(_11512_ ), .Z(_11637_ ) );
MUX2_X1 _18343_ ( .A(\icache.icache_reg_0_2 [15] ), .B(_11637_ ), .S(_11549_ ), .Z(_11638_ ) );
MUX2_X1 _18344_ ( .A(\icache.icache_reg_0_3 [15] ), .B(_11638_ ), .S(_11553_ ), .Z(_11639_ ) );
MUX2_X1 _18345_ ( .A(\icache.icache_reg_1_0 [15] ), .B(_11639_ ), .S(_11524_ ), .Z(_11640_ ) );
MUX2_X1 _18346_ ( .A(\icache.icache_reg_1_1 [15] ), .B(_11640_ ), .S(_11529_ ), .Z(_11641_ ) );
NAND2_X1 _18347_ ( .A1(_11641_ ), .A2(_11534_ ), .ZN(_11642_ ) );
BUF_X2 _18348_ ( .A(_10840_ ), .Z(_11643_ ) );
NAND3_X1 _18349_ ( .A1(_11643_ ), .A2(\icache.icache_reg_1_2 [15] ), .A3(_11518_ ), .ZN(_11644_ ) );
AOI21_X1 _18350_ ( .A(_11560_ ), .B1(_11642_ ), .B2(_11644_ ), .ZN(_11645_ ) );
AOI221_X4 _18351_ ( .A(_11645_ ), .B1(\icache.icache_reg_1_3 [15] ), .B2(_11575_ ), .C1(_11577_ ), .C2(_11578_ ), .ZN(_11646_ ) );
AOI211_X1 _18352_ ( .A(\io_master_rdata [15] ), .B(_11580_ ), .C1(_11582_ ), .C2(_11584_ ), .ZN(_11647_ ) );
NOR3_X1 _18353_ ( .A1(_11646_ ), .A2(fanout_net_20 ), .A3(_11647_ ), .ZN(_00142_ ) );
BUF_X4 _18354_ ( .A(_11300_ ), .Z(_11648_ ) );
AOI211_X1 _18355_ ( .A(\io_master_rdata [14] ), .B(_11648_ ), .C1(_11489_ ), .C2(_11493_ ), .ZN(_11649_ ) );
AND3_X1 _18356_ ( .A1(\arbiter.io_ifu_araddr [4] ), .A2(\icache.icache_reg_1_3 [14] ), .A3(_11503_ ), .ZN(_11650_ ) );
MUX2_X1 _18357_ ( .A(\icache.icache_reg_0_0 [14] ), .B(\icache.icache_reg_0_1 [14] ), .S(_11513_ ), .Z(_11651_ ) );
MUX2_X1 _18358_ ( .A(\icache.icache_reg_0_2 [14] ), .B(_11651_ ), .S(_11550_ ), .Z(_11652_ ) );
MUX2_X1 _18359_ ( .A(\icache.icache_reg_0_3 [14] ), .B(_11652_ ), .S(_11554_ ), .Z(_11653_ ) );
MUX2_X1 _18360_ ( .A(\icache.icache_reg_1_0 [14] ), .B(_11653_ ), .S(_11525_ ), .Z(_11654_ ) );
MUX2_X1 _18361_ ( .A(\icache.icache_reg_1_1 [14] ), .B(_11654_ ), .S(_11530_ ), .Z(_11655_ ) );
MUX2_X1 _18362_ ( .A(\icache.icache_reg_1_2 [14] ), .B(_11655_ ), .S(_11535_ ), .Z(_11656_ ) );
AOI21_X1 _18363_ ( .A(_11650_ ), .B1(_11656_ ), .B2(_11540_ ), .ZN(_11657_ ) );
AOI211_X1 _18364_ ( .A(fanout_net_20 ), .B(_11649_ ), .C1(_11500_ ), .C2(_11657_ ), .ZN(_00143_ ) );
AOI211_X1 _18365_ ( .A(\icache.icache_reg_1_2 [13] ), .B(_11547_ ), .C1(_11561_ ), .C2(_11562_ ), .ZN(_11658_ ) );
OR3_X1 _18366_ ( .A1(_11505_ ), .A2(\icache.icache_reg_0_2 [13] ), .A3(_11547_ ), .ZN(_11659_ ) );
MUX2_X1 _18367_ ( .A(\icache.icache_reg_0_0 [13] ), .B(\icache.icache_reg_0_1 [13] ), .S(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_ANDNOT__B_Y ), .Z(_11660_ ) );
OAI211_X1 _18368_ ( .A(_11567_ ), .B(_11659_ ), .C1(_11660_ ), .C2(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_ANDNOT__B_Y ), .ZN(_11661_ ) );
NAND4_X1 _18369_ ( .A1(_11561_ ), .A2(\icache.icache_reg_0_3 [13] ), .A3(_11562_ ), .A4(_11501_ ), .ZN(_11662_ ) );
AOI21_X1 _18370_ ( .A(\icache.offset_buf_$_OR__A_Y_$_NOR__A_Y ), .B1(_11661_ ), .B2(_11662_ ), .ZN(_11663_ ) );
AND3_X1 _18371_ ( .A1(_10840_ ), .A2(\icache.icache_reg_1_0 [13] ), .A3(_11523_ ), .ZN(_11664_ ) );
OAI21_X1 _18372_ ( .A(_11530_ ), .B1(_11663_ ), .B2(_11664_ ), .ZN(_11665_ ) );
AOI22_X1 _18373_ ( .A1(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_NOR__A_Y ), .A2(\icache.icache_reg_1_1 [13] ), .B1(_11572_ ), .B2(_11518_ ), .ZN(_11666_ ) );
AOI211_X1 _18374_ ( .A(_11560_ ), .B(_11658_ ), .C1(_11665_ ), .C2(_11666_ ), .ZN(_11667_ ) );
AOI221_X4 _18375_ ( .A(_11667_ ), .B1(\icache.icache_reg_1_3 [13] ), .B2(_11575_ ), .C1(_11577_ ), .C2(_11578_ ), .ZN(_11668_ ) );
AOI211_X1 _18376_ ( .A(\io_master_rdata [13] ), .B(_11301_ ), .C1(_11582_ ), .C2(_11584_ ), .ZN(_11669_ ) );
NOR3_X1 _18377_ ( .A1(_11668_ ), .A2(fanout_net_20 ), .A3(_11669_ ), .ZN(_00144_ ) );
AOI211_X1 _18378_ ( .A(\io_master_rdata [12] ), .B(_11648_ ), .C1(_11489_ ), .C2(_11493_ ), .ZN(_11670_ ) );
AND3_X1 _18379_ ( .A1(\arbiter.io_ifu_araddr [4] ), .A2(\icache.icache_reg_1_3 [12] ), .A3(_11503_ ), .ZN(_11671_ ) );
NOR4_X1 _18380_ ( .A1(_10836_ ), .A2(\icache.icache_reg_1_0 [12] ), .A3(\icache.offset_buf [1] ), .A4(\icache.offset_buf [0] ), .ZN(_11672_ ) );
INV_X1 _18381_ ( .A(\icache.icache_reg_0_3 [12] ), .ZN(_11673_ ) );
OR3_X1 _18382_ ( .A1(_11505_ ), .A2(\icache.icache_reg_0_2 [12] ), .A3(_11547_ ), .ZN(_11674_ ) );
MUX2_X1 _18383_ ( .A(\icache.icache_reg_0_0 [12] ), .B(\icache.icache_reg_0_1 [12] ), .S(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_ANDNOT__B_Y ), .Z(_11675_ ) );
OAI21_X1 _18384_ ( .A(_11674_ ), .B1(_11675_ ), .B2(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_ANDNOT__B_Y ), .ZN(_11676_ ) );
MUX2_X1 _18385_ ( .A(_11673_ ), .B(_11676_ ), .S(_11567_ ), .Z(_11677_ ) );
AOI211_X1 _18386_ ( .A(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_NOR__A_Y ), .B(_11672_ ), .C1(_11677_ ), .C2(_11525_ ), .ZN(_11678_ ) );
AOI211_X1 _18387_ ( .A(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_NOR__A_Y ), .B(_11678_ ), .C1(\icache.icache_reg_1_1 [12] ), .C2(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_NOR__A_Y ), .ZN(_11679_ ) );
AOI211_X1 _18388_ ( .A(\icache.icache_reg_1_2 [12] ), .B(_11547_ ), .C1(_11561_ ), .C2(_11562_ ), .ZN(_11680_ ) );
NOR2_X1 _18389_ ( .A1(_11679_ ), .A2(_11680_ ), .ZN(_11681_ ) );
AOI21_X1 _18390_ ( .A(_11671_ ), .B1(_11681_ ), .B2(_11540_ ), .ZN(_11682_ ) );
AOI211_X1 _18391_ ( .A(fanout_net_20 ), .B(_11670_ ), .C1(_11500_ ), .C2(_11682_ ), .ZN(_00145_ ) );
AND3_X1 _18392_ ( .A1(_10841_ ), .A2(\icache.icache_reg_1_3 [29] ), .A3(_11502_ ), .ZN(_11683_ ) );
MUX2_X1 _18393_ ( .A(\icache.icache_reg_0_0 [29] ), .B(\icache.icache_reg_0_1 [29] ), .S(_11511_ ), .Z(_11684_ ) );
MUX2_X1 _18394_ ( .A(\icache.icache_reg_0_2 [29] ), .B(_11684_ ), .S(_11548_ ), .Z(_11685_ ) );
MUX2_X1 _18395_ ( .A(\icache.icache_reg_0_3 [29] ), .B(_11685_ ), .S(_11552_ ), .Z(_11686_ ) );
MUX2_X1 _18396_ ( .A(\icache.icache_reg_1_0 [29] ), .B(_11686_ ), .S(_11524_ ), .Z(_11687_ ) );
MUX2_X1 _18397_ ( .A(\icache.icache_reg_1_1 [29] ), .B(_11687_ ), .S(_11528_ ), .Z(_11688_ ) );
MUX2_X1 _18398_ ( .A(\icache.icache_reg_1_2 [29] ), .B(_11688_ ), .S(_11533_ ), .Z(_11689_ ) );
AOI221_X4 _18399_ ( .A(_11683_ ), .B1(_11539_ ), .B2(_11689_ ), .C1(_11576_ ), .C2(_11578_ ), .ZN(_11690_ ) );
AOI211_X1 _18400_ ( .A(\io_master_rdata [29] ), .B(_11301_ ), .C1(_11582_ ), .C2(_11584_ ), .ZN(_11691_ ) );
NOR3_X1 _18401_ ( .A1(_11690_ ), .A2(fanout_net_20 ), .A3(_11691_ ), .ZN(_00146_ ) );
AOI211_X1 _18402_ ( .A(\io_master_rdata [11] ), .B(_11648_ ), .C1(_11489_ ), .C2(_11493_ ), .ZN(_11692_ ) );
OR3_X1 _18403_ ( .A1(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__A_Y ), .A2(\icache.icache_reg_1_3 [11] ), .A3(_11506_ ), .ZN(_11693_ ) );
MUX2_X1 _18404_ ( .A(\icache.icache_reg_0_0 [11] ), .B(\icache.icache_reg_0_1 [11] ), .S(_11513_ ), .Z(_11694_ ) );
MUX2_X1 _18405_ ( .A(\icache.icache_reg_0_2 [11] ), .B(_11694_ ), .S(_11550_ ), .Z(_11695_ ) );
MUX2_X1 _18406_ ( .A(\icache.icache_reg_0_3 [11] ), .B(_11695_ ), .S(_11554_ ), .Z(_11696_ ) );
MUX2_X1 _18407_ ( .A(\icache.icache_reg_1_0 [11] ), .B(_11696_ ), .S(_11612_ ), .Z(_11697_ ) );
MUX2_X1 _18408_ ( .A(\icache.icache_reg_1_1 [11] ), .B(_11697_ ), .S(_11530_ ), .Z(_11698_ ) );
MUX2_X1 _18409_ ( .A(\icache.icache_reg_1_2 [11] ), .B(_11698_ ), .S(_11535_ ), .Z(_11699_ ) );
OAI21_X1 _18410_ ( .A(_11693_ ), .B1(_11699_ ), .B2(_11575_ ), .ZN(_11700_ ) );
AOI211_X1 _18411_ ( .A(fanout_net_20 ), .B(_11692_ ), .C1(_11500_ ), .C2(_11700_ ), .ZN(_00147_ ) );
AND3_X1 _18412_ ( .A1(_11643_ ), .A2(\icache.icache_reg_1_3 [10] ), .A3(_11502_ ), .ZN(_11701_ ) );
MUX2_X1 _18413_ ( .A(\icache.icache_reg_0_0 [10] ), .B(\icache.icache_reg_0_1 [10] ), .S(_11511_ ), .Z(_11702_ ) );
MUX2_X1 _18414_ ( .A(\icache.icache_reg_0_2 [10] ), .B(_11702_ ), .S(_11548_ ), .Z(_11703_ ) );
MUX2_X1 _18415_ ( .A(\icache.icache_reg_0_3 [10] ), .B(_11703_ ), .S(_11552_ ), .Z(_11704_ ) );
MUX2_X1 _18416_ ( .A(\icache.icache_reg_1_0 [10] ), .B(_11704_ ), .S(_11524_ ), .Z(_11705_ ) );
MUX2_X1 _18417_ ( .A(\icache.icache_reg_1_1 [10] ), .B(_11705_ ), .S(_11528_ ), .Z(_11706_ ) );
MUX2_X1 _18418_ ( .A(\icache.icache_reg_1_2 [10] ), .B(_11706_ ), .S(_11533_ ), .Z(_11707_ ) );
AOI221_X4 _18419_ ( .A(_11701_ ), .B1(_11539_ ), .B2(_11707_ ), .C1(_11576_ ), .C2(_11497_ ), .ZN(_11708_ ) );
AOI211_X1 _18420_ ( .A(\io_master_rdata [10] ), .B(_11301_ ), .C1(_11582_ ), .C2(_11584_ ), .ZN(_11709_ ) );
NOR3_X1 _18421_ ( .A1(_11708_ ), .A2(fanout_net_20 ), .A3(_11709_ ), .ZN(_00148_ ) );
OR3_X1 _18422_ ( .A1(_11495_ ), .A2(\io_master_rdata [9] ), .A3(_11300_ ), .ZN(_11710_ ) );
NAND3_X1 _18423_ ( .A1(\arbiter.io_ifu_araddr [4] ), .A2(\icache.icache_reg_1_3 [9] ), .A3(_11503_ ), .ZN(_11711_ ) );
NAND3_X1 _18424_ ( .A1(_10836_ ), .A2(\icache.icache_reg_0_2 [9] ), .A3(_11518_ ), .ZN(_11712_ ) );
AND4_X1 _18425_ ( .A1(\icache.icache_reg_0_1 [9] ), .A2(_09335_ ), .A3(_09337_ ), .A4(_11509_ ), .ZN(_11713_ ) );
INV_X1 _18426_ ( .A(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_ANDNOT__B_Y ), .ZN(_11714_ ) );
AOI21_X1 _18427_ ( .A(_11713_ ), .B1(_11714_ ), .B2(\icache.icache_reg_0_0 [9] ), .ZN(_11715_ ) );
OAI211_X1 _18428_ ( .A(_11567_ ), .B(_11712_ ), .C1(_11715_ ), .C2(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_ANDNOT__B_Y ), .ZN(_11716_ ) );
OAI211_X1 _18429_ ( .A(_11716_ ), .B(_11525_ ), .C1(\icache.icache_reg_0_3 [9] ), .C2(_11567_ ), .ZN(_11717_ ) );
NAND3_X1 _18430_ ( .A1(_11643_ ), .A2(\icache.icache_reg_1_0 [9] ), .A3(_11523_ ), .ZN(_11718_ ) );
AOI21_X1 _18431_ ( .A(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_NOR__A_Y ), .B1(_11717_ ), .B2(_11718_ ), .ZN(_11719_ ) );
NAND3_X1 _18432_ ( .A1(_11643_ ), .A2(\icache.icache_reg_1_1 [9] ), .A3(_11509_ ), .ZN(_11720_ ) );
OAI21_X1 _18433_ ( .A(_11720_ ), .B1(_10836_ ), .B2(_11547_ ), .ZN(_11721_ ) );
OAI221_X1 _18434_ ( .A(_11539_ ), .B1(\icache.icache_reg_1_2 [9] ), .B2(_11534_ ), .C1(_11719_ ), .C2(_11721_ ), .ZN(_11722_ ) );
OAI211_X1 _18435_ ( .A(_11711_ ), .B(_11722_ ), .C1(_11495_ ), .C2(_11580_ ), .ZN(_11723_ ) );
AND3_X1 _18436_ ( .A1(_11710_ ), .A2(_10992_ ), .A3(_11723_ ), .ZN(_00149_ ) );
AOI211_X1 _18437_ ( .A(\io_master_rdata [8] ), .B(_11648_ ), .C1(_11581_ ), .C2(_11583_ ), .ZN(_11724_ ) );
OR3_X1 _18438_ ( .A1(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__A_Y ), .A2(\icache.icache_reg_1_3 [8] ), .A3(_11506_ ), .ZN(_11725_ ) );
MUX2_X1 _18439_ ( .A(\icache.icache_reg_0_0 [8] ), .B(\icache.icache_reg_0_1 [8] ), .S(_11513_ ), .Z(_11726_ ) );
MUX2_X1 _18440_ ( .A(\icache.icache_reg_0_2 [8] ), .B(_11726_ ), .S(_11549_ ), .Z(_11727_ ) );
MUX2_X1 _18441_ ( .A(\icache.icache_reg_0_3 [8] ), .B(_11727_ ), .S(_11554_ ), .Z(_11728_ ) );
MUX2_X1 _18442_ ( .A(\icache.icache_reg_1_0 [8] ), .B(_11728_ ), .S(_11612_ ), .Z(_11729_ ) );
MUX2_X1 _18443_ ( .A(\icache.icache_reg_1_1 [8] ), .B(_11729_ ), .S(_11529_ ), .Z(_11730_ ) );
MUX2_X1 _18444_ ( .A(\icache.icache_reg_1_2 [8] ), .B(_11730_ ), .S(_11534_ ), .Z(_11731_ ) );
OAI21_X1 _18445_ ( .A(_11725_ ), .B1(_11731_ ), .B2(_11575_ ), .ZN(_11732_ ) );
AOI211_X1 _18446_ ( .A(fanout_net_20 ), .B(_11724_ ), .C1(_11500_ ), .C2(_11732_ ), .ZN(_00150_ ) );
AOI211_X1 _18447_ ( .A(\io_master_rdata [7] ), .B(_11648_ ), .C1(_11581_ ), .C2(_11583_ ), .ZN(_11733_ ) );
AND3_X1 _18448_ ( .A1(\arbiter.io_ifu_araddr [4] ), .A2(\icache.icache_reg_1_3 [7] ), .A3(_11503_ ), .ZN(_11734_ ) );
MUX2_X1 _18449_ ( .A(\icache.icache_reg_0_0 [7] ), .B(\icache.icache_reg_0_1 [7] ), .S(_11513_ ), .Z(_11735_ ) );
MUX2_X1 _18450_ ( .A(\icache.icache_reg_0_2 [7] ), .B(_11735_ ), .S(_11550_ ), .Z(_11736_ ) );
MUX2_X1 _18451_ ( .A(\icache.icache_reg_0_3 [7] ), .B(_11736_ ), .S(_11554_ ), .Z(_11737_ ) );
MUX2_X1 _18452_ ( .A(\icache.icache_reg_1_0 [7] ), .B(_11737_ ), .S(_11525_ ), .Z(_11738_ ) );
MUX2_X1 _18453_ ( .A(\icache.icache_reg_1_1 [7] ), .B(_11738_ ), .S(_11530_ ), .Z(_11739_ ) );
MUX2_X1 _18454_ ( .A(\icache.icache_reg_1_2 [7] ), .B(_11739_ ), .S(_11535_ ), .Z(_11740_ ) );
AOI21_X1 _18455_ ( .A(_11734_ ), .B1(_11740_ ), .B2(_11540_ ), .ZN(_11741_ ) );
AOI211_X1 _18456_ ( .A(fanout_net_20 ), .B(_11733_ ), .C1(_11500_ ), .C2(_11741_ ), .ZN(_00151_ ) );
MUX2_X1 _18457_ ( .A(\icache.icache_reg_0_0 [6] ), .B(\icache.icache_reg_0_1 [6] ), .S(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_ANDNOT__B_Y ), .Z(_11742_ ) );
AND2_X1 _18458_ ( .A1(_11742_ ), .A2(_11550_ ), .ZN(_11743_ ) );
INV_X1 _18459_ ( .A(\icache.icache_reg_0_2 [6] ), .ZN(_11744_ ) );
AOI211_X1 _18460_ ( .A(_11516_ ), .B(_10840_ ), .C1(_11744_ ), .C2(_11508_ ), .ZN(_11745_ ) );
OAI221_X1 _18461_ ( .A(_11525_ ), .B1(\icache.icache_reg_0_3 [6] ), .B2(_11567_ ), .C1(_11743_ ), .C2(_11745_ ), .ZN(_11746_ ) );
NAND3_X1 _18462_ ( .A1(_10841_ ), .A2(\icache.icache_reg_1_0 [6] ), .A3(_11523_ ), .ZN(_11747_ ) );
AOI21_X1 _18463_ ( .A(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_NOR__A_Y ), .B1(_11746_ ), .B2(_11747_ ), .ZN(_11748_ ) );
NAND3_X1 _18464_ ( .A1(_10841_ ), .A2(\icache.icache_reg_1_1 [6] ), .A3(_11509_ ), .ZN(_11749_ ) );
OAI21_X1 _18465_ ( .A(_11749_ ), .B1(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__A_Y ), .B2(_11547_ ), .ZN(_11750_ ) );
OAI221_X1 _18466_ ( .A(_11539_ ), .B1(\icache.icache_reg_1_2 [6] ), .B2(_11535_ ), .C1(_11748_ ), .C2(_11750_ ), .ZN(_11751_ ) );
NAND3_X1 _18467_ ( .A1(\arbiter.io_ifu_araddr [4] ), .A2(\icache.icache_reg_1_3 [6] ), .A3(_11503_ ), .ZN(_11752_ ) );
AND3_X1 _18468_ ( .A1(_11499_ ), .A2(_11751_ ), .A3(_11752_ ), .ZN(_11753_ ) );
AOI211_X1 _18469_ ( .A(\io_master_rdata [6] ), .B(_11301_ ), .C1(_11489_ ), .C2(_11493_ ), .ZN(_11754_ ) );
NOR3_X1 _18470_ ( .A1(_11753_ ), .A2(fanout_net_20 ), .A3(_11754_ ), .ZN(_00152_ ) );
AND3_X1 _18471_ ( .A1(_11643_ ), .A2(\icache.icache_reg_1_3 [5] ), .A3(_11502_ ), .ZN(_11755_ ) );
AND3_X1 _18472_ ( .A1(_11505_ ), .A2(\icache.icache_reg_1_0 [5] ), .A3(_11523_ ), .ZN(_11756_ ) );
MUX2_X1 _18473_ ( .A(\icache.icache_reg_0_0 [5] ), .B(\icache.icache_reg_0_1 [5] ), .S(_11512_ ), .Z(_11757_ ) );
MUX2_X1 _18474_ ( .A(\icache.icache_reg_0_2 [5] ), .B(_11757_ ), .S(_11549_ ), .Z(_11758_ ) );
MUX2_X1 _18475_ ( .A(\icache.icache_reg_0_3 [5] ), .B(_11758_ ), .S(_11553_ ), .Z(_11759_ ) );
AOI211_X1 _18476_ ( .A(_11527_ ), .B(_11756_ ), .C1(_11759_ ), .C2(_11612_ ), .ZN(_11760_ ) );
AOI211_X1 _18477_ ( .A(\icache.icache_reg_1_1 [5] ), .B(_11510_ ), .C1(_11561_ ), .C2(_11562_ ), .ZN(_11761_ ) );
NOR2_X1 _18478_ ( .A1(_11760_ ), .A2(_11761_ ), .ZN(_11762_ ) );
MUX2_X1 _18479_ ( .A(\icache.icache_reg_1_2 [5] ), .B(_11762_ ), .S(_11533_ ), .Z(_11763_ ) );
AOI221_X4 _18480_ ( .A(_11755_ ), .B1(_11539_ ), .B2(_11763_ ), .C1(_11576_ ), .C2(_11497_ ), .ZN(_11764_ ) );
AOI211_X1 _18481_ ( .A(\io_master_rdata [5] ), .B(_11301_ ), .C1(_11489_ ), .C2(_11493_ ), .ZN(_11765_ ) );
NOR3_X1 _18482_ ( .A1(_11764_ ), .A2(fanout_net_20 ), .A3(_11765_ ), .ZN(_00153_ ) );
NAND3_X1 _18483_ ( .A1(_10835_ ), .A2(\icache.icache_reg_0_2 [4] ), .A3(_11518_ ), .ZN(_11766_ ) );
OAI22_X1 _18484_ ( .A1(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_ANDNOT__B_Y ), .A2(\icache.icache_reg_0_0 [4] ), .B1(_11505_ ), .B2(_11547_ ), .ZN(_11767_ ) );
NOR3_X1 _18485_ ( .A1(_11505_ ), .A2(\icache.icache_reg_0_1 [4] ), .A3(_11510_ ), .ZN(_11768_ ) );
OAI211_X1 _18486_ ( .A(_11567_ ), .B(_11766_ ), .C1(_11767_ ), .C2(_11768_ ), .ZN(_11769_ ) );
OAI211_X1 _18487_ ( .A(_11769_ ), .B(_11525_ ), .C1(\icache.icache_reg_0_3 [4] ), .C2(_11567_ ), .ZN(_11770_ ) );
NAND3_X1 _18488_ ( .A1(_10840_ ), .A2(\icache.icache_reg_1_0 [4] ), .A3(_11523_ ), .ZN(_11771_ ) );
AOI21_X1 _18489_ ( .A(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_NOR__A_Y ), .B1(_11770_ ), .B2(_11771_ ), .ZN(_11772_ ) );
INV_X1 _18490_ ( .A(\icache.icache_reg_1_1 [4] ), .ZN(_11773_ ) );
AOI211_X1 _18491_ ( .A(_11773_ ), .B(_11510_ ), .C1(_11561_ ), .C2(_11562_ ), .ZN(_11774_ ) );
OAI21_X1 _18492_ ( .A(_11533_ ), .B1(_11772_ ), .B2(_11774_ ), .ZN(_11775_ ) );
NAND3_X1 _18493_ ( .A1(_11643_ ), .A2(\icache.icache_reg_1_2 [4] ), .A3(_11518_ ), .ZN(_11776_ ) );
AOI21_X1 _18494_ ( .A(_11560_ ), .B1(_11775_ ), .B2(_11776_ ), .ZN(_11777_ ) );
AOI221_X4 _18495_ ( .A(_11777_ ), .B1(\icache.icache_reg_1_3 [4] ), .B2(_11560_ ), .C1(_11576_ ), .C2(_11497_ ), .ZN(_11778_ ) );
AOI211_X1 _18496_ ( .A(\io_master_rdata [4] ), .B(_11301_ ), .C1(_11489_ ), .C2(_11493_ ), .ZN(_11779_ ) );
NOR3_X1 _18497_ ( .A1(_11778_ ), .A2(fanout_net_20 ), .A3(_11779_ ), .ZN(_00154_ ) );
OR3_X1 _18498_ ( .A1(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__A_Y ), .A2(\icache.icache_reg_1_3 [3] ), .A3(_11506_ ), .ZN(_11780_ ) );
MUX2_X1 _18499_ ( .A(\icache.icache_reg_0_0 [3] ), .B(\icache.icache_reg_0_1 [3] ), .S(_11512_ ), .Z(_11781_ ) );
MUX2_X1 _18500_ ( .A(\icache.icache_reg_0_2 [3] ), .B(_11781_ ), .S(_11549_ ), .Z(_11782_ ) );
MUX2_X1 _18501_ ( .A(\icache.icache_reg_0_3 [3] ), .B(_11782_ ), .S(_11553_ ), .Z(_11783_ ) );
MUX2_X1 _18502_ ( .A(\icache.icache_reg_1_0 [3] ), .B(_11783_ ), .S(_11612_ ), .Z(_11784_ ) );
MUX2_X1 _18503_ ( .A(\icache.icache_reg_1_1 [3] ), .B(_11784_ ), .S(_11529_ ), .Z(_11785_ ) );
MUX2_X1 _18504_ ( .A(\icache.icache_reg_1_2 [3] ), .B(_11785_ ), .S(_11534_ ), .Z(_11786_ ) );
OAI221_X1 _18505_ ( .A(_11780_ ), .B1(_11575_ ), .B2(_11786_ ), .C1(_11495_ ), .C2(_11580_ ), .ZN(_11787_ ) );
NAND3_X1 _18506_ ( .A1(_11577_ ), .A2(\io_master_rdata [3] ), .A3(_11578_ ), .ZN(_11788_ ) );
AOI21_X1 _18507_ ( .A(fanout_net_20 ), .B1(_11787_ ), .B2(_11788_ ), .ZN(_00155_ ) );
OR3_X1 _18508_ ( .A1(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__A_Y ), .A2(\icache.icache_reg_1_3 [2] ), .A3(_11506_ ), .ZN(_11789_ ) );
MUX2_X1 _18509_ ( .A(\icache.icache_reg_0_0 [2] ), .B(\icache.icache_reg_0_1 [2] ), .S(_11512_ ), .Z(_11790_ ) );
MUX2_X1 _18510_ ( .A(\icache.icache_reg_0_2 [2] ), .B(_11790_ ), .S(_11549_ ), .Z(_11791_ ) );
MUX2_X1 _18511_ ( .A(\icache.icache_reg_0_3 [2] ), .B(_11791_ ), .S(_11553_ ), .Z(_11792_ ) );
MUX2_X1 _18512_ ( .A(\icache.icache_reg_1_0 [2] ), .B(_11792_ ), .S(_11612_ ), .Z(_11793_ ) );
MUX2_X1 _18513_ ( .A(\icache.icache_reg_1_1 [2] ), .B(_11793_ ), .S(_11529_ ), .Z(_11794_ ) );
MUX2_X1 _18514_ ( .A(\icache.icache_reg_1_2 [2] ), .B(_11794_ ), .S(_11534_ ), .Z(_11795_ ) );
OAI221_X1 _18515_ ( .A(_11789_ ), .B1(_11575_ ), .B2(_11795_ ), .C1(_11495_ ), .C2(_11580_ ), .ZN(_11796_ ) );
NAND3_X1 _18516_ ( .A1(_11577_ ), .A2(\io_master_rdata [2] ), .A3(_11578_ ), .ZN(_11797_ ) );
AOI21_X1 _18517_ ( .A(fanout_net_20 ), .B1(_11796_ ), .B2(_11797_ ), .ZN(_00156_ ) );
AOI211_X1 _18518_ ( .A(\io_master_rdata [28] ), .B(_11648_ ), .C1(_11581_ ), .C2(_11583_ ), .ZN(_11798_ ) );
AND3_X1 _18519_ ( .A1(_10841_ ), .A2(\icache.icache_reg_1_3 [28] ), .A3(_11503_ ), .ZN(_11799_ ) );
MUX2_X1 _18520_ ( .A(\icache.icache_reg_0_0 [28] ), .B(\icache.icache_reg_0_1 [28] ), .S(_11513_ ), .Z(_11800_ ) );
MUX2_X1 _18521_ ( .A(\icache.icache_reg_0_2 [28] ), .B(_11800_ ), .S(_11550_ ), .Z(_11801_ ) );
MUX2_X1 _18522_ ( .A(\icache.icache_reg_0_3 [28] ), .B(_11801_ ), .S(_11554_ ), .Z(_11802_ ) );
MUX2_X1 _18523_ ( .A(\icache.icache_reg_1_0 [28] ), .B(_11802_ ), .S(_11525_ ), .Z(_11803_ ) );
MUX2_X1 _18524_ ( .A(\icache.icache_reg_1_1 [28] ), .B(_11803_ ), .S(_11530_ ), .Z(_11804_ ) );
MUX2_X1 _18525_ ( .A(\icache.icache_reg_1_2 [28] ), .B(_11804_ ), .S(_11535_ ), .Z(_11805_ ) );
AOI21_X1 _18526_ ( .A(_11799_ ), .B1(_11805_ ), .B2(_11540_ ), .ZN(_11806_ ) );
AOI211_X1 _18527_ ( .A(fanout_net_20 ), .B(_11798_ ), .C1(_11500_ ), .C2(_11806_ ), .ZN(_00157_ ) );
AND3_X1 _18528_ ( .A1(_11643_ ), .A2(\icache.icache_reg_1_3 [1] ), .A3(_11502_ ), .ZN(_11807_ ) );
NAND3_X1 _18529_ ( .A1(_11571_ ), .A2(\icache.icache_reg_1_1 [1] ), .A3(_11509_ ), .ZN(_11808_ ) );
AND3_X1 _18530_ ( .A1(_11505_ ), .A2(\icache.icache_reg_1_0 [1] ), .A3(_11523_ ), .ZN(_11809_ ) );
MUX2_X1 _18531_ ( .A(\icache.icache_reg_0_0 [1] ), .B(\icache.icache_reg_0_1 [1] ), .S(_11512_ ), .Z(_11810_ ) );
MUX2_X1 _18532_ ( .A(\icache.icache_reg_0_2 [1] ), .B(_11810_ ), .S(_11549_ ), .Z(_11811_ ) );
MUX2_X1 _18533_ ( .A(\icache.icache_reg_0_3 [1] ), .B(_11811_ ), .S(_11553_ ), .Z(_11812_ ) );
AOI21_X1 _18534_ ( .A(_11809_ ), .B1(_11812_ ), .B2(_11612_ ), .ZN(_11813_ ) );
OAI21_X1 _18535_ ( .A(_11808_ ), .B1(_11813_ ), .B2(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_NOR__A_Y ), .ZN(_11814_ ) );
MUX2_X1 _18536_ ( .A(\icache.icache_reg_1_2 [1] ), .B(_11814_ ), .S(_11533_ ), .Z(_11815_ ) );
AOI221_X4 _18537_ ( .A(_11807_ ), .B1(_11539_ ), .B2(_11815_ ), .C1(_11576_ ), .C2(_11497_ ), .ZN(_11816_ ) );
AOI211_X1 _18538_ ( .A(\io_master_rdata [1] ), .B(_11301_ ), .C1(_11489_ ), .C2(_11493_ ), .ZN(_11817_ ) );
NOR3_X1 _18539_ ( .A1(_11816_ ), .A2(fanout_net_20 ), .A3(_11817_ ), .ZN(_00158_ ) );
OR3_X1 _18540_ ( .A1(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__A_Y ), .A2(\icache.icache_reg_1_3 [0] ), .A3(_11506_ ), .ZN(_11818_ ) );
MUX2_X1 _18541_ ( .A(\icache.icache_reg_0_0 [0] ), .B(\icache.icache_reg_0_1 [0] ), .S(_11512_ ), .Z(_11819_ ) );
MUX2_X1 _18542_ ( .A(\icache.icache_reg_0_2 [0] ), .B(_11819_ ), .S(_11549_ ), .Z(_11820_ ) );
MUX2_X1 _18543_ ( .A(\icache.icache_reg_0_3 [0] ), .B(_11820_ ), .S(_11553_ ), .Z(_11821_ ) );
MUX2_X1 _18544_ ( .A(\icache.icache_reg_1_0 [0] ), .B(_11821_ ), .S(_11612_ ), .Z(_11822_ ) );
MUX2_X1 _18545_ ( .A(\icache.icache_reg_1_1 [0] ), .B(_11822_ ), .S(_11529_ ), .Z(_11823_ ) );
MUX2_X1 _18546_ ( .A(\icache.icache_reg_1_2 [0] ), .B(_11823_ ), .S(_11534_ ), .Z(_11824_ ) );
OAI221_X1 _18547_ ( .A(_11818_ ), .B1(_11575_ ), .B2(_11824_ ), .C1(_11495_ ), .C2(_11580_ ), .ZN(_11825_ ) );
NAND3_X1 _18548_ ( .A1(_11577_ ), .A2(\io_master_rdata [0] ), .A3(_11578_ ), .ZN(_11826_ ) );
AOI21_X1 _18549_ ( .A(fanout_net_20 ), .B1(_11825_ ), .B2(_11826_ ), .ZN(_00159_ ) );
AOI211_X1 _18550_ ( .A(\io_master_rdata [27] ), .B(_11648_ ), .C1(_11581_ ), .C2(_11583_ ), .ZN(_11827_ ) );
AND3_X1 _18551_ ( .A1(_10841_ ), .A2(\icache.icache_reg_1_3 [27] ), .A3(_11503_ ), .ZN(_11828_ ) );
MUX2_X1 _18552_ ( .A(\icache.icache_reg_0_0 [27] ), .B(\icache.icache_reg_0_1 [27] ), .S(_11513_ ), .Z(_11829_ ) );
MUX2_X1 _18553_ ( .A(\icache.icache_reg_0_2 [27] ), .B(_11829_ ), .S(_11550_ ), .Z(_11830_ ) );
MUX2_X1 _18554_ ( .A(\icache.icache_reg_0_3 [27] ), .B(_11830_ ), .S(_11554_ ), .Z(_11831_ ) );
MUX2_X1 _18555_ ( .A(\icache.icache_reg_1_0 [27] ), .B(_11831_ ), .S(_11525_ ), .Z(_11832_ ) );
MUX2_X1 _18556_ ( .A(\icache.icache_reg_1_1 [27] ), .B(_11832_ ), .S(_11530_ ), .Z(_11833_ ) );
MUX2_X1 _18557_ ( .A(\icache.icache_reg_1_2 [27] ), .B(_11833_ ), .S(_11535_ ), .Z(_11834_ ) );
AOI21_X1 _18558_ ( .A(_11828_ ), .B1(_11834_ ), .B2(_11540_ ), .ZN(_11835_ ) );
AOI211_X1 _18559_ ( .A(fanout_net_20 ), .B(_11827_ ), .C1(_11500_ ), .C2(_11835_ ), .ZN(_00160_ ) );
AOI211_X1 _18560_ ( .A(\io_master_rdata [26] ), .B(_11648_ ), .C1(_11581_ ), .C2(_11583_ ), .ZN(_11836_ ) );
AND3_X1 _18561_ ( .A1(_10841_ ), .A2(\icache.icache_reg_1_3 [26] ), .A3(_11502_ ), .ZN(_11837_ ) );
NAND3_X1 _18562_ ( .A1(_11643_ ), .A2(\icache.icache_reg_1_1 [26] ), .A3(_11509_ ), .ZN(_11838_ ) );
NAND3_X1 _18563_ ( .A1(_10836_ ), .A2(\icache.icache_reg_0_2 [26] ), .A3(_11518_ ), .ZN(_11839_ ) );
AND4_X1 _18564_ ( .A1(\icache.icache_reg_0_1 [26] ), .A2(_11561_ ), .A3(_11562_ ), .A4(_11509_ ), .ZN(_11840_ ) );
AOI21_X1 _18565_ ( .A(_11840_ ), .B1(_11714_ ), .B2(\icache.icache_reg_0_0 [26] ), .ZN(_11841_ ) );
OAI211_X1 _18566_ ( .A(_11567_ ), .B(_11839_ ), .C1(_11841_ ), .C2(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_ANDNOT__B_Y ), .ZN(_11842_ ) );
OR3_X1 _18567_ ( .A1(_10840_ ), .A2(\icache.icache_reg_0_3 [26] ), .A3(_11506_ ), .ZN(_11843_ ) );
AOI21_X1 _18568_ ( .A(\icache.offset_buf_$_OR__A_Y_$_NOR__A_Y ), .B1(_11842_ ), .B2(_11843_ ), .ZN(_11844_ ) );
AOI221_X4 _18569_ ( .A(\icache.offset_buf [1] ), .B1(\icache.icache_reg_1_0 [26] ), .B2(_11508_ ), .C1(_11561_ ), .C2(_11562_ ), .ZN(_11845_ ) );
OAI21_X1 _18570_ ( .A(_11838_ ), .B1(_11844_ ), .B2(_11845_ ), .ZN(_11846_ ) );
MUX2_X1 _18571_ ( .A(\icache.icache_reg_1_2 [26] ), .B(_11846_ ), .S(_11535_ ), .Z(_11847_ ) );
AOI21_X1 _18572_ ( .A(_11837_ ), .B1(_11847_ ), .B2(_11540_ ), .ZN(_11848_ ) );
AOI211_X1 _18573_ ( .A(fanout_net_20 ), .B(_11836_ ), .C1(_11500_ ), .C2(_11848_ ), .ZN(_00161_ ) );
AOI211_X1 _18574_ ( .A(\io_master_rdata [25] ), .B(_11648_ ), .C1(_11581_ ), .C2(_11583_ ), .ZN(_11849_ ) );
OR3_X1 _18575_ ( .A1(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__A_Y ), .A2(\icache.icache_reg_1_3 [25] ), .A3(_11506_ ), .ZN(_11850_ ) );
MUX2_X1 _18576_ ( .A(\icache.icache_reg_0_0 [25] ), .B(\icache.icache_reg_0_1 [25] ), .S(_11512_ ), .Z(_11851_ ) );
MUX2_X1 _18577_ ( .A(\icache.icache_reg_0_2 [25] ), .B(_11851_ ), .S(_11549_ ), .Z(_11852_ ) );
MUX2_X1 _18578_ ( .A(\icache.icache_reg_0_3 [25] ), .B(_11852_ ), .S(_11554_ ), .Z(_11853_ ) );
MUX2_X1 _18579_ ( .A(\icache.icache_reg_1_0 [25] ), .B(_11853_ ), .S(_11612_ ), .Z(_11854_ ) );
MUX2_X1 _18580_ ( .A(\icache.icache_reg_1_1 [25] ), .B(_11854_ ), .S(_11529_ ), .Z(_11855_ ) );
MUX2_X1 _18581_ ( .A(\icache.icache_reg_1_2 [25] ), .B(_11855_ ), .S(_11534_ ), .Z(_11856_ ) );
OAI21_X1 _18582_ ( .A(_11850_ ), .B1(_11856_ ), .B2(_11575_ ), .ZN(_11857_ ) );
AOI211_X1 _18583_ ( .A(fanout_net_20 ), .B(_11849_ ), .C1(_11499_ ), .C2(_11857_ ), .ZN(_00162_ ) );
AOI211_X1 _18584_ ( .A(\io_master_rdata [24] ), .B(_11648_ ), .C1(_11581_ ), .C2(_11583_ ), .ZN(_11858_ ) );
AND3_X1 _18585_ ( .A1(_10841_ ), .A2(\icache.icache_reg_1_3 [24] ), .A3(_11502_ ), .ZN(_11859_ ) );
MUX2_X1 _18586_ ( .A(\icache.icache_reg_0_0 [24] ), .B(\icache.icache_reg_0_1 [24] ), .S(_11513_ ), .Z(_11860_ ) );
MUX2_X1 _18587_ ( .A(\icache.icache_reg_0_2 [24] ), .B(_11860_ ), .S(_11550_ ), .Z(_11861_ ) );
MUX2_X1 _18588_ ( .A(\icache.icache_reg_0_3 [24] ), .B(_11861_ ), .S(_11554_ ), .Z(_11862_ ) );
MUX2_X1 _18589_ ( .A(\icache.icache_reg_1_0 [24] ), .B(_11862_ ), .S(_11612_ ), .Z(_11863_ ) );
MUX2_X1 _18590_ ( .A(\icache.icache_reg_1_1 [24] ), .B(_11863_ ), .S(_11530_ ), .Z(_11864_ ) );
MUX2_X1 _18591_ ( .A(\icache.icache_reg_1_2 [24] ), .B(_11864_ ), .S(_11535_ ), .Z(_11865_ ) );
AOI21_X1 _18592_ ( .A(_11859_ ), .B1(_11865_ ), .B2(_11540_ ), .ZN(_11866_ ) );
AOI211_X1 _18593_ ( .A(fanout_net_20 ), .B(_11858_ ), .C1(_11499_ ), .C2(_11866_ ), .ZN(_00163_ ) );
AOI211_X1 _18594_ ( .A(\icache.icache_reg_1_2 [23] ), .B(_11547_ ), .C1(_11561_ ), .C2(_11562_ ), .ZN(_11867_ ) );
NAND3_X1 _18595_ ( .A1(_11571_ ), .A2(\icache.icache_reg_1_0 [23] ), .A3(_11523_ ), .ZN(_11868_ ) );
AND4_X1 _18596_ ( .A1(\icache.icache_reg_0_3 [23] ), .A2(_09335_ ), .A3(_09337_ ), .A4(_11501_ ), .ZN(_11869_ ) );
MUX2_X1 _18597_ ( .A(\icache.icache_reg_0_0 [23] ), .B(\icache.icache_reg_0_1 [23] ), .S(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_ANDNOT__B_Y ), .Z(_11870_ ) );
MUX2_X1 _18598_ ( .A(\icache.icache_reg_0_2 [23] ), .B(_11870_ ), .S(_11550_ ), .Z(_11871_ ) );
AOI21_X1 _18599_ ( .A(_11869_ ), .B1(_11871_ ), .B2(_11567_ ), .ZN(_11872_ ) );
OAI211_X1 _18600_ ( .A(_11529_ ), .B(_11868_ ), .C1(_11872_ ), .C2(\icache.offset_buf_$_OR__A_Y_$_NOR__A_Y ), .ZN(_11873_ ) );
OAI21_X1 _18601_ ( .A(_11873_ ), .B1(\icache.icache_reg_1_1 [23] ), .B2(_11530_ ), .ZN(_11874_ ) );
AOI211_X1 _18602_ ( .A(_11560_ ), .B(_11867_ ), .C1(_11874_ ), .C2(_11534_ ), .ZN(_11875_ ) );
AOI221_X4 _18603_ ( .A(_11875_ ), .B1(\icache.icache_reg_1_3 [23] ), .B2(_11560_ ), .C1(_11576_ ), .C2(_11497_ ), .ZN(_11876_ ) );
AOI211_X1 _18604_ ( .A(\io_master_rdata [23] ), .B(_11301_ ), .C1(_11489_ ), .C2(_11493_ ), .ZN(_11877_ ) );
NOR3_X1 _18605_ ( .A1(_11876_ ), .A2(fanout_net_20 ), .A3(_11877_ ), .ZN(_00164_ ) );
AND3_X1 _18606_ ( .A1(_11572_ ), .A2(\icache.icache_reg_1_3 [22] ), .A3(_11501_ ), .ZN(_11878_ ) );
MUX2_X1 _18607_ ( .A(\icache.icache_reg_0_0 [22] ), .B(\icache.icache_reg_0_1 [22] ), .S(_11511_ ), .Z(_11879_ ) );
MUX2_X1 _18608_ ( .A(\icache.icache_reg_0_2 [22] ), .B(_11879_ ), .S(_11548_ ), .Z(_11880_ ) );
MUX2_X1 _18609_ ( .A(\icache.icache_reg_0_3 [22] ), .B(_11880_ ), .S(_11552_ ), .Z(_11881_ ) );
MUX2_X1 _18610_ ( .A(\icache.icache_reg_1_0 [22] ), .B(_11881_ ), .S(_11524_ ), .Z(_11882_ ) );
MUX2_X1 _18611_ ( .A(\icache.icache_reg_1_1 [22] ), .B(_11882_ ), .S(_11528_ ), .Z(_11883_ ) );
MUX2_X1 _18612_ ( .A(\icache.icache_reg_1_2 [22] ), .B(_11883_ ), .S(_11532_ ), .Z(_11884_ ) );
AOI221_X4 _18613_ ( .A(_11878_ ), .B1(_11538_ ), .B2(_11884_ ), .C1(_11576_ ), .C2(_11497_ ), .ZN(_11885_ ) );
INV_X1 _18614_ ( .A(\io_master_rdata [22] ), .ZN(_11886_ ) );
AOI211_X1 _18615_ ( .A(fanout_net_20 ), .B(_11885_ ), .C1(_11886_ ), .C2(_11498_ ), .ZN(_00165_ ) );
AND3_X1 _18616_ ( .A1(_10987_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [31] ), .ZN(_00166_ ) );
AND3_X1 _18617_ ( .A1(_10987_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [30] ), .ZN(_00167_ ) );
AND3_X1 _18618_ ( .A1(_10987_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [21] ), .ZN(_00168_ ) );
AND3_X1 _18619_ ( .A1(_10987_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [20] ), .ZN(_00169_ ) );
AND3_X1 _18620_ ( .A1(_10987_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [19] ), .ZN(_00170_ ) );
CLKBUF_X2 _18621_ ( .A(_10846_ ), .Z(_11887_ ) );
AND3_X1 _18622_ ( .A1(_11887_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [18] ), .ZN(_00171_ ) );
AND3_X1 _18623_ ( .A1(_11887_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [17] ), .ZN(_00172_ ) );
AND3_X1 _18624_ ( .A1(_11887_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [16] ), .ZN(_00173_ ) );
AND3_X1 _18625_ ( .A1(_11887_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [15] ), .ZN(_00174_ ) );
AND3_X1 _18626_ ( .A1(_11887_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [14] ), .ZN(_00175_ ) );
AND3_X1 _18627_ ( .A1(_11887_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [13] ), .ZN(_00176_ ) );
NAND2_X1 _18628_ ( .A1(fanout_net_2 ), .A2(\io_master_rdata [12] ), .ZN(_11888_ ) );
NOR2_X1 _18629_ ( .A1(_11888_ ), .A2(fanout_net_20 ), .ZN(_00177_ ) );
AND3_X1 _18630_ ( .A1(_11887_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [29] ), .ZN(_00178_ ) );
AND3_X1 _18631_ ( .A1(_11887_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [11] ), .ZN(_00179_ ) );
AND3_X1 _18632_ ( .A1(_11887_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [10] ), .ZN(_00180_ ) );
AND3_X1 _18633_ ( .A1(_11887_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [9] ), .ZN(_00181_ ) );
CLKBUF_X2 _18634_ ( .A(_10846_ ), .Z(_11889_ ) );
AND3_X1 _18635_ ( .A1(_11889_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [8] ), .ZN(_00182_ ) );
AND3_X1 _18636_ ( .A1(_11889_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [7] ), .ZN(_00183_ ) );
AND3_X1 _18637_ ( .A1(_11889_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [6] ), .ZN(_00184_ ) );
AND3_X1 _18638_ ( .A1(_11889_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [5] ), .ZN(_00185_ ) );
AND3_X1 _18639_ ( .A1(_11889_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [4] ), .ZN(_00186_ ) );
AND3_X1 _18640_ ( .A1(_11889_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [3] ), .ZN(_00187_ ) );
AND3_X1 _18641_ ( .A1(_11889_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [2] ), .ZN(_00188_ ) );
AND3_X1 _18642_ ( .A1(_11889_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [28] ), .ZN(_00189_ ) );
AND3_X1 _18643_ ( .A1(_11889_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [1] ), .ZN(_00190_ ) );
AND3_X1 _18644_ ( .A1(_11889_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [0] ), .ZN(_00191_ ) );
AND3_X1 _18645_ ( .A1(_10847_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [27] ), .ZN(_00192_ ) );
AND3_X1 _18646_ ( .A1(_10847_ ), .A2(fanout_net_2 ), .A3(\io_master_rdata [26] ), .ZN(_00193_ ) );
AND3_X1 _18647_ ( .A1(_10847_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [25] ), .ZN(_00194_ ) );
AND3_X1 _18648_ ( .A1(_10847_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [24] ), .ZN(_00195_ ) );
AND3_X1 _18649_ ( .A1(_10847_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [23] ), .ZN(_00196_ ) );
AND3_X1 _18650_ ( .A1(_10847_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [22] ), .ZN(_00197_ ) );
NAND2_X1 _18651_ ( .A1(fanout_net_3 ), .A2(io_master_rlast ), .ZN(_11890_ ) );
OAI211_X1 _18652_ ( .A(\icache.offset_buf_$_SDFFE_PP0P__Q_E ), .B(_11890_ ), .C1(_11518_ ), .C2(_11509_ ), .ZN(_11891_ ) );
NOR2_X1 _18653_ ( .A1(_11891_ ), .A2(fanout_net_20 ), .ZN(_00198_ ) );
BUF_X2 _18654_ ( .A(_10846_ ), .Z(_11892_ ) );
AND4_X1 _18655_ ( .A1(_11892_ ), .A2(\icache.offset_buf_$_SDFFE_PP0P__Q_E ), .A3(_11508_ ), .A4(_11890_ ), .ZN(_00199_ ) );
AOI21_X1 _18656_ ( .A(fanout_net_20 ), .B1(_09770_ ), .B2(_09771_ ), .ZN(_00200_ ) );
AOI21_X1 _18657_ ( .A(fanout_net_20 ), .B1(_09715_ ), .B2(_09716_ ), .ZN(_00201_ ) );
AND3_X1 _18658_ ( .A1(_09609_ ), .A2(_10992_ ), .A3(_09610_ ), .ZN(_00202_ ) );
AND3_X1 _18659_ ( .A1(_10054_ ), .A2(_10992_ ), .A3(_10056_ ), .ZN(_00203_ ) );
AND3_X1 _18660_ ( .A1(_09967_ ), .A2(_10992_ ), .A3(_09968_ ), .ZN(_00204_ ) );
AND3_X1 _18661_ ( .A1(_10010_ ), .A2(_10992_ ), .A3(_10012_ ), .ZN(_00205_ ) );
AND3_X1 _18662_ ( .A1(_10102_ ), .A2(_10992_ ), .A3(_10103_ ), .ZN(_00206_ ) );
AND3_X1 _18663_ ( .A1(_09915_ ), .A2(_10992_ ), .A3(_09917_ ), .ZN(_00207_ ) );
AND3_X1 _18664_ ( .A1(_09867_ ), .A2(_10992_ ), .A3(_09868_ ), .ZN(_00208_ ) );
CLKBUF_X2 _18665_ ( .A(_10846_ ), .Z(_11893_ ) );
AND3_X1 _18666_ ( .A1(_10150_ ), .A2(_11893_ ), .A3(_10152_ ), .ZN(_00209_ ) );
AND3_X1 _18667_ ( .A1(_10199_ ), .A2(_11893_ ), .A3(_10201_ ), .ZN(_00210_ ) );
AND3_X1 _18668_ ( .A1(_10388_ ), .A2(_11893_ ), .A3(_10389_ ), .ZN(_00211_ ) );
AOI21_X1 _18669_ ( .A(fanout_net_20 ), .B1(_09816_ ), .B2(_09817_ ), .ZN(_00212_ ) );
AND3_X1 _18670_ ( .A1(_10347_ ), .A2(_11893_ ), .A3(_10348_ ), .ZN(_00213_ ) );
AND3_X1 _18671_ ( .A1(_10248_ ), .A2(_11893_ ), .A3(_10249_ ), .ZN(_00214_ ) );
AND3_X1 _18672_ ( .A1(_10293_ ), .A2(_11893_ ), .A3(_10294_ ), .ZN(_00215_ ) );
AND3_X1 _18673_ ( .A1(_10559_ ), .A2(_11893_ ), .A3(_10560_ ), .ZN(_00216_ ) );
AND3_X1 _18674_ ( .A1(_10518_ ), .A2(_11893_ ), .A3(_10519_ ), .ZN(_00217_ ) );
AND3_X1 _18675_ ( .A1(_10431_ ), .A2(_11893_ ), .A3(_10432_ ), .ZN(_00218_ ) );
AND3_X1 _18676_ ( .A1(_10473_ ), .A2(_11893_ ), .A3(_10474_ ), .ZN(_00219_ ) );
AOI21_X1 _18677_ ( .A(fanout_net_20 ), .B1(_09404_ ), .B2(_09405_ ), .ZN(_00220_ ) );
AND3_X1 _18678_ ( .A1(_09468_ ), .A2(_10917_ ), .A3(_09469_ ), .ZN(_00221_ ) );
AND3_X1 _18679_ ( .A1(_09187_ ), .A2(_10917_ ), .A3(_09188_ ), .ZN(_00222_ ) );
AND3_X1 _18680_ ( .A1(_09330_ ), .A2(_10917_ ), .A3(_09331_ ), .ZN(_00223_ ) );
AOI21_X1 _18681_ ( .A(fanout_net_20 ), .B1(_09647_ ), .B2(_09649_ ), .ZN(_00224_ ) );
AND3_X1 _18682_ ( .A1(_09521_ ), .A2(_10917_ ), .A3(_09522_ ), .ZN(_00225_ ) );
AND3_X1 _18683_ ( .A1(_09561_ ), .A2(_10917_ ), .A3(_09562_ ), .ZN(_00226_ ) );
AND2_X1 _18684_ ( .A1(_10709_ ), .A2(\icache._icache_reg_T ), .ZN(_11894_ ) );
BUF_X4 _18685_ ( .A(_11894_ ), .Z(_11895_ ) );
AOI21_X1 _18686_ ( .A(_10705_ ), .B1(_11577_ ), .B2(_11895_ ), .ZN(_11896_ ) );
AND3_X1 _18687_ ( .A1(_10623_ ), .A2(\idu.io_in_valid ), .A3(_10648_ ), .ZN(_11897_ ) );
NOR3_X1 _18688_ ( .A1(_11896_ ), .A2(fanout_net_21 ), .A3(_11897_ ), .ZN(_00227_ ) );
AOI211_X1 _18689_ ( .A(fanout_net_21 ), .B(_10828_ ), .C1(_11543_ ), .C2(_10830_ ), .ZN(_00228_ ) );
AND2_X1 _18690_ ( .A1(_11361_ ), .A2(_11362_ ), .ZN(_11898_ ) );
CLKBUF_X2 _18691_ ( .A(_09040_ ), .Z(_11899_ ) );
AOI211_X1 _18692_ ( .A(fanout_net_21 ), .B(_11898_ ), .C1(_idu_io_in_bits_T ), .C2(_11899_ ), .ZN(_00229_ ) );
NOR3_X1 _18693_ ( .A1(_10712_ ), .A2(fanout_net_21 ), .A3(_10832_ ), .ZN(_00230_ ) );
NOR2_X1 _18694_ ( .A1(_09656_ ), .A2(_09823_ ), .ZN(_11900_ ) );
AND3_X2 _18695_ ( .A1(_11900_ ), .A2(_10705_ ), .A3(_10569_ ), .ZN(_11901_ ) );
BUF_X2 _18696_ ( .A(_11901_ ), .Z(_11902_ ) );
CLKBUF_X2 _18697_ ( .A(_10704_ ), .Z(_11903_ ) );
INV_X1 _18698_ ( .A(_11437_ ), .ZN(_11904_ ) );
INV_X1 _18699_ ( .A(_11479_ ), .ZN(_11905_ ) );
NOR4_X1 _18700_ ( .A1(_11904_ ), .A2(\icache.icache_reg_0_3 [31] ), .A3(_10837_ ), .A4(_11905_ ), .ZN(_11906_ ) );
AOI21_X1 _18701_ ( .A(_11905_ ), .B1(_11435_ ), .B2(_11436_ ), .ZN(_11907_ ) );
AND2_X2 _18702_ ( .A1(_11907_ ), .A2(_09870_ ), .ZN(_11908_ ) );
AND3_X2 _18703_ ( .A1(_11435_ ), .A2(_11905_ ), .A3(_11436_ ), .ZN(_11909_ ) );
AND2_X2 _18704_ ( .A1(_11909_ ), .A2(_09870_ ), .ZN(_11910_ ) );
BUF_X4 _18705_ ( .A(_11910_ ), .Z(_11911_ ) );
BUF_X4 _18706_ ( .A(_11911_ ), .Z(_11912_ ) );
AOI21_X1 _18707_ ( .A(_11908_ ), .B1(_11912_ ), .B2(_11514_ ), .ZN(_11913_ ) );
OAI21_X1 _18708_ ( .A(_11913_ ), .B1(\icache.icache_reg_0_0 [31] ), .B2(_11912_ ), .ZN(_11914_ ) );
OAI211_X1 _18709_ ( .A(_10834_ ), .B(_11479_ ), .C1(_11437_ ), .C2(\icache.icache_reg_0_2 [31] ), .ZN(_11915_ ) );
AOI21_X1 _18710_ ( .A(_11906_ ), .B1(_11914_ ), .B2(_11915_ ), .ZN(_11916_ ) );
AND2_X2 _18711_ ( .A1(_11480_ ), .A2(_09818_ ), .ZN(_11917_ ) );
INV_X1 _18712_ ( .A(_11917_ ), .ZN(_11918_ ) );
BUF_X4 _18713_ ( .A(_11918_ ), .Z(_11919_ ) );
MUX2_X1 _18714_ ( .A(\icache.icache_reg_1_0 [31] ), .B(_11916_ ), .S(_11919_ ), .Z(_11920_ ) );
AND2_X2 _18715_ ( .A1(_11909_ ), .A2(_09818_ ), .ZN(_11921_ ) );
INV_X1 _18716_ ( .A(_11921_ ), .ZN(_11922_ ) );
BUF_X4 _18717_ ( .A(_11922_ ), .Z(_11923_ ) );
MUX2_X1 _18718_ ( .A(\icache.icache_reg_1_1 [31] ), .B(_11920_ ), .S(_11923_ ), .Z(_11924_ ) );
AND2_X2 _18719_ ( .A1(_11907_ ), .A2(_10837_ ), .ZN(_11925_ ) );
INV_X1 _18720_ ( .A(_11925_ ), .ZN(_11926_ ) );
BUF_X4 _18721_ ( .A(_11926_ ), .Z(_11927_ ) );
MUX2_X1 _18722_ ( .A(\icache.icache_reg_1_2 [31] ), .B(_11924_ ), .S(_11927_ ), .Z(_11928_ ) );
AND2_X1 _18723_ ( .A1(_11437_ ), .A2(_11479_ ), .ZN(_11929_ ) );
AND2_X1 _18724_ ( .A1(_11929_ ), .A2(_10838_ ), .ZN(_11930_ ) );
BUF_X4 _18725_ ( .A(_11930_ ), .Z(_11931_ ) );
NOR2_X1 _18726_ ( .A1(_11928_ ), .A2(_11931_ ), .ZN(_11932_ ) );
BUF_X2 _18727_ ( .A(_11904_ ), .Z(_11933_ ) );
BUF_X2 _18728_ ( .A(_11933_ ), .Z(_11934_ ) );
BUF_X4 _18729_ ( .A(_11905_ ), .Z(_11935_ ) );
BUF_X2 _18730_ ( .A(_11935_ ), .Z(_11936_ ) );
NOR4_X1 _18731_ ( .A1(_11934_ ), .A2(\icache.icache_reg_1_3 [31] ), .A3(_10836_ ), .A4(_11936_ ), .ZN(_11937_ ) );
NOR2_X1 _18732_ ( .A1(_11932_ ), .A2(_11937_ ), .ZN(_11938_ ) );
NAND4_X1 _18733_ ( .A1(_11902_ ), .A2(fanout_net_13 ), .A3(_11903_ ), .A4(_11938_ ), .ZN(_11939_ ) );
BUF_X2 _18734_ ( .A(_11929_ ), .Z(_11940_ ) );
AND2_X1 _18735_ ( .A1(_11940_ ), .A2(_11894_ ), .ZN(_11941_ ) );
BUF_X2 _18736_ ( .A(_11941_ ), .Z(_11942_ ) );
AND3_X1 _18737_ ( .A1(_11942_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [31] ), .ZN(_11943_ ) );
INV_X1 _18738_ ( .A(_11894_ ), .ZN(_11944_ ) );
NOR2_X1 _18739_ ( .A1(_11929_ ), .A2(_11944_ ), .ZN(_11945_ ) );
BUF_X4 _18740_ ( .A(_11945_ ), .Z(_11946_ ) );
AOI21_X1 _18741_ ( .A(_11943_ ), .B1(_11938_ ), .B2(_11946_ ), .ZN(_11947_ ) );
OAI21_X1 _18742_ ( .A(_11939_ ), .B1(_10708_ ), .B2(_11947_ ), .ZN(_11948_ ) );
CLKBUF_X2 _18743_ ( .A(_10709_ ), .Z(_11949_ ) );
BUF_X2 _18744_ ( .A(_11949_ ), .Z(_11950_ ) );
NAND2_X1 _18745_ ( .A1(_11495_ ), .A2(_11950_ ), .ZN(_11951_ ) );
BUF_X4 _18746_ ( .A(_10710_ ), .Z(_11952_ ) );
AOI22_X1 _18747_ ( .A1(_11948_ ), .A2(_11951_ ), .B1(_11952_ ), .B2(\ifu.inst [31] ), .ZN(_11953_ ) );
INV_X1 _18748_ ( .A(_10433_ ), .ZN(_11954_ ) );
NAND4_X1 _18749_ ( .A1(_11482_ ), .A2(_11326_ ), .A3(_11954_ ), .A4(_11405_ ), .ZN(_11955_ ) );
INV_X1 _18750_ ( .A(_10475_ ), .ZN(_11956_ ) );
NAND4_X1 _18751_ ( .A1(_11956_ ), .A2(_11327_ ), .A3(_11484_ ), .A4(_11365_ ), .ZN(_11957_ ) );
AND4_X1 _18752_ ( .A1(_10153_ ), .A2(_11480_ ), .A3(_10199_ ), .A4(_10201_ ), .ZN(_11958_ ) );
NAND4_X1 _18753_ ( .A1(_11958_ ), .A2(_09870_ ), .A3(_11483_ ), .A4(_10349_ ), .ZN(_11959_ ) );
NOR3_X1 _18754_ ( .A1(_11955_ ), .A2(_11957_ ), .A3(_11959_ ), .ZN(_11960_ ) );
NAND3_X1 _18755_ ( .A1(_11960_ ), .A2(_09869_ ), .A3(_09918_ ), .ZN(_11961_ ) );
NAND2_X1 _18756_ ( .A1(_11317_ ), .A2(_11961_ ), .ZN(_11962_ ) );
AND3_X1 _18757_ ( .A1(_11962_ ), .A2(_10013_ ), .A3(_10057_ ), .ZN(_11963_ ) );
NAND4_X1 _18758_ ( .A1(_11963_ ), .A2(_11304_ ), .A3(_09969_ ), .A4(_10104_ ), .ZN(_11964_ ) );
NAND4_X1 _18759_ ( .A1(_11308_ ), .A2(_09189_ ), .A3(_09563_ ), .A4(_09650_ ), .ZN(_11965_ ) );
NOR2_X1 _18760_ ( .A1(_11964_ ), .A2(_11965_ ), .ZN(_11966_ ) );
OR3_X1 _18761_ ( .A1(\ifu.pc [31] ), .A2(\ifu.pc [30] ), .A3(\ifu.pc [29] ), .ZN(_11967_ ) );
OAI21_X1 _18762_ ( .A(_09609_ ), .B1(_09610_ ), .B2(_11967_ ), .ZN(_11968_ ) );
AND4_X1 _18763_ ( .A1(_09406_ ), .A2(_11966_ ), .A3(_11305_ ), .A4(_11968_ ), .ZN(_11969_ ) );
NAND2_X1 _18764_ ( .A1(_09712_ ), .A2(_09714_ ), .ZN(_11970_ ) );
OAI21_X1 _18765_ ( .A(_09775_ ), .B1(_09763_ ), .B2(_09768_ ), .ZN(_11971_ ) );
OAI21_X1 _18766_ ( .A(\ifu.pc [31] ), .B1(_09402_ ), .B2(exu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_11972_ ) );
AND2_X1 _18767_ ( .A1(_11971_ ), .A2(_11972_ ), .ZN(_11973_ ) );
NAND2_X1 _18768_ ( .A1(_09813_ ), .A2(_09815_ ), .ZN(_11974_ ) );
NAND3_X1 _18769_ ( .A1(_11970_ ), .A2(_11973_ ), .A3(_11974_ ), .ZN(_11975_ ) );
NAND2_X1 _18770_ ( .A1(_11975_ ), .A2(_09466_ ), .ZN(_11976_ ) );
AND2_X2 _18771_ ( .A1(_11969_ ), .A2(_11976_ ), .ZN(_11977_ ) );
NAND4_X1 _18772_ ( .A1(_11977_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [31] ), .A4(_11950_ ), .ZN(_11978_ ) );
NAND2_X1 _18773_ ( .A1(_11953_ ), .A2(_11978_ ), .ZN(\ifu.io_out_bits_inst [31] ) );
AOI21_X1 _18774_ ( .A(fanout_net_21 ), .B1(_11953_ ), .B2(_11978_ ), .ZN(_00231_ ) );
AND4_X1 _18775_ ( .A1(_09969_ ), .A2(_11963_ ), .A3(_10104_ ), .A4(_09650_ ), .ZN(_11979_ ) );
AOI221_X4 _18776_ ( .A(_09611_ ), .B1(_09609_ ), .B2(_11967_ ), .C1(_09561_ ), .C2(_09562_ ), .ZN(_11980_ ) );
AND4_X1 _18777_ ( .A1(_11304_ ), .A2(_11979_ ), .A3(_11308_ ), .A4(_11980_ ), .ZN(_11981_ ) );
AND4_X2 _18778_ ( .A1(_09406_ ), .A2(_11981_ ), .A3(_11305_ ), .A4(_09189_ ), .ZN(_11982_ ) );
CLKBUF_X2 _18779_ ( .A(_11982_ ), .Z(_11983_ ) );
CLKBUF_X2 _18780_ ( .A(_11976_ ), .Z(_11984_ ) );
AND2_X1 _18781_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [30] ), .ZN(_11985_ ) );
AND4_X1 _18782_ ( .A1(_11950_ ), .A2(_11983_ ), .A3(_11984_ ), .A4(_11985_ ), .ZN(_11986_ ) );
BUF_X4 _18783_ ( .A(_10710_ ), .Z(_11987_ ) );
AOI21_X1 _18784_ ( .A(_11986_ ), .B1(_11987_ ), .B2(\ifu.inst [30] ), .ZN(_11988_ ) );
NAND2_X1 _18785_ ( .A1(_11977_ ), .A2(_11949_ ), .ZN(_11989_ ) );
BUF_X4 _18786_ ( .A(_11989_ ), .Z(_11990_ ) );
BUF_X4 _18787_ ( .A(_10706_ ), .Z(_11991_ ) );
NAND3_X1 _18788_ ( .A1(_11940_ ), .A2(_11985_ ), .A3(_11895_ ), .ZN(_11992_ ) );
BUF_X2 _18789_ ( .A(_11437_ ), .Z(_11993_ ) );
BUF_X2 _18790_ ( .A(_11993_ ), .Z(_11994_ ) );
BUF_X2 _18791_ ( .A(_11479_ ), .Z(_11995_ ) );
BUF_X2 _18792_ ( .A(_11995_ ), .Z(_11996_ ) );
BUF_X2 _18793_ ( .A(_11996_ ), .Z(_11997_ ) );
AND4_X1 _18794_ ( .A1(\icache.icache_reg_1_3 [30] ), .A2(_11994_ ), .A3(_11571_ ), .A4(_11997_ ), .ZN(_11998_ ) );
MUX2_X1 _18795_ ( .A(\icache.icache_reg_0_0 [30] ), .B(\icache.icache_reg_0_1 [30] ), .S(_11911_ ), .Z(_11999_ ) );
INV_X2 _18796_ ( .A(_11908_ ), .ZN(_12000_ ) );
BUF_X4 _18797_ ( .A(_12000_ ), .Z(_12001_ ) );
MUX2_X1 _18798_ ( .A(\icache.icache_reg_0_2 [30] ), .B(_11999_ ), .S(_12001_ ), .Z(_12002_ ) );
AND2_X1 _18799_ ( .A1(_11929_ ), .A2(_09870_ ), .ZN(_12003_ ) );
BUF_X4 _18800_ ( .A(_12003_ ), .Z(_12004_ ) );
INV_X2 _18801_ ( .A(_12004_ ), .ZN(_12005_ ) );
BUF_X4 _18802_ ( .A(_12005_ ), .Z(_12006_ ) );
MUX2_X1 _18803_ ( .A(\icache.icache_reg_0_3 [30] ), .B(_12002_ ), .S(_12006_ ), .Z(_12007_ ) );
MUX2_X1 _18804_ ( .A(\icache.icache_reg_1_0 [30] ), .B(_12007_ ), .S(_11919_ ), .Z(_12008_ ) );
MUX2_X1 _18805_ ( .A(\icache.icache_reg_1_1 [30] ), .B(_12008_ ), .S(_11923_ ), .Z(_12009_ ) );
MUX2_X1 _18806_ ( .A(\icache.icache_reg_1_2 [30] ), .B(_12009_ ), .S(_11927_ ), .Z(_12010_ ) );
INV_X1 _18807_ ( .A(_11930_ ), .ZN(_12011_ ) );
BUF_X4 _18808_ ( .A(_12011_ ), .Z(_12012_ ) );
AOI21_X1 _18809_ ( .A(_11998_ ), .B1(_12010_ ), .B2(_12012_ ), .ZN(_12013_ ) );
INV_X1 _18810_ ( .A(_11945_ ), .ZN(_12014_ ) );
OR2_X1 _18811_ ( .A1(_12013_ ), .A2(_12014_ ), .ZN(_12015_ ) );
AOI22_X1 _18812_ ( .A1(_11991_ ), .A2(fanout_net_13 ), .B1(_11992_ ), .B2(_12015_ ), .ZN(_12016_ ) );
NAND3_X1 _18813_ ( .A1(_11900_ ), .A2(_10705_ ), .A3(_10569_ ), .ZN(_12017_ ) );
INV_X1 _18814_ ( .A(fanout_net_13 ), .ZN(_12018_ ) );
BUF_X4 _18815_ ( .A(_12018_ ), .Z(_12019_ ) );
BUF_X4 _18816_ ( .A(_10703_ ), .Z(_12020_ ) );
NOR4_X1 _18817_ ( .A1(_12017_ ), .A2(_12019_ ), .A3(_12020_ ), .A4(_12013_ ), .ZN(_12021_ ) );
OAI21_X1 _18818_ ( .A(_11990_ ), .B1(_12016_ ), .B2(_12021_ ), .ZN(_12022_ ) );
NAND2_X1 _18819_ ( .A1(_11988_ ), .A2(_12022_ ), .ZN(\ifu.io_out_bits_inst [30] ) );
AOI21_X1 _18820_ ( .A(fanout_net_21 ), .B1(_11988_ ), .B2(_12022_ ), .ZN(_00232_ ) );
CLKBUF_X2 _18821_ ( .A(_11949_ ), .Z(_12023_ ) );
AND2_X1 _18822_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [21] ), .ZN(_12024_ ) );
AND4_X1 _18823_ ( .A1(_12023_ ), .A2(_11983_ ), .A3(_11984_ ), .A4(_12024_ ), .ZN(_12025_ ) );
AOI21_X1 _18824_ ( .A(_12025_ ), .B1(_11987_ ), .B2(\ifu.inst [21] ), .ZN(_12026_ ) );
NAND3_X1 _18825_ ( .A1(_11940_ ), .A2(_12024_ ), .A3(_11895_ ), .ZN(_12027_ ) );
OR4_X1 _18826_ ( .A1(\icache.icache_reg_0_2 [21] ), .A2(_11437_ ), .A3(_10837_ ), .A4(_11905_ ), .ZN(_12028_ ) );
MUX2_X1 _18827_ ( .A(\icache.icache_reg_0_0 [21] ), .B(\icache.icache_reg_0_1 [21] ), .S(_11912_ ), .Z(_12029_ ) );
OAI211_X1 _18828_ ( .A(_12006_ ), .B(_12028_ ), .C1(_12029_ ), .C2(_11908_ ), .ZN(_12030_ ) );
NAND4_X1 _18829_ ( .A1(_11437_ ), .A2(\icache.icache_reg_0_3 [21] ), .A3(_11515_ ), .A4(_11479_ ), .ZN(_12031_ ) );
NAND3_X1 _18830_ ( .A1(_12030_ ), .A2(_11919_ ), .A3(_12031_ ), .ZN(_12032_ ) );
NOR2_X1 _18831_ ( .A1(_11919_ ), .A2(\icache.icache_reg_1_0 [21] ), .ZN(_12033_ ) );
NOR2_X1 _18832_ ( .A1(_12033_ ), .A2(_11921_ ), .ZN(_12034_ ) );
AOI221_X4 _18833_ ( .A(_11925_ ), .B1(\icache.icache_reg_1_1 [21] ), .B2(_11921_ ), .C1(_12032_ ), .C2(_12034_ ), .ZN(_12035_ ) );
BUF_X2 _18834_ ( .A(_11993_ ), .Z(_12036_ ) );
BUF_X2 _18835_ ( .A(_11515_ ), .Z(_12037_ ) );
NOR4_X1 _18836_ ( .A1(_12036_ ), .A2(\icache.icache_reg_1_2 [21] ), .A3(_12037_ ), .A4(_11935_ ), .ZN(_12038_ ) );
NOR3_X1 _18837_ ( .A1(_12035_ ), .A2(_11931_ ), .A3(_12038_ ), .ZN(_12039_ ) );
AOI21_X1 _18838_ ( .A(_12039_ ), .B1(\icache.icache_reg_1_3 [21] ), .B2(_11931_ ), .ZN(_12040_ ) );
OR2_X1 _18839_ ( .A1(_12040_ ), .A2(_12014_ ), .ZN(_12041_ ) );
AOI22_X1 _18840_ ( .A1(_11991_ ), .A2(fanout_net_13 ), .B1(_12027_ ), .B2(_12041_ ), .ZN(_12042_ ) );
NOR4_X1 _18841_ ( .A1(_12017_ ), .A2(_12019_ ), .A3(_12020_ ), .A4(_12040_ ), .ZN(_12043_ ) );
OAI21_X1 _18842_ ( .A(_11990_ ), .B1(_12042_ ), .B2(_12043_ ), .ZN(_12044_ ) );
NAND2_X1 _18843_ ( .A1(_12026_ ), .A2(_12044_ ), .ZN(\ifu.io_out_bits_inst [21] ) );
AOI21_X1 _18844_ ( .A(fanout_net_21 ), .B1(_12026_ ), .B2(_12044_ ), .ZN(_00233_ ) );
AND2_X1 _18845_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [20] ), .ZN(_12045_ ) );
AND4_X1 _18846_ ( .A1(_12023_ ), .A2(_11983_ ), .A3(_11984_ ), .A4(_12045_ ), .ZN(_12046_ ) );
AOI21_X1 _18847_ ( .A(_12046_ ), .B1(_11987_ ), .B2(\ifu.inst [20] ), .ZN(_12047_ ) );
CLKBUF_X2 _18848_ ( .A(_10704_ ), .Z(_12048_ ) );
MUX2_X1 _18849_ ( .A(\icache.icache_reg_0_0 [20] ), .B(\icache.icache_reg_0_1 [20] ), .S(_11911_ ), .Z(_12049_ ) );
MUX2_X1 _18850_ ( .A(\icache.icache_reg_0_2 [20] ), .B(_12049_ ), .S(_12000_ ), .Z(_12050_ ) );
MUX2_X1 _18851_ ( .A(\icache.icache_reg_0_3 [20] ), .B(_12050_ ), .S(_12005_ ), .Z(_12051_ ) );
BUF_X4 _18852_ ( .A(_11918_ ), .Z(_12052_ ) );
MUX2_X1 _18853_ ( .A(\icache.icache_reg_1_0 [20] ), .B(_12051_ ), .S(_12052_ ), .Z(_12053_ ) );
BUF_X4 _18854_ ( .A(_11922_ ), .Z(_12054_ ) );
MUX2_X1 _18855_ ( .A(\icache.icache_reg_1_1 [20] ), .B(_12053_ ), .S(_12054_ ), .Z(_12055_ ) );
BUF_X4 _18856_ ( .A(_11926_ ), .Z(_12056_ ) );
MUX2_X1 _18857_ ( .A(\icache.icache_reg_1_2 [20] ), .B(_12055_ ), .S(_12056_ ), .Z(_12057_ ) );
MUX2_X1 _18858_ ( .A(\icache.icache_reg_1_3 [20] ), .B(_12057_ ), .S(_12012_ ), .Z(_12058_ ) );
AND4_X1 _18859_ ( .A1(fanout_net_13 ), .A2(_11902_ ), .A3(_12048_ ), .A4(_12058_ ), .ZN(_12059_ ) );
BUF_X4 _18860_ ( .A(_11941_ ), .Z(_12060_ ) );
AOI22_X1 _18861_ ( .A1(_12058_ ), .A2(_11946_ ), .B1(_12045_ ), .B2(_12060_ ), .ZN(_12061_ ) );
AOI21_X1 _18862_ ( .A(_12061_ ), .B1(_11991_ ), .B2(fanout_net_13 ), .ZN(_12062_ ) );
OAI21_X1 _18863_ ( .A(_11990_ ), .B1(_12059_ ), .B2(_12062_ ), .ZN(_12063_ ) );
NAND2_X1 _18864_ ( .A1(_12047_ ), .A2(_12063_ ), .ZN(\ifu.io_out_bits_inst [20] ) );
AOI21_X1 _18865_ ( .A(fanout_net_21 ), .B1(_12047_ ), .B2(_12063_ ), .ZN(_00234_ ) );
AND2_X1 _18866_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [19] ), .ZN(_12064_ ) );
AND4_X1 _18867_ ( .A1(_12023_ ), .A2(_11983_ ), .A3(_11984_ ), .A4(_12064_ ), .ZN(_12065_ ) );
AOI21_X1 _18868_ ( .A(_12065_ ), .B1(_11987_ ), .B2(\ifu.inst [19] ), .ZN(_12066_ ) );
NAND4_X1 _18869_ ( .A1(_11994_ ), .A2(\icache.icache_reg_1_3 [19] ), .A3(_11572_ ), .A4(_11997_ ), .ZN(_12067_ ) );
NAND4_X1 _18870_ ( .A1(_11934_ ), .A2(\icache.icache_reg_1_0 [19] ), .A3(_10839_ ), .A4(_11936_ ), .ZN(_12068_ ) );
OR4_X1 _18871_ ( .A1(\icache.icache_reg_0_1 [19] ), .A2(_11933_ ), .A3(_10837_ ), .A4(_11479_ ), .ZN(_12069_ ) );
BUF_X4 _18872_ ( .A(_12001_ ), .Z(_12070_ ) );
BUF_X4 _18873_ ( .A(_11912_ ), .Z(_12071_ ) );
OAI211_X1 _18874_ ( .A(_12069_ ), .B(_12070_ ), .C1(\icache.icache_reg_0_0 [19] ), .C2(_12071_ ), .ZN(_12072_ ) );
BUF_X2 _18875_ ( .A(_12006_ ), .Z(_12073_ ) );
BUF_X2 _18876_ ( .A(_11907_ ), .Z(_12074_ ) );
NAND3_X1 _18877_ ( .A1(_12074_ ), .A2(\icache.icache_reg_0_2 [19] ), .A3(_10835_ ), .ZN(_12075_ ) );
AND3_X1 _18878_ ( .A1(_12072_ ), .A2(_12073_ ), .A3(_12075_ ), .ZN(_12076_ ) );
OAI21_X1 _18879_ ( .A(_11919_ ), .B1(_12073_ ), .B2(\icache.icache_reg_0_3 [19] ), .ZN(_12077_ ) );
OAI211_X1 _18880_ ( .A(_11923_ ), .B(_12068_ ), .C1(_12076_ ), .C2(_12077_ ), .ZN(_12078_ ) );
OR4_X1 _18881_ ( .A1(\icache.icache_reg_1_1 [19] ), .A2(_11934_ ), .A3(_12037_ ), .A4(_11996_ ), .ZN(_12079_ ) );
AOI21_X1 _18882_ ( .A(_11925_ ), .B1(_12078_ ), .B2(_12079_ ), .ZN(_12080_ ) );
AOI211_X1 _18883_ ( .A(_10836_ ), .B(_11936_ ), .C1(_11934_ ), .C2(\icache.icache_reg_1_2 [19] ), .ZN(_12081_ ) );
OAI21_X1 _18884_ ( .A(_12067_ ), .B1(_12080_ ), .B2(_12081_ ), .ZN(_12082_ ) );
AND4_X1 _18885_ ( .A1(fanout_net_13 ), .A2(_11902_ ), .A3(_12048_ ), .A4(_12082_ ), .ZN(_12083_ ) );
AOI22_X1 _18886_ ( .A1(_12082_ ), .A2(_11946_ ), .B1(_12064_ ), .B2(_12060_ ), .ZN(_12084_ ) );
AOI21_X1 _18887_ ( .A(_12084_ ), .B1(_11991_ ), .B2(fanout_net_13 ), .ZN(_12085_ ) );
OAI21_X1 _18888_ ( .A(_11990_ ), .B1(_12083_ ), .B2(_12085_ ), .ZN(_12086_ ) );
NAND2_X1 _18889_ ( .A1(_12066_ ), .A2(_12086_ ), .ZN(\ifu.io_out_bits_inst [19] ) );
AOI21_X1 _18890_ ( .A(fanout_net_21 ), .B1(_12066_ ), .B2(_12086_ ), .ZN(_00235_ ) );
AND2_X1 _18891_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [18] ), .ZN(_12087_ ) );
AND4_X1 _18892_ ( .A1(_12023_ ), .A2(_11983_ ), .A3(_11984_ ), .A4(_12087_ ), .ZN(_12088_ ) );
AOI21_X1 _18893_ ( .A(_12088_ ), .B1(_11987_ ), .B2(\ifu.inst [18] ), .ZN(_12089_ ) );
AND2_X1 _18894_ ( .A1(_11982_ ), .A2(_11976_ ), .ZN(_12090_ ) );
NAND2_X1 _18895_ ( .A1(_12090_ ), .A2(_11950_ ), .ZN(_12091_ ) );
BUF_X2 _18896_ ( .A(_10706_ ), .Z(_12092_ ) );
AND4_X1 _18897_ ( .A1(_11607_ ), .A2(_11994_ ), .A3(_10840_ ), .A4(_11997_ ), .ZN(_12093_ ) );
NAND4_X1 _18898_ ( .A1(_11934_ ), .A2(\icache.icache_reg_1_0 [18] ), .A3(_10839_ ), .A4(_11936_ ), .ZN(_12094_ ) );
INV_X1 _18899_ ( .A(_11912_ ), .ZN(_12095_ ) );
OR2_X1 _18900_ ( .A1(_12095_ ), .A2(\icache.icache_reg_0_1 [18] ), .ZN(_12096_ ) );
OAI211_X1 _18901_ ( .A(_12096_ ), .B(_12070_ ), .C1(\icache.icache_reg_0_0 [18] ), .C2(_12071_ ), .ZN(_12097_ ) );
NAND3_X1 _18902_ ( .A1(_12074_ ), .A2(\icache.icache_reg_0_2 [18] ), .A3(_10835_ ), .ZN(_12098_ ) );
AND3_X1 _18903_ ( .A1(_12097_ ), .A2(_12073_ ), .A3(_12098_ ), .ZN(_12099_ ) );
OAI21_X1 _18904_ ( .A(_11919_ ), .B1(_12073_ ), .B2(\icache.icache_reg_0_3 [18] ), .ZN(_12100_ ) );
OAI211_X1 _18905_ ( .A(_11923_ ), .B(_12094_ ), .C1(_12099_ ), .C2(_12100_ ), .ZN(_12101_ ) );
BUF_X4 _18906_ ( .A(_11927_ ), .Z(_12102_ ) );
OR4_X1 _18907_ ( .A1(\icache.icache_reg_1_1 [18] ), .A2(_11934_ ), .A3(_12037_ ), .A4(_11996_ ), .ZN(_12103_ ) );
NAND3_X1 _18908_ ( .A1(_12101_ ), .A2(_12102_ ), .A3(_12103_ ), .ZN(_12104_ ) );
OAI211_X1 _18909_ ( .A(_10840_ ), .B(_11997_ ), .C1(_11994_ ), .C2(\icache.icache_reg_1_2 [18] ), .ZN(_12105_ ) );
AOI21_X1 _18910_ ( .A(_12093_ ), .B1(_12104_ ), .B2(_12105_ ), .ZN(_12106_ ) );
AND3_X1 _18911_ ( .A1(_12092_ ), .A2(fanout_net_13 ), .A3(_12106_ ), .ZN(_12107_ ) );
AOI22_X1 _18912_ ( .A1(_12106_ ), .A2(_11946_ ), .B1(_12087_ ), .B2(_12060_ ), .ZN(_12108_ ) );
BUF_X4 _18913_ ( .A(_10706_ ), .Z(_12109_ ) );
AOI21_X1 _18914_ ( .A(_12108_ ), .B1(_12109_ ), .B2(fanout_net_13 ), .ZN(_12110_ ) );
OAI21_X1 _18915_ ( .A(_12091_ ), .B1(_12107_ ), .B2(_12110_ ), .ZN(_12111_ ) );
NAND2_X1 _18916_ ( .A1(_12089_ ), .A2(_12111_ ), .ZN(\ifu.io_out_bits_inst [18] ) );
AOI21_X1 _18917_ ( .A(fanout_net_21 ), .B1(_12089_ ), .B2(_12111_ ), .ZN(_00236_ ) );
BUF_X4 _18918_ ( .A(_11917_ ), .Z(_12112_ ) );
AND4_X1 _18919_ ( .A1(\icache.icache_reg_0_3 [17] ), .A2(_11993_ ), .A3(_10835_ ), .A4(_11995_ ), .ZN(_12113_ ) );
MUX2_X1 _18920_ ( .A(\icache.icache_reg_0_0 [17] ), .B(\icache.icache_reg_0_1 [17] ), .S(_12071_ ), .Z(_12114_ ) );
MUX2_X1 _18921_ ( .A(\icache.icache_reg_0_2 [17] ), .B(_12114_ ), .S(_12070_ ), .Z(_12115_ ) );
AOI211_X1 _18922_ ( .A(_12112_ ), .B(_12113_ ), .C1(_12115_ ), .C2(_12073_ ), .ZN(_12116_ ) );
BUF_X4 _18923_ ( .A(_11921_ ), .Z(_12117_ ) );
NOR4_X1 _18924_ ( .A1(_12036_ ), .A2(\icache.icache_reg_1_0 [17] ), .A3(_12037_ ), .A4(_11996_ ), .ZN(_12118_ ) );
NOR3_X1 _18925_ ( .A1(_12116_ ), .A2(_12117_ ), .A3(_12118_ ), .ZN(_12119_ ) );
NAND3_X1 _18926_ ( .A1(_11909_ ), .A2(\icache.icache_reg_1_1 [17] ), .A3(_10840_ ), .ZN(_12120_ ) );
NAND2_X1 _18927_ ( .A1(_12102_ ), .A2(_12120_ ), .ZN(_12121_ ) );
OAI221_X1 _18928_ ( .A(_12012_ ), .B1(\icache.icache_reg_1_2 [17] ), .B2(_12102_ ), .C1(_12119_ ), .C2(_12121_ ), .ZN(_12122_ ) );
NAND4_X1 _18929_ ( .A1(_11994_ ), .A2(\icache.icache_reg_1_3 [17] ), .A3(_11643_ ), .A4(_11997_ ), .ZN(_12123_ ) );
NAND2_X1 _18930_ ( .A1(_12122_ ), .A2(_12123_ ), .ZN(_12124_ ) );
NAND4_X1 _18931_ ( .A1(_11902_ ), .A2(fanout_net_13 ), .A3(_11903_ ), .A4(_12124_ ), .ZN(_12125_ ) );
AND3_X1 _18932_ ( .A1(_11942_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [17] ), .ZN(_12126_ ) );
AOI21_X1 _18933_ ( .A(_12126_ ), .B1(_12124_ ), .B2(_11946_ ), .ZN(_12127_ ) );
OAI21_X1 _18934_ ( .A(_12125_ ), .B1(_10708_ ), .B2(_12127_ ), .ZN(_12128_ ) );
AOI22_X1 _18935_ ( .A1(_12128_ ), .A2(_11951_ ), .B1(_11952_ ), .B2(\ifu.inst [17] ), .ZN(_12129_ ) );
NAND4_X1 _18936_ ( .A1(_11977_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [17] ), .A4(_11950_ ), .ZN(_12130_ ) );
NAND2_X1 _18937_ ( .A1(_12129_ ), .A2(_12130_ ), .ZN(\ifu.io_out_bits_inst [17] ) );
AOI21_X1 _18938_ ( .A(fanout_net_21 ), .B1(_12129_ ), .B2(_12130_ ), .ZN(_00237_ ) );
AND2_X1 _18939_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [16] ), .ZN(_12131_ ) );
AND4_X1 _18940_ ( .A1(_12023_ ), .A2(_11983_ ), .A3(_11984_ ), .A4(_12131_ ), .ZN(_12132_ ) );
AOI21_X1 _18941_ ( .A(_12132_ ), .B1(_11987_ ), .B2(\ifu.inst [16] ), .ZN(_12133_ ) );
NOR4_X1 _18942_ ( .A1(_12036_ ), .A2(\icache.icache_reg_1_2 [16] ), .A3(_12037_ ), .A4(_11936_ ), .ZN(_12134_ ) );
NOR4_X1 _18943_ ( .A1(_11993_ ), .A2(\icache.icache_reg_1_0 [16] ), .A3(_11515_ ), .A4(_11995_ ), .ZN(_12135_ ) );
NOR2_X1 _18944_ ( .A1(_12135_ ), .A2(_11921_ ), .ZN(_12136_ ) );
MUX2_X1 _18945_ ( .A(\icache.icache_reg_0_0 [16] ), .B(\icache.icache_reg_0_1 [16] ), .S(_11912_ ), .Z(_12137_ ) );
MUX2_X1 _18946_ ( .A(\icache.icache_reg_0_2 [16] ), .B(_12137_ ), .S(_12001_ ), .Z(_12138_ ) );
MUX2_X1 _18947_ ( .A(\icache.icache_reg_0_3 [16] ), .B(_12138_ ), .S(_12073_ ), .Z(_12139_ ) );
OAI21_X1 _18948_ ( .A(_12136_ ), .B1(_12139_ ), .B2(_12112_ ), .ZN(_12140_ ) );
AOI21_X1 _18949_ ( .A(_11925_ ), .B1(_12117_ ), .B2(\icache.icache_reg_1_1 [16] ), .ZN(_12141_ ) );
AOI21_X1 _18950_ ( .A(_12134_ ), .B1(_12140_ ), .B2(_12141_ ), .ZN(_12142_ ) );
BUF_X4 _18951_ ( .A(_12011_ ), .Z(_12143_ ) );
MUX2_X1 _18952_ ( .A(\icache.icache_reg_1_3 [16] ), .B(_12142_ ), .S(_12143_ ), .Z(_12144_ ) );
AND4_X1 _18953_ ( .A1(fanout_net_13 ), .A2(_11902_ ), .A3(_12048_ ), .A4(_12144_ ), .ZN(_12145_ ) );
AOI22_X1 _18954_ ( .A1(_12144_ ), .A2(_11946_ ), .B1(_12131_ ), .B2(_12060_ ), .ZN(_12146_ ) );
AOI21_X1 _18955_ ( .A(_12146_ ), .B1(_12109_ ), .B2(fanout_net_13 ), .ZN(_12147_ ) );
OAI21_X1 _18956_ ( .A(_11990_ ), .B1(_12145_ ), .B2(_12147_ ), .ZN(_12148_ ) );
NAND2_X1 _18957_ ( .A1(_12133_ ), .A2(_12148_ ), .ZN(\ifu.io_out_bits_inst [16] ) );
AOI21_X1 _18958_ ( .A(fanout_net_21 ), .B1(_12133_ ), .B2(_12148_ ), .ZN(_00238_ ) );
AND2_X1 _18959_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [15] ), .ZN(_12149_ ) );
AND4_X1 _18960_ ( .A1(_12023_ ), .A2(_11983_ ), .A3(_11984_ ), .A4(_12149_ ), .ZN(_12150_ ) );
AOI21_X1 _18961_ ( .A(_12150_ ), .B1(_11987_ ), .B2(\ifu.inst [15] ), .ZN(_12151_ ) );
MUX2_X1 _18962_ ( .A(\icache.icache_reg_0_0 [15] ), .B(\icache.icache_reg_0_1 [15] ), .S(_11910_ ), .Z(_12152_ ) );
MUX2_X1 _18963_ ( .A(\icache.icache_reg_0_2 [15] ), .B(_12152_ ), .S(_12000_ ), .Z(_12153_ ) );
MUX2_X1 _18964_ ( .A(\icache.icache_reg_0_3 [15] ), .B(_12153_ ), .S(_12005_ ), .Z(_12154_ ) );
MUX2_X1 _18965_ ( .A(\icache.icache_reg_1_0 [15] ), .B(_12154_ ), .S(_12052_ ), .Z(_12155_ ) );
MUX2_X1 _18966_ ( .A(\icache.icache_reg_1_1 [15] ), .B(_12155_ ), .S(_12054_ ), .Z(_12156_ ) );
MUX2_X1 _18967_ ( .A(\icache.icache_reg_1_2 [15] ), .B(_12156_ ), .S(_12056_ ), .Z(_12157_ ) );
MUX2_X1 _18968_ ( .A(\icache.icache_reg_1_3 [15] ), .B(_12157_ ), .S(_12011_ ), .Z(_12158_ ) );
AND3_X1 _18969_ ( .A1(_12092_ ), .A2(fanout_net_13 ), .A3(_12158_ ), .ZN(_12159_ ) );
AOI22_X1 _18970_ ( .A1(_12158_ ), .A2(_11946_ ), .B1(_12149_ ), .B2(_12060_ ), .ZN(_12160_ ) );
AOI21_X1 _18971_ ( .A(_12160_ ), .B1(_12109_ ), .B2(fanout_net_13 ), .ZN(_12161_ ) );
OAI21_X1 _18972_ ( .A(_12091_ ), .B1(_12159_ ), .B2(_12161_ ), .ZN(_12162_ ) );
NAND2_X1 _18973_ ( .A1(_12151_ ), .A2(_12162_ ), .ZN(\ifu.io_out_bits_inst [15] ) );
AOI21_X1 _18974_ ( .A(fanout_net_21 ), .B1(_12151_ ), .B2(_12162_ ), .ZN(_00239_ ) );
AND2_X1 _18975_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [14] ), .ZN(_12163_ ) );
AND4_X1 _18976_ ( .A1(_12023_ ), .A2(_11983_ ), .A3(_11984_ ), .A4(_12163_ ), .ZN(_12164_ ) );
AOI21_X1 _18977_ ( .A(_12164_ ), .B1(_11987_ ), .B2(\ifu.inst [14] ), .ZN(_12165_ ) );
NOR4_X1 _18978_ ( .A1(_11933_ ), .A2(\icache.icache_reg_1_1 [14] ), .A3(_11515_ ), .A4(_11995_ ), .ZN(_12166_ ) );
NOR4_X1 _18979_ ( .A1(_11933_ ), .A2(\icache.icache_reg_0_3 [14] ), .A3(_10837_ ), .A4(_11905_ ), .ZN(_12167_ ) );
NOR2_X1 _18980_ ( .A1(_12167_ ), .A2(_11917_ ), .ZN(_12168_ ) );
MUX2_X1 _18981_ ( .A(\icache.icache_reg_0_0 [14] ), .B(\icache.icache_reg_0_1 [14] ), .S(_11912_ ), .Z(_12169_ ) );
MUX2_X1 _18982_ ( .A(\icache.icache_reg_0_2 [14] ), .B(_12169_ ), .S(_12001_ ), .Z(_12170_ ) );
OAI21_X1 _18983_ ( .A(_12168_ ), .B1(_12170_ ), .B2(_12004_ ), .ZN(_12171_ ) );
OAI211_X1 _18984_ ( .A(_11505_ ), .B(_11935_ ), .C1(_11993_ ), .C2(\icache.icache_reg_1_0 [14] ), .ZN(_12172_ ) );
AOI21_X1 _18985_ ( .A(_12166_ ), .B1(_12171_ ), .B2(_12172_ ), .ZN(_12173_ ) );
MUX2_X1 _18986_ ( .A(\icache.icache_reg_1_2 [14] ), .B(_12173_ ), .S(_12056_ ), .Z(_12174_ ) );
MUX2_X1 _18987_ ( .A(\icache.icache_reg_1_3 [14] ), .B(_12174_ ), .S(_12143_ ), .Z(_12175_ ) );
AND4_X1 _18988_ ( .A1(fanout_net_13 ), .A2(_11902_ ), .A3(_12048_ ), .A4(_12175_ ), .ZN(_12176_ ) );
BUF_X4 _18989_ ( .A(_11945_ ), .Z(_12177_ ) );
AOI22_X1 _18990_ ( .A1(_12175_ ), .A2(_12177_ ), .B1(_12163_ ), .B2(_12060_ ), .ZN(_12178_ ) );
AOI21_X1 _18991_ ( .A(_12178_ ), .B1(_12109_ ), .B2(fanout_net_13 ), .ZN(_12179_ ) );
OAI21_X1 _18992_ ( .A(_11990_ ), .B1(_12176_ ), .B2(_12179_ ), .ZN(_12180_ ) );
NAND2_X1 _18993_ ( .A1(_12165_ ), .A2(_12180_ ), .ZN(\ifu.io_out_bits_inst [14] ) );
AOI21_X1 _18994_ ( .A(fanout_net_21 ), .B1(_12165_ ), .B2(_12180_ ), .ZN(_00240_ ) );
AND2_X1 _18995_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [13] ), .ZN(_12181_ ) );
AND4_X1 _18996_ ( .A1(_12023_ ), .A2(_11983_ ), .A3(_11984_ ), .A4(_12181_ ), .ZN(_12182_ ) );
AOI21_X1 _18997_ ( .A(_12182_ ), .B1(_11987_ ), .B2(\ifu.inst [13] ), .ZN(_12183_ ) );
NAND3_X1 _18998_ ( .A1(_11940_ ), .A2(_12181_ ), .A3(_11895_ ), .ZN(_12184_ ) );
NOR4_X1 _18999_ ( .A1(_11993_ ), .A2(\icache.icache_reg_1_2 [13] ), .A3(_10835_ ), .A4(_11935_ ), .ZN(_12185_ ) );
AND3_X1 _19000_ ( .A1(_12074_ ), .A2(\icache.icache_reg_0_2 [13] ), .A3(_10834_ ), .ZN(_12186_ ) );
MUX2_X1 _19001_ ( .A(\icache.icache_reg_0_0 [13] ), .B(\icache.icache_reg_0_1 [13] ), .S(_12071_ ), .Z(_12187_ ) );
AOI211_X1 _19002_ ( .A(_12004_ ), .B(_12186_ ), .C1(_12187_ ), .C2(_12070_ ), .ZN(_12188_ ) );
NOR4_X1 _19003_ ( .A1(_11933_ ), .A2(\icache.icache_reg_0_3 [13] ), .A3(_10838_ ), .A4(_11935_ ), .ZN(_12189_ ) );
NOR3_X1 _19004_ ( .A1(_12188_ ), .A2(_12112_ ), .A3(_12189_ ), .ZN(_12190_ ) );
AND3_X1 _19005_ ( .A1(_11480_ ), .A2(\icache.icache_reg_1_0 [13] ), .A3(_11505_ ), .ZN(_12191_ ) );
OAI21_X1 _19006_ ( .A(_11923_ ), .B1(_12190_ ), .B2(_12191_ ), .ZN(_12192_ ) );
AOI21_X1 _19007_ ( .A(_11925_ ), .B1(_12117_ ), .B2(\icache.icache_reg_1_1 [13] ), .ZN(_12193_ ) );
AOI211_X1 _19008_ ( .A(_11931_ ), .B(_12185_ ), .C1(_12192_ ), .C2(_12193_ ), .ZN(_12194_ ) );
AOI21_X1 _19009_ ( .A(_12194_ ), .B1(\icache.icache_reg_1_3 [13] ), .B2(_11931_ ), .ZN(_12195_ ) );
OR2_X1 _19010_ ( .A1(_12195_ ), .A2(_12014_ ), .ZN(_12196_ ) );
AOI22_X1 _19011_ ( .A1(_11991_ ), .A2(fanout_net_13 ), .B1(_12184_ ), .B2(_12196_ ), .ZN(_12197_ ) );
NOR4_X1 _19012_ ( .A1(_12017_ ), .A2(_12019_ ), .A3(_12020_ ), .A4(_12195_ ), .ZN(_12198_ ) );
OAI21_X1 _19013_ ( .A(_11990_ ), .B1(_12197_ ), .B2(_12198_ ), .ZN(_12199_ ) );
NAND2_X1 _19014_ ( .A1(_12183_ ), .A2(_12199_ ), .ZN(\ifu.io_out_bits_inst [13] ) );
AOI21_X1 _19015_ ( .A(fanout_net_21 ), .B1(_12183_ ), .B2(_12199_ ), .ZN(_00241_ ) );
INV_X1 _19016_ ( .A(_10708_ ), .ZN(_12200_ ) );
INV_X1 _19017_ ( .A(_11949_ ), .ZN(_12201_ ) );
NAND3_X1 _19018_ ( .A1(_12200_ ), .A2(\ifu.inst [12] ), .A3(_12201_ ), .ZN(_12202_ ) );
NAND4_X1 _19019_ ( .A1(_11977_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [12] ), .A4(_11950_ ), .ZN(_12203_ ) );
INV_X1 _19020_ ( .A(_10706_ ), .ZN(_12204_ ) );
AND3_X1 _19021_ ( .A1(_12074_ ), .A2(\icache.icache_reg_1_2 [12] ), .A3(_10839_ ), .ZN(_12205_ ) );
NOR4_X1 _19022_ ( .A1(_11933_ ), .A2(\icache.icache_reg_1_1 [12] ), .A3(_10835_ ), .A4(_11995_ ), .ZN(_12206_ ) );
AOI21_X1 _19023_ ( .A(_11917_ ), .B1(_12004_ ), .B2(_11673_ ), .ZN(_12207_ ) );
MUX2_X1 _19024_ ( .A(\icache.icache_reg_0_0 [12] ), .B(\icache.icache_reg_0_1 [12] ), .S(_12071_ ), .Z(_12208_ ) );
MUX2_X1 _19025_ ( .A(\icache.icache_reg_0_2 [12] ), .B(_12208_ ), .S(_12070_ ), .Z(_12209_ ) );
OAI21_X1 _19026_ ( .A(_12207_ ), .B1(_12209_ ), .B2(_12004_ ), .ZN(_12210_ ) );
OAI211_X1 _19027_ ( .A(_10839_ ), .B(_11935_ ), .C1(_11993_ ), .C2(\icache.icache_reg_1_0 [12] ), .ZN(_12211_ ) );
AOI21_X1 _19028_ ( .A(_12206_ ), .B1(_12210_ ), .B2(_12211_ ), .ZN(_12212_ ) );
AOI211_X1 _19029_ ( .A(_11931_ ), .B(_12205_ ), .C1(_12212_ ), .C2(_11927_ ), .ZN(_12213_ ) );
NOR4_X1 _19030_ ( .A1(_11934_ ), .A2(\icache.icache_reg_1_3 [12] ), .A3(_12037_ ), .A4(_11936_ ), .ZN(_12214_ ) );
NOR4_X1 _19031_ ( .A1(_12204_ ), .A2(_12019_ ), .A3(_12213_ ), .A4(_12214_ ), .ZN(_12215_ ) );
OR3_X1 _19032_ ( .A1(_12213_ ), .A2(_12014_ ), .A3(_12214_ ), .ZN(_12216_ ) );
INV_X1 _19033_ ( .A(_11942_ ), .ZN(_12217_ ) );
OAI21_X1 _19034_ ( .A(_12216_ ), .B1(_11888_ ), .B2(_12217_ ), .ZN(_12218_ ) );
AOI21_X1 _19035_ ( .A(_12215_ ), .B1(_12200_ ), .B2(_12218_ ), .ZN(_12219_ ) );
AND2_X1 _19036_ ( .A1(_11977_ ), .A2(_11950_ ), .ZN(_12220_ ) );
OAI211_X1 _19037_ ( .A(_12202_ ), .B(_12203_ ), .C1(_12219_ ), .C2(_12220_ ), .ZN(\ifu.io_out_bits_inst [12] ) );
AND2_X1 _19038_ ( .A1(\ifu.io_out_bits_inst [12] ), .A2(_10987_ ), .ZN(_00242_ ) );
AND2_X1 _19039_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [29] ), .ZN(_12221_ ) );
AND4_X1 _19040_ ( .A1(_12023_ ), .A2(_11983_ ), .A3(_11984_ ), .A4(_12221_ ), .ZN(_12222_ ) );
AOI21_X1 _19041_ ( .A(_12222_ ), .B1(_11987_ ), .B2(\ifu.inst [29] ), .ZN(_12223_ ) );
NAND3_X1 _19042_ ( .A1(_11480_ ), .A2(\icache.icache_reg_1_0 [29] ), .A3(_10838_ ), .ZN(_12224_ ) );
AND3_X1 _19043_ ( .A1(_11909_ ), .A2(\icache.icache_reg_0_1 [29] ), .A3(_10834_ ), .ZN(_12225_ ) );
AOI211_X1 _19044_ ( .A(_11908_ ), .B(_12225_ ), .C1(_12095_ ), .C2(\icache.icache_reg_0_0 [29] ), .ZN(_12226_ ) );
NOR4_X1 _19045_ ( .A1(_11437_ ), .A2(\icache.icache_reg_0_2 [29] ), .A3(_09818_ ), .A4(_11905_ ), .ZN(_12227_ ) );
OAI21_X1 _19046_ ( .A(_12006_ ), .B1(_12226_ ), .B2(_12227_ ), .ZN(_12228_ ) );
OAI21_X1 _19047_ ( .A(_12228_ ), .B1(\icache.icache_reg_0_3 [29] ), .B2(_12006_ ), .ZN(_12229_ ) );
OAI21_X1 _19048_ ( .A(_12224_ ), .B1(_12229_ ), .B2(_11917_ ), .ZN(_12230_ ) );
MUX2_X1 _19049_ ( .A(\icache.icache_reg_1_1 [29] ), .B(_12230_ ), .S(_12054_ ), .Z(_12231_ ) );
MUX2_X1 _19050_ ( .A(\icache.icache_reg_1_2 [29] ), .B(_12231_ ), .S(_12056_ ), .Z(_12232_ ) );
MUX2_X1 _19051_ ( .A(\icache.icache_reg_1_3 [29] ), .B(_12232_ ), .S(_12143_ ), .Z(_12233_ ) );
AND4_X1 _19052_ ( .A1(fanout_net_13 ), .A2(_11902_ ), .A3(_12048_ ), .A4(_12233_ ), .ZN(_12234_ ) );
AOI22_X1 _19053_ ( .A1(_12233_ ), .A2(_12177_ ), .B1(_12221_ ), .B2(_12060_ ), .ZN(_12235_ ) );
AOI21_X1 _19054_ ( .A(_12235_ ), .B1(_12109_ ), .B2(fanout_net_13 ), .ZN(_12236_ ) );
OAI21_X1 _19055_ ( .A(_11990_ ), .B1(_12234_ ), .B2(_12236_ ), .ZN(_12237_ ) );
NAND2_X1 _19056_ ( .A1(_12223_ ), .A2(_12237_ ), .ZN(\ifu.io_out_bits_inst [29] ) );
AOI21_X1 _19057_ ( .A(fanout_net_21 ), .B1(_12223_ ), .B2(_12237_ ), .ZN(_00243_ ) );
CLKBUF_X2 _19058_ ( .A(_11982_ ), .Z(_12238_ ) );
CLKBUF_X2 _19059_ ( .A(_11976_ ), .Z(_12239_ ) );
AND2_X1 _19060_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [11] ), .ZN(_12240_ ) );
AND4_X1 _19061_ ( .A1(_12023_ ), .A2(_12238_ ), .A3(_12239_ ), .A4(_12240_ ), .ZN(_12241_ ) );
BUF_X4 _19062_ ( .A(_10710_ ), .Z(_12242_ ) );
AOI21_X1 _19063_ ( .A(_12241_ ), .B1(_12242_ ), .B2(\ifu.inst [11] ), .ZN(_12243_ ) );
MUX2_X1 _19064_ ( .A(\icache.icache_reg_0_0 [11] ), .B(\icache.icache_reg_0_1 [11] ), .S(_11911_ ), .Z(_12244_ ) );
MUX2_X1 _19065_ ( .A(\icache.icache_reg_0_2 [11] ), .B(_12244_ ), .S(_12000_ ), .Z(_12245_ ) );
MUX2_X1 _19066_ ( .A(\icache.icache_reg_0_3 [11] ), .B(_12245_ ), .S(_12005_ ), .Z(_12246_ ) );
MUX2_X1 _19067_ ( .A(\icache.icache_reg_1_0 [11] ), .B(_12246_ ), .S(_12052_ ), .Z(_12247_ ) );
MUX2_X1 _19068_ ( .A(\icache.icache_reg_1_1 [11] ), .B(_12247_ ), .S(_12054_ ), .Z(_12248_ ) );
MUX2_X1 _19069_ ( .A(\icache.icache_reg_1_2 [11] ), .B(_12248_ ), .S(_12056_ ), .Z(_12249_ ) );
MUX2_X1 _19070_ ( .A(\icache.icache_reg_1_3 [11] ), .B(_12249_ ), .S(_12143_ ), .Z(_12250_ ) );
AND4_X1 _19071_ ( .A1(fanout_net_13 ), .A2(_11901_ ), .A3(_12048_ ), .A4(_12250_ ), .ZN(_12251_ ) );
AOI22_X1 _19072_ ( .A1(_12250_ ), .A2(_12177_ ), .B1(_12240_ ), .B2(_12060_ ), .ZN(_12252_ ) );
AOI21_X1 _19073_ ( .A(_12252_ ), .B1(_12109_ ), .B2(fanout_net_13 ), .ZN(_12253_ ) );
OAI21_X1 _19074_ ( .A(_11990_ ), .B1(_12251_ ), .B2(_12253_ ), .ZN(_12254_ ) );
NAND2_X1 _19075_ ( .A1(_12243_ ), .A2(_12254_ ), .ZN(\ifu.io_out_bits_inst [11] ) );
AOI21_X1 _19076_ ( .A(fanout_net_21 ), .B1(_12243_ ), .B2(_12254_ ), .ZN(_00244_ ) );
CLKBUF_X2 _19077_ ( .A(_11949_ ), .Z(_12255_ ) );
AND2_X1 _19078_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [10] ), .ZN(_12256_ ) );
AND4_X1 _19079_ ( .A1(_12255_ ), .A2(_12238_ ), .A3(_12239_ ), .A4(_12256_ ), .ZN(_12257_ ) );
AOI21_X1 _19080_ ( .A(_12257_ ), .B1(_12242_ ), .B2(\ifu.inst [10] ), .ZN(_12258_ ) );
OR4_X1 _19081_ ( .A1(\icache.icache_reg_1_3 [10] ), .A2(_11934_ ), .A3(_10836_ ), .A4(_11936_ ), .ZN(_12259_ ) );
NAND3_X1 _19082_ ( .A1(_12074_ ), .A2(\icache.icache_reg_1_2 [10] ), .A3(_11572_ ), .ZN(_12260_ ) );
OR4_X1 _19083_ ( .A1(\icache.icache_reg_0_3 [10] ), .A2(_11933_ ), .A3(_10838_ ), .A4(_11935_ ), .ZN(_12261_ ) );
MUX2_X1 _19084_ ( .A(\icache.icache_reg_0_0 [10] ), .B(\icache.icache_reg_0_1 [10] ), .S(_12071_ ), .Z(_12262_ ) );
MUX2_X1 _19085_ ( .A(\icache.icache_reg_0_2 [10] ), .B(_12262_ ), .S(_12070_ ), .Z(_12263_ ) );
OAI211_X1 _19086_ ( .A(_11919_ ), .B(_12261_ ), .C1(_12263_ ), .C2(_12004_ ), .ZN(_12264_ ) );
NAND4_X1 _19087_ ( .A1(_11934_ ), .A2(\icache.icache_reg_1_0 [10] ), .A3(_10839_ ), .A4(_11936_ ), .ZN(_12265_ ) );
AND3_X1 _19088_ ( .A1(_12264_ ), .A2(_11923_ ), .A3(_12265_ ), .ZN(_12266_ ) );
OAI21_X1 _19089_ ( .A(_12102_ ), .B1(_11923_ ), .B2(\icache.icache_reg_1_1 [10] ), .ZN(_12267_ ) );
OAI211_X1 _19090_ ( .A(_12012_ ), .B(_12260_ ), .C1(_12266_ ), .C2(_12267_ ), .ZN(_12268_ ) );
AND4_X1 _19091_ ( .A1(fanout_net_13 ), .A2(_10706_ ), .A3(_12259_ ), .A4(_12268_ ), .ZN(_12269_ ) );
NAND3_X1 _19092_ ( .A1(_11940_ ), .A2(_12256_ ), .A3(_11895_ ), .ZN(_12270_ ) );
NAND3_X1 _19093_ ( .A1(_12268_ ), .A2(_11945_ ), .A3(_12259_ ), .ZN(_12271_ ) );
AOI22_X1 _19094_ ( .A1(_12092_ ), .A2(fanout_net_13 ), .B1(_12270_ ), .B2(_12271_ ), .ZN(_12272_ ) );
OAI21_X1 _19095_ ( .A(_12091_ ), .B1(_12269_ ), .B2(_12272_ ), .ZN(_12273_ ) );
NAND2_X1 _19096_ ( .A1(_12258_ ), .A2(_12273_ ), .ZN(\ifu.io_out_bits_inst [10] ) );
AOI21_X1 _19097_ ( .A(fanout_net_21 ), .B1(_12258_ ), .B2(_12273_ ), .ZN(_00245_ ) );
AND2_X1 _19098_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [9] ), .ZN(_12274_ ) );
AND4_X1 _19099_ ( .A1(_12255_ ), .A2(_12238_ ), .A3(_12239_ ), .A4(_12274_ ), .ZN(_12275_ ) );
AOI21_X1 _19100_ ( .A(_12275_ ), .B1(_12242_ ), .B2(\ifu.inst [9] ), .ZN(_12276_ ) );
NOR4_X1 _19101_ ( .A1(_12036_ ), .A2(\icache.icache_reg_1_2 [9] ), .A3(_12037_ ), .A4(_11936_ ), .ZN(_12277_ ) );
NOR4_X1 _19102_ ( .A1(_11993_ ), .A2(\icache.icache_reg_1_0 [9] ), .A3(_11515_ ), .A4(_11995_ ), .ZN(_12278_ ) );
NOR2_X1 _19103_ ( .A1(_12278_ ), .A2(_11921_ ), .ZN(_12279_ ) );
MUX2_X1 _19104_ ( .A(\icache.icache_reg_0_0 [9] ), .B(\icache.icache_reg_0_1 [9] ), .S(_11912_ ), .Z(_12280_ ) );
MUX2_X1 _19105_ ( .A(\icache.icache_reg_0_2 [9] ), .B(_12280_ ), .S(_12001_ ), .Z(_12281_ ) );
MUX2_X1 _19106_ ( .A(\icache.icache_reg_0_3 [9] ), .B(_12281_ ), .S(_12073_ ), .Z(_12282_ ) );
OAI21_X1 _19107_ ( .A(_12279_ ), .B1(_12282_ ), .B2(_12112_ ), .ZN(_12283_ ) );
AOI21_X1 _19108_ ( .A(_11925_ ), .B1(_12117_ ), .B2(\icache.icache_reg_1_1 [9] ), .ZN(_12284_ ) );
AOI21_X1 _19109_ ( .A(_12277_ ), .B1(_12283_ ), .B2(_12284_ ), .ZN(_12285_ ) );
MUX2_X1 _19110_ ( .A(\icache.icache_reg_1_3 [9] ), .B(_12285_ ), .S(_12143_ ), .Z(_12286_ ) );
AND4_X1 _19111_ ( .A1(fanout_net_13 ), .A2(_11901_ ), .A3(_11903_ ), .A4(_12286_ ), .ZN(_12287_ ) );
AOI22_X1 _19112_ ( .A1(_12286_ ), .A2(_12177_ ), .B1(_12274_ ), .B2(_12060_ ), .ZN(_12288_ ) );
AOI21_X1 _19113_ ( .A(_12288_ ), .B1(_12109_ ), .B2(fanout_net_13 ), .ZN(_12289_ ) );
OAI21_X1 _19114_ ( .A(_11990_ ), .B1(_12287_ ), .B2(_12289_ ), .ZN(_12290_ ) );
NAND2_X1 _19115_ ( .A1(_12276_ ), .A2(_12290_ ), .ZN(\ifu.io_out_bits_inst [9] ) );
AOI21_X1 _19116_ ( .A(fanout_net_21 ), .B1(_12276_ ), .B2(_12290_ ), .ZN(_00246_ ) );
AND2_X1 _19117_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [8] ), .ZN(_12291_ ) );
AND4_X1 _19118_ ( .A1(_12255_ ), .A2(_12238_ ), .A3(_12239_ ), .A4(_12291_ ), .ZN(_12292_ ) );
AOI21_X1 _19119_ ( .A(_12292_ ), .B1(_12242_ ), .B2(\ifu.inst [8] ), .ZN(_12293_ ) );
MUX2_X1 _19120_ ( .A(\icache.icache_reg_0_0 [8] ), .B(\icache.icache_reg_0_1 [8] ), .S(_11910_ ), .Z(_12294_ ) );
MUX2_X1 _19121_ ( .A(\icache.icache_reg_0_2 [8] ), .B(_12294_ ), .S(_12000_ ), .Z(_12295_ ) );
MUX2_X1 _19122_ ( .A(\icache.icache_reg_0_3 [8] ), .B(_12295_ ), .S(_12005_ ), .Z(_12296_ ) );
MUX2_X1 _19123_ ( .A(\icache.icache_reg_1_0 [8] ), .B(_12296_ ), .S(_12052_ ), .Z(_12297_ ) );
MUX2_X1 _19124_ ( .A(\icache.icache_reg_1_1 [8] ), .B(_12297_ ), .S(_11922_ ), .Z(_12298_ ) );
MUX2_X1 _19125_ ( .A(\icache.icache_reg_1_2 [8] ), .B(_12298_ ), .S(_12056_ ), .Z(_12299_ ) );
MUX2_X1 _19126_ ( .A(\icache.icache_reg_1_3 [8] ), .B(_12299_ ), .S(_12011_ ), .Z(_12300_ ) );
AND3_X1 _19127_ ( .A1(_12092_ ), .A2(fanout_net_13 ), .A3(_12300_ ), .ZN(_12301_ ) );
AOI22_X1 _19128_ ( .A1(_12300_ ), .A2(_12177_ ), .B1(_12291_ ), .B2(_12060_ ), .ZN(_12302_ ) );
AOI21_X1 _19129_ ( .A(_12302_ ), .B1(_12109_ ), .B2(fanout_net_13 ), .ZN(_12303_ ) );
OAI21_X1 _19130_ ( .A(_12091_ ), .B1(_12301_ ), .B2(_12303_ ), .ZN(_12304_ ) );
NAND2_X1 _19131_ ( .A1(_12293_ ), .A2(_12304_ ), .ZN(\ifu.io_out_bits_inst [8] ) );
AOI21_X1 _19132_ ( .A(fanout_net_21 ), .B1(_12293_ ), .B2(_12304_ ), .ZN(_00247_ ) );
AND2_X1 _19133_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [7] ), .ZN(_12305_ ) );
AND4_X1 _19134_ ( .A1(_12255_ ), .A2(_12238_ ), .A3(_12239_ ), .A4(_12305_ ), .ZN(_12306_ ) );
AOI21_X1 _19135_ ( .A(_12306_ ), .B1(_12242_ ), .B2(\ifu.inst [7] ), .ZN(_12307_ ) );
MUX2_X1 _19136_ ( .A(\icache.icache_reg_0_0 [7] ), .B(\icache.icache_reg_0_1 [7] ), .S(_11910_ ), .Z(_12308_ ) );
MUX2_X1 _19137_ ( .A(\icache.icache_reg_0_2 [7] ), .B(_12308_ ), .S(_12000_ ), .Z(_12309_ ) );
MUX2_X1 _19138_ ( .A(\icache.icache_reg_0_3 [7] ), .B(_12309_ ), .S(_12005_ ), .Z(_12310_ ) );
MUX2_X1 _19139_ ( .A(\icache.icache_reg_1_0 [7] ), .B(_12310_ ), .S(_12052_ ), .Z(_12311_ ) );
MUX2_X1 _19140_ ( .A(\icache.icache_reg_1_1 [7] ), .B(_12311_ ), .S(_11922_ ), .Z(_12312_ ) );
MUX2_X1 _19141_ ( .A(\icache.icache_reg_1_2 [7] ), .B(_12312_ ), .S(_11926_ ), .Z(_12313_ ) );
MUX2_X1 _19142_ ( .A(\icache.icache_reg_1_3 [7] ), .B(_12313_ ), .S(_12011_ ), .Z(_12314_ ) );
AND3_X1 _19143_ ( .A1(_12092_ ), .A2(fanout_net_13 ), .A3(_12314_ ), .ZN(_12315_ ) );
AOI22_X1 _19144_ ( .A1(_12314_ ), .A2(_12177_ ), .B1(_12305_ ), .B2(_11942_ ), .ZN(_12316_ ) );
AOI21_X1 _19145_ ( .A(_12316_ ), .B1(_12109_ ), .B2(\icache._io_out_arvalid_T ), .ZN(_12317_ ) );
OAI21_X1 _19146_ ( .A(_12091_ ), .B1(_12315_ ), .B2(_12317_ ), .ZN(_12318_ ) );
NAND2_X1 _19147_ ( .A1(_12307_ ), .A2(_12318_ ), .ZN(\ifu.io_out_bits_inst [7] ) );
AOI21_X1 _19148_ ( .A(fanout_net_21 ), .B1(_12307_ ), .B2(_12318_ ), .ZN(_00248_ ) );
AND4_X1 _19149_ ( .A1(\icache.icache_reg_0_3 [6] ), .A2(_11993_ ), .A3(_10835_ ), .A4(_11995_ ), .ZN(_12319_ ) );
NAND3_X1 _19150_ ( .A1(_12074_ ), .A2(\icache.icache_reg_0_2 [6] ), .A3(_10835_ ), .ZN(_12320_ ) );
AND3_X1 _19151_ ( .A1(_11909_ ), .A2(\icache.icache_reg_0_1 [6] ), .A3(_11515_ ), .ZN(_12321_ ) );
AOI21_X1 _19152_ ( .A(_12321_ ), .B1(_12095_ ), .B2(\icache.icache_reg_0_0 [6] ), .ZN(_12322_ ) );
OAI21_X1 _19153_ ( .A(_12320_ ), .B1(_12322_ ), .B2(_11908_ ), .ZN(_12323_ ) );
AOI211_X1 _19154_ ( .A(_12112_ ), .B(_12319_ ), .C1(_12323_ ), .C2(_12073_ ), .ZN(_12324_ ) );
NOR4_X1 _19155_ ( .A1(_12036_ ), .A2(\icache.icache_reg_1_0 [6] ), .A3(_12037_ ), .A4(_11996_ ), .ZN(_12325_ ) );
NOR3_X1 _19156_ ( .A1(_12324_ ), .A2(_12117_ ), .A3(_12325_ ), .ZN(_12326_ ) );
NAND3_X1 _19157_ ( .A1(_11909_ ), .A2(\icache.icache_reg_1_1 [6] ), .A3(_10840_ ), .ZN(_12327_ ) );
NAND2_X1 _19158_ ( .A1(_12102_ ), .A2(_12327_ ), .ZN(_12328_ ) );
OAI221_X1 _19159_ ( .A(_12012_ ), .B1(\icache.icache_reg_1_2 [6] ), .B2(_12102_ ), .C1(_12326_ ), .C2(_12328_ ), .ZN(_12329_ ) );
NAND4_X1 _19160_ ( .A1(_11994_ ), .A2(\icache.icache_reg_1_3 [6] ), .A3(_11643_ ), .A4(_11997_ ), .ZN(_12330_ ) );
NAND2_X1 _19161_ ( .A1(_12329_ ), .A2(_12330_ ), .ZN(_12331_ ) );
NAND4_X1 _19162_ ( .A1(_11902_ ), .A2(\icache._io_out_arvalid_T ), .A3(_11903_ ), .A4(_12331_ ), .ZN(_12332_ ) );
AND3_X1 _19163_ ( .A1(_11941_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [6] ), .ZN(_12333_ ) );
AOI21_X1 _19164_ ( .A(_12333_ ), .B1(_12331_ ), .B2(_11946_ ), .ZN(_12334_ ) );
OAI21_X1 _19165_ ( .A(_12332_ ), .B1(_10708_ ), .B2(_12334_ ), .ZN(_12335_ ) );
AOI22_X1 _19166_ ( .A1(_12335_ ), .A2(_11951_ ), .B1(_11952_ ), .B2(\ifu.inst [6] ), .ZN(_12336_ ) );
NAND4_X1 _19167_ ( .A1(_11977_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [6] ), .A4(_11950_ ), .ZN(_12337_ ) );
NAND2_X1 _19168_ ( .A1(_12336_ ), .A2(_12337_ ), .ZN(\ifu.io_out_bits_inst [6] ) );
AOI21_X1 _19169_ ( .A(fanout_net_21 ), .B1(_12336_ ), .B2(_12337_ ), .ZN(_00249_ ) );
AND4_X1 _19170_ ( .A1(\icache.icache_reg_0_3 [5] ), .A2(_11437_ ), .A3(_11515_ ), .A4(_11995_ ), .ZN(_12338_ ) );
MUX2_X1 _19171_ ( .A(\icache.icache_reg_0_0 [5] ), .B(\icache.icache_reg_0_1 [5] ), .S(_12071_ ), .Z(_12339_ ) );
MUX2_X1 _19172_ ( .A(\icache.icache_reg_0_2 [5] ), .B(_12339_ ), .S(_12070_ ), .Z(_12340_ ) );
AOI211_X1 _19173_ ( .A(_12112_ ), .B(_12338_ ), .C1(_12340_ ), .C2(_12073_ ), .ZN(_12341_ ) );
NOR4_X1 _19174_ ( .A1(_12036_ ), .A2(\icache.icache_reg_1_0 [5] ), .A3(_12037_ ), .A4(_11996_ ), .ZN(_12342_ ) );
NOR3_X1 _19175_ ( .A1(_12341_ ), .A2(_12117_ ), .A3(_12342_ ), .ZN(_12343_ ) );
NAND3_X1 _19176_ ( .A1(_11909_ ), .A2(\icache.icache_reg_1_1 [5] ), .A3(_11571_ ), .ZN(_12344_ ) );
NAND2_X1 _19177_ ( .A1(_12102_ ), .A2(_12344_ ), .ZN(_12345_ ) );
OAI221_X1 _19178_ ( .A(_12012_ ), .B1(\icache.icache_reg_1_2 [5] ), .B2(_12102_ ), .C1(_12343_ ), .C2(_12345_ ), .ZN(_12346_ ) );
NAND4_X1 _19179_ ( .A1(_11994_ ), .A2(\icache.icache_reg_1_3 [5] ), .A3(_11572_ ), .A4(_11997_ ), .ZN(_12347_ ) );
NAND2_X1 _19180_ ( .A1(_12346_ ), .A2(_12347_ ), .ZN(_12348_ ) );
NAND4_X1 _19181_ ( .A1(_11902_ ), .A2(\icache._io_out_arvalid_T ), .A3(_10704_ ), .A4(_12348_ ), .ZN(_12349_ ) );
AND3_X1 _19182_ ( .A1(_11941_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [5] ), .ZN(_12350_ ) );
AOI21_X1 _19183_ ( .A(_12350_ ), .B1(_12348_ ), .B2(_11946_ ), .ZN(_12351_ ) );
OAI21_X1 _19184_ ( .A(_12349_ ), .B1(_10708_ ), .B2(_12351_ ), .ZN(_12352_ ) );
AOI22_X1 _19185_ ( .A1(_12352_ ), .A2(_11951_ ), .B1(_11952_ ), .B2(\ifu.inst [5] ), .ZN(_12353_ ) );
NAND4_X1 _19186_ ( .A1(_11977_ ), .A2(fanout_net_3 ), .A3(\io_master_rdata [5] ), .A4(_11950_ ), .ZN(_12354_ ) );
NAND2_X1 _19187_ ( .A1(_12353_ ), .A2(_12354_ ), .ZN(\ifu.io_out_bits_inst [5] ) );
AOI21_X1 _19188_ ( .A(fanout_net_21 ), .B1(_12353_ ), .B2(_12354_ ), .ZN(_00250_ ) );
AND2_X1 _19189_ ( .A1(fanout_net_3 ), .A2(\io_master_rdata [4] ), .ZN(_12355_ ) );
AND4_X1 _19190_ ( .A1(_12255_ ), .A2(_12238_ ), .A3(_12239_ ), .A4(_12355_ ), .ZN(_12356_ ) );
AOI21_X1 _19191_ ( .A(_12356_ ), .B1(_12242_ ), .B2(\ifu.inst [4] ), .ZN(_12357_ ) );
BUF_X4 _19192_ ( .A(_11989_ ), .Z(_12358_ ) );
NOR4_X1 _19193_ ( .A1(_11934_ ), .A2(\icache.icache_reg_1_3 [4] ), .A3(_10836_ ), .A4(_11936_ ), .ZN(_12359_ ) );
AOI21_X1 _19194_ ( .A(_11925_ ), .B1(_12117_ ), .B2(_11773_ ), .ZN(_12360_ ) );
MUX2_X1 _19195_ ( .A(\icache.icache_reg_0_0 [4] ), .B(\icache.icache_reg_0_1 [4] ), .S(_11912_ ), .Z(_12361_ ) );
MUX2_X1 _19196_ ( .A(\icache.icache_reg_0_2 [4] ), .B(_12361_ ), .S(_12001_ ), .Z(_12362_ ) );
MUX2_X1 _19197_ ( .A(\icache.icache_reg_0_3 [4] ), .B(_12362_ ), .S(_12006_ ), .Z(_12363_ ) );
MUX2_X1 _19198_ ( .A(\icache.icache_reg_1_0 [4] ), .B(_12363_ ), .S(_11919_ ), .Z(_12364_ ) );
OAI21_X1 _19199_ ( .A(_12360_ ), .B1(_12364_ ), .B2(_12117_ ), .ZN(_12365_ ) );
OAI211_X1 _19200_ ( .A(_11572_ ), .B(_11997_ ), .C1(_11994_ ), .C2(\icache.icache_reg_1_2 [4] ), .ZN(_12366_ ) );
AOI21_X1 _19201_ ( .A(_12359_ ), .B1(_12365_ ), .B2(_12366_ ), .ZN(_12367_ ) );
AND4_X1 _19202_ ( .A1(\icache._io_out_arvalid_T ), .A2(_11901_ ), .A3(_11903_ ), .A4(_12367_ ), .ZN(_12368_ ) );
AOI22_X1 _19203_ ( .A1(_12367_ ), .A2(_12177_ ), .B1(_12355_ ), .B2(_11942_ ), .ZN(_12369_ ) );
AOI21_X1 _19204_ ( .A(_12369_ ), .B1(_12109_ ), .B2(\icache._io_out_arvalid_T ), .ZN(_12370_ ) );
OAI21_X1 _19205_ ( .A(_12358_ ), .B1(_12368_ ), .B2(_12370_ ), .ZN(_12371_ ) );
NAND2_X1 _19206_ ( .A1(_12357_ ), .A2(_12371_ ), .ZN(\ifu.io_out_bits_inst [4] ) );
AOI21_X1 _19207_ ( .A(fanout_net_21 ), .B1(_12357_ ), .B2(_12371_ ), .ZN(_00251_ ) );
AND4_X1 _19208_ ( .A1(\icache.icache_reg_0_3 [3] ), .A2(_11437_ ), .A3(_11515_ ), .A4(_11995_ ), .ZN(_12372_ ) );
MUX2_X1 _19209_ ( .A(\icache.icache_reg_0_0 [3] ), .B(\icache.icache_reg_0_1 [3] ), .S(_12071_ ), .Z(_12373_ ) );
MUX2_X1 _19210_ ( .A(\icache.icache_reg_0_2 [3] ), .B(_12373_ ), .S(_12070_ ), .Z(_12374_ ) );
AOI211_X1 _19211_ ( .A(_12112_ ), .B(_12372_ ), .C1(_12374_ ), .C2(_12073_ ), .ZN(_12375_ ) );
NOR4_X1 _19212_ ( .A1(_12036_ ), .A2(\icache.icache_reg_1_0 [3] ), .A3(_12037_ ), .A4(_11996_ ), .ZN(_12376_ ) );
NOR3_X1 _19213_ ( .A1(_12375_ ), .A2(_12117_ ), .A3(_12376_ ), .ZN(_12377_ ) );
NAND3_X1 _19214_ ( .A1(_11909_ ), .A2(\icache.icache_reg_1_1 [3] ), .A3(_11571_ ), .ZN(_12378_ ) );
NAND2_X1 _19215_ ( .A1(_12102_ ), .A2(_12378_ ), .ZN(_12379_ ) );
OAI221_X1 _19216_ ( .A(_12012_ ), .B1(\icache.icache_reg_1_2 [3] ), .B2(_12102_ ), .C1(_12377_ ), .C2(_12379_ ), .ZN(_12380_ ) );
NAND4_X1 _19217_ ( .A1(_11994_ ), .A2(\icache.icache_reg_1_3 [3] ), .A3(_11572_ ), .A4(_11997_ ), .ZN(_12381_ ) );
NAND2_X1 _19218_ ( .A1(_12380_ ), .A2(_12381_ ), .ZN(_12382_ ) );
NAND4_X1 _19219_ ( .A1(_11902_ ), .A2(\icache._io_out_arvalid_T ), .A3(_10704_ ), .A4(_12382_ ), .ZN(_12383_ ) );
AND3_X1 _19220_ ( .A1(_11941_ ), .A2(\arbiter._io_axi_araddr_T_6 ), .A3(\io_master_rdata [3] ), .ZN(_12384_ ) );
AOI21_X1 _19221_ ( .A(_12384_ ), .B1(_12382_ ), .B2(_11946_ ), .ZN(_12385_ ) );
OAI21_X1 _19222_ ( .A(_12383_ ), .B1(_10708_ ), .B2(_12385_ ), .ZN(_12386_ ) );
AOI22_X1 _19223_ ( .A1(_12386_ ), .A2(_11951_ ), .B1(_10710_ ), .B2(\ifu.inst [3] ), .ZN(_12387_ ) );
NAND4_X1 _19224_ ( .A1(_11977_ ), .A2(\arbiter._io_axi_araddr_T_6 ), .A3(\io_master_rdata [3] ), .A4(_11950_ ), .ZN(_12388_ ) );
NAND2_X1 _19225_ ( .A1(_12387_ ), .A2(_12388_ ), .ZN(\ifu.io_out_bits_inst [3] ) );
AOI21_X1 _19226_ ( .A(fanout_net_21 ), .B1(_12387_ ), .B2(_12388_ ), .ZN(_00252_ ) );
AND2_X1 _19227_ ( .A1(\arbiter._io_axi_araddr_T_6 ), .A2(\io_master_rdata [2] ), .ZN(_12389_ ) );
AND4_X1 _19228_ ( .A1(_12255_ ), .A2(_12238_ ), .A3(_12239_ ), .A4(_12389_ ), .ZN(_12390_ ) );
AOI21_X1 _19229_ ( .A(_12390_ ), .B1(_12242_ ), .B2(\ifu.inst [2] ), .ZN(_12391_ ) );
NAND3_X1 _19230_ ( .A1(_11940_ ), .A2(_12389_ ), .A3(_11895_ ), .ZN(_12392_ ) );
NAND4_X1 _19231_ ( .A1(_11933_ ), .A2(\icache.icache_reg_1_0 [2] ), .A3(_10838_ ), .A4(_11935_ ), .ZN(_12393_ ) );
OR4_X1 _19232_ ( .A1(\icache.icache_reg_0_1 [2] ), .A2(_11904_ ), .A3(_09818_ ), .A4(_11479_ ), .ZN(_12394_ ) );
OAI211_X1 _19233_ ( .A(_12394_ ), .B(_12001_ ), .C1(\icache.icache_reg_0_0 [2] ), .C2(_12071_ ), .ZN(_12395_ ) );
NAND3_X1 _19234_ ( .A1(_12074_ ), .A2(\icache.icache_reg_0_2 [2] ), .A3(_10834_ ), .ZN(_12396_ ) );
AOI21_X1 _19235_ ( .A(_12004_ ), .B1(_12395_ ), .B2(_12396_ ), .ZN(_12397_ ) );
AOI21_X1 _19236_ ( .A(_12397_ ), .B1(\icache.icache_reg_0_3 [2] ), .B2(_12004_ ), .ZN(_12398_ ) );
OAI211_X1 _19237_ ( .A(_11923_ ), .B(_12393_ ), .C1(_12398_ ), .C2(_12112_ ), .ZN(_12399_ ) );
OAI211_X1 _19238_ ( .A(_12399_ ), .B(_11927_ ), .C1(\icache.icache_reg_1_1 [2] ), .C2(_11923_ ), .ZN(_12400_ ) );
NAND3_X1 _19239_ ( .A1(_12074_ ), .A2(\icache.icache_reg_1_2 [2] ), .A3(_11571_ ), .ZN(_12401_ ) );
AOI21_X1 _19240_ ( .A(_11931_ ), .B1(_12400_ ), .B2(_12401_ ), .ZN(_12402_ ) );
AOI21_X1 _19241_ ( .A(_12402_ ), .B1(\icache.icache_reg_1_3 [2] ), .B2(_11931_ ), .ZN(_12403_ ) );
OR2_X1 _19242_ ( .A1(_12403_ ), .A2(_12014_ ), .ZN(_12404_ ) );
AOI22_X1 _19243_ ( .A1(_11991_ ), .A2(\icache._io_out_arvalid_T ), .B1(_12392_ ), .B2(_12404_ ), .ZN(_12405_ ) );
NOR4_X1 _19244_ ( .A1(_12017_ ), .A2(_12019_ ), .A3(_12020_ ), .A4(_12403_ ), .ZN(_12406_ ) );
OAI21_X1 _19245_ ( .A(_12358_ ), .B1(_12405_ ), .B2(_12406_ ), .ZN(_12407_ ) );
NAND2_X1 _19246_ ( .A1(_12391_ ), .A2(_12407_ ), .ZN(\ifu.io_out_bits_inst [2] ) );
AOI21_X1 _19247_ ( .A(fanout_net_21 ), .B1(_12391_ ), .B2(_12407_ ), .ZN(_00253_ ) );
AND2_X1 _19248_ ( .A1(\arbiter._io_axi_araddr_T_6 ), .A2(\io_master_rdata [28] ), .ZN(_12408_ ) );
AND4_X1 _19249_ ( .A1(_12255_ ), .A2(_12238_ ), .A3(_12239_ ), .A4(_12408_ ), .ZN(_12409_ ) );
AOI21_X1 _19250_ ( .A(_12409_ ), .B1(_12242_ ), .B2(\ifu.inst [28] ), .ZN(_12410_ ) );
NAND3_X1 _19251_ ( .A1(_12074_ ), .A2(\icache.icache_reg_1_2 [28] ), .A3(_11571_ ), .ZN(_12411_ ) );
AND3_X1 _19252_ ( .A1(_11907_ ), .A2(\icache.icache_reg_0_2 [28] ), .A3(_10834_ ), .ZN(_12412_ ) );
MUX2_X1 _19253_ ( .A(\icache.icache_reg_0_0 [28] ), .B(\icache.icache_reg_0_1 [28] ), .S(_12071_ ), .Z(_12413_ ) );
AOI211_X1 _19254_ ( .A(_12004_ ), .B(_12412_ ), .C1(_12413_ ), .C2(_12070_ ), .ZN(_12414_ ) );
NOR4_X1 _19255_ ( .A1(_11933_ ), .A2(\icache.icache_reg_0_3 [28] ), .A3(_10838_ ), .A4(_11935_ ), .ZN(_12415_ ) );
NOR3_X1 _19256_ ( .A1(_12414_ ), .A2(_11917_ ), .A3(_12415_ ), .ZN(_12416_ ) );
AOI211_X1 _19257_ ( .A(_11921_ ), .B(_12416_ ), .C1(\icache.icache_reg_1_0 [28] ), .C2(_12112_ ), .ZN(_12417_ ) );
OAI21_X1 _19258_ ( .A(_11927_ ), .B1(_11923_ ), .B2(\icache.icache_reg_1_1 [28] ), .ZN(_12418_ ) );
OAI21_X1 _19259_ ( .A(_12411_ ), .B1(_12417_ ), .B2(_12418_ ), .ZN(_12419_ ) );
MUX2_X1 _19260_ ( .A(\icache.icache_reg_1_3 [28] ), .B(_12419_ ), .S(_12143_ ), .Z(_12420_ ) );
AND4_X1 _19261_ ( .A1(\icache._io_out_arvalid_T ), .A2(_11901_ ), .A3(_11903_ ), .A4(_12420_ ), .ZN(_12421_ ) );
AOI22_X1 _19262_ ( .A1(_12420_ ), .A2(_12177_ ), .B1(_12408_ ), .B2(_11942_ ), .ZN(_12422_ ) );
AOI21_X1 _19263_ ( .A(_12422_ ), .B1(_12092_ ), .B2(\icache._io_out_arvalid_T ), .ZN(_12423_ ) );
OAI21_X1 _19264_ ( .A(_12358_ ), .B1(_12421_ ), .B2(_12423_ ), .ZN(_12424_ ) );
NAND2_X1 _19265_ ( .A1(_12410_ ), .A2(_12424_ ), .ZN(\ifu.io_out_bits_inst [28] ) );
AOI21_X1 _19266_ ( .A(fanout_net_21 ), .B1(_12410_ ), .B2(_12424_ ), .ZN(_00254_ ) );
AND2_X1 _19267_ ( .A1(\arbiter._io_axi_araddr_T_6 ), .A2(\io_master_rdata [1] ), .ZN(_12425_ ) );
AND4_X1 _19268_ ( .A1(_12255_ ), .A2(_12238_ ), .A3(_12239_ ), .A4(_12425_ ), .ZN(_12426_ ) );
AOI21_X1 _19269_ ( .A(_12426_ ), .B1(_12242_ ), .B2(\ifu.inst [1] ), .ZN(_12427_ ) );
NAND3_X1 _19270_ ( .A1(_11940_ ), .A2(_12425_ ), .A3(_11895_ ), .ZN(_12428_ ) );
AND4_X1 _19271_ ( .A1(\icache.icache_reg_1_3 [1] ), .A2(_12036_ ), .A3(_11571_ ), .A4(_11996_ ), .ZN(_12429_ ) );
NAND4_X1 _19272_ ( .A1(_11993_ ), .A2(\icache.icache_reg_1_1 [1] ), .A3(_11505_ ), .A4(_11935_ ), .ZN(_12430_ ) );
NOR4_X1 _19273_ ( .A1(_11904_ ), .A2(\icache.icache_reg_0_3 [1] ), .A3(_10837_ ), .A4(_11905_ ), .ZN(_12431_ ) );
AND3_X1 _19274_ ( .A1(_11907_ ), .A2(\icache.icache_reg_0_2 [1] ), .A3(_10834_ ), .ZN(_12432_ ) );
MUX2_X1 _19275_ ( .A(\icache.icache_reg_0_0 [1] ), .B(\icache.icache_reg_0_1 [1] ), .S(_11912_ ), .Z(_12433_ ) );
AOI21_X1 _19276_ ( .A(_12432_ ), .B1(_12433_ ), .B2(_12070_ ), .ZN(_12434_ ) );
AOI211_X1 _19277_ ( .A(_11917_ ), .B(_12431_ ), .C1(_12434_ ), .C2(_12006_ ), .ZN(_12435_ ) );
AOI21_X1 _19278_ ( .A(_12435_ ), .B1(\icache.icache_reg_1_0 [1] ), .B2(_12112_ ), .ZN(_12436_ ) );
OAI21_X1 _19279_ ( .A(_12430_ ), .B1(_12436_ ), .B2(_11921_ ), .ZN(_12437_ ) );
MUX2_X1 _19280_ ( .A(\icache.icache_reg_1_2 [1] ), .B(_12437_ ), .S(_11927_ ), .Z(_12438_ ) );
AOI21_X1 _19281_ ( .A(_12429_ ), .B1(_12438_ ), .B2(_12012_ ), .ZN(_12439_ ) );
OR2_X1 _19282_ ( .A1(_12439_ ), .A2(_12014_ ), .ZN(_12440_ ) );
AOI22_X1 _19283_ ( .A1(_11991_ ), .A2(\icache._io_out_arvalid_T ), .B1(_12428_ ), .B2(_12440_ ), .ZN(_12441_ ) );
NOR4_X1 _19284_ ( .A1(_12017_ ), .A2(_12019_ ), .A3(_12020_ ), .A4(_12439_ ), .ZN(_12442_ ) );
OAI21_X1 _19285_ ( .A(_12358_ ), .B1(_12441_ ), .B2(_12442_ ), .ZN(_12443_ ) );
NAND2_X1 _19286_ ( .A1(_12427_ ), .A2(_12443_ ), .ZN(\ifu.io_out_bits_inst [1] ) );
AOI21_X1 _19287_ ( .A(fanout_net_21 ), .B1(_12427_ ), .B2(_12443_ ), .ZN(_00255_ ) );
AND2_X1 _19288_ ( .A1(\arbiter._io_axi_araddr_T_6 ), .A2(\io_master_rdata [0] ), .ZN(_12444_ ) );
AND4_X1 _19289_ ( .A1(_12255_ ), .A2(_12238_ ), .A3(_12239_ ), .A4(_12444_ ), .ZN(_12445_ ) );
AOI21_X1 _19290_ ( .A(_12445_ ), .B1(_12242_ ), .B2(\ifu.inst [0] ), .ZN(_12446_ ) );
NAND3_X1 _19291_ ( .A1(_11940_ ), .A2(_12444_ ), .A3(_11895_ ), .ZN(_12447_ ) );
OR4_X1 _19292_ ( .A1(\icache.icache_reg_1_1 [0] ), .A2(_11933_ ), .A3(_11515_ ), .A4(_11995_ ), .ZN(_12448_ ) );
MUX2_X1 _19293_ ( .A(\icache.icache_reg_0_0 [0] ), .B(\icache.icache_reg_0_1 [0] ), .S(_11911_ ), .Z(_12449_ ) );
MUX2_X1 _19294_ ( .A(\icache.icache_reg_0_2 [0] ), .B(_12449_ ), .S(_12001_ ), .Z(_12450_ ) );
MUX2_X1 _19295_ ( .A(\icache.icache_reg_0_3 [0] ), .B(_12450_ ), .S(_12006_ ), .Z(_12451_ ) );
MUX2_X1 _19296_ ( .A(\icache.icache_reg_1_0 [0] ), .B(_12451_ ), .S(_11919_ ), .Z(_12452_ ) );
OAI211_X1 _19297_ ( .A(_11927_ ), .B(_12448_ ), .C1(_12452_ ), .C2(_12117_ ), .ZN(_12453_ ) );
NAND3_X1 _19298_ ( .A1(_12074_ ), .A2(\icache.icache_reg_1_2 [0] ), .A3(_11571_ ), .ZN(_12454_ ) );
AOI21_X1 _19299_ ( .A(_11931_ ), .B1(_12453_ ), .B2(_12454_ ), .ZN(_12455_ ) );
AOI21_X1 _19300_ ( .A(_12455_ ), .B1(\icache.icache_reg_1_3 [0] ), .B2(_11931_ ), .ZN(_12456_ ) );
OR2_X1 _19301_ ( .A1(_12456_ ), .A2(_12014_ ), .ZN(_12457_ ) );
AOI22_X1 _19302_ ( .A1(_11991_ ), .A2(\icache._io_out_arvalid_T ), .B1(_12447_ ), .B2(_12457_ ), .ZN(_12458_ ) );
NOR4_X1 _19303_ ( .A1(_12017_ ), .A2(_12019_ ), .A3(_12020_ ), .A4(_12456_ ), .ZN(_12459_ ) );
OAI21_X1 _19304_ ( .A(_12358_ ), .B1(_12458_ ), .B2(_12459_ ), .ZN(_12460_ ) );
NAND2_X1 _19305_ ( .A1(_12446_ ), .A2(_12460_ ), .ZN(\ifu.io_out_bits_inst [0] ) );
AOI21_X1 _19306_ ( .A(fanout_net_21 ), .B1(_12446_ ), .B2(_12460_ ), .ZN(_00256_ ) );
AND2_X1 _19307_ ( .A1(\arbiter._io_axi_araddr_T_6 ), .A2(\io_master_rdata [27] ), .ZN(_12461_ ) );
AND4_X1 _19308_ ( .A1(_12255_ ), .A2(_11982_ ), .A3(_11976_ ), .A4(_12461_ ), .ZN(_12462_ ) );
AOI21_X1 _19309_ ( .A(_12462_ ), .B1(_11952_ ), .B2(\ifu.inst [27] ), .ZN(_12463_ ) );
MUX2_X1 _19310_ ( .A(\icache.icache_reg_0_0 [27] ), .B(\icache.icache_reg_0_1 [27] ), .S(_11911_ ), .Z(_12464_ ) );
MUX2_X1 _19311_ ( .A(\icache.icache_reg_0_2 [27] ), .B(_12464_ ), .S(_12000_ ), .Z(_12465_ ) );
MUX2_X1 _19312_ ( .A(\icache.icache_reg_0_3 [27] ), .B(_12465_ ), .S(_12005_ ), .Z(_12466_ ) );
MUX2_X1 _19313_ ( .A(\icache.icache_reg_1_0 [27] ), .B(_12466_ ), .S(_12052_ ), .Z(_12467_ ) );
MUX2_X1 _19314_ ( .A(\icache.icache_reg_1_1 [27] ), .B(_12467_ ), .S(_12054_ ), .Z(_12468_ ) );
MUX2_X1 _19315_ ( .A(\icache.icache_reg_1_2 [27] ), .B(_12468_ ), .S(_12056_ ), .Z(_12469_ ) );
MUX2_X1 _19316_ ( .A(\icache.icache_reg_1_3 [27] ), .B(_12469_ ), .S(_12143_ ), .Z(_12470_ ) );
AND4_X1 _19317_ ( .A1(\icache._io_out_arvalid_T ), .A2(_11901_ ), .A3(_11903_ ), .A4(_12470_ ), .ZN(_12471_ ) );
AOI22_X1 _19318_ ( .A1(_12470_ ), .A2(_12177_ ), .B1(_12461_ ), .B2(_11942_ ), .ZN(_12472_ ) );
AOI21_X1 _19319_ ( .A(_12472_ ), .B1(_12092_ ), .B2(\icache._io_out_arvalid_T ), .ZN(_12473_ ) );
OAI21_X1 _19320_ ( .A(_12358_ ), .B1(_12471_ ), .B2(_12473_ ), .ZN(_12474_ ) );
NAND2_X1 _19321_ ( .A1(_12463_ ), .A2(_12474_ ), .ZN(\ifu.io_out_bits_inst [27] ) );
AOI21_X1 _19322_ ( .A(fanout_net_21 ), .B1(_12463_ ), .B2(_12474_ ), .ZN(_00257_ ) );
AND2_X1 _19323_ ( .A1(\arbiter._io_axi_araddr_T_6 ), .A2(\io_master_rdata [26] ), .ZN(_12475_ ) );
AND4_X1 _19324_ ( .A1(_11949_ ), .A2(_11982_ ), .A3(_11976_ ), .A4(_12475_ ), .ZN(_12476_ ) );
AOI21_X1 _19325_ ( .A(_12476_ ), .B1(_11952_ ), .B2(\ifu.inst [26] ), .ZN(_12477_ ) );
MUX2_X1 _19326_ ( .A(\icache.icache_reg_0_0 [26] ), .B(\icache.icache_reg_0_1 [26] ), .S(_11911_ ), .Z(_12478_ ) );
MUX2_X1 _19327_ ( .A(\icache.icache_reg_0_2 [26] ), .B(_12478_ ), .S(_12000_ ), .Z(_12479_ ) );
MUX2_X1 _19328_ ( .A(\icache.icache_reg_0_3 [26] ), .B(_12479_ ), .S(_12005_ ), .Z(_12480_ ) );
MUX2_X1 _19329_ ( .A(\icache.icache_reg_1_0 [26] ), .B(_12480_ ), .S(_12052_ ), .Z(_12481_ ) );
MUX2_X1 _19330_ ( .A(\icache.icache_reg_1_1 [26] ), .B(_12481_ ), .S(_12054_ ), .Z(_12482_ ) );
MUX2_X1 _19331_ ( .A(\icache.icache_reg_1_2 [26] ), .B(_12482_ ), .S(_12056_ ), .Z(_12483_ ) );
MUX2_X1 _19332_ ( .A(\icache.icache_reg_1_3 [26] ), .B(_12483_ ), .S(_12143_ ), .Z(_12484_ ) );
AND4_X1 _19333_ ( .A1(\icache._io_out_arvalid_T ), .A2(_11901_ ), .A3(_11903_ ), .A4(_12484_ ), .ZN(_12485_ ) );
AOI22_X1 _19334_ ( .A1(_12484_ ), .A2(_12177_ ), .B1(_12475_ ), .B2(_11942_ ), .ZN(_12486_ ) );
AOI21_X1 _19335_ ( .A(_12486_ ), .B1(_12092_ ), .B2(\icache._io_out_arvalid_T ), .ZN(_12487_ ) );
OAI21_X1 _19336_ ( .A(_12358_ ), .B1(_12485_ ), .B2(_12487_ ), .ZN(_12488_ ) );
NAND2_X1 _19337_ ( .A1(_12477_ ), .A2(_12488_ ), .ZN(\ifu.io_out_bits_inst [26] ) );
AOI21_X1 _19338_ ( .A(fanout_net_22 ), .B1(_12477_ ), .B2(_12488_ ), .ZN(_00258_ ) );
AND2_X1 _19339_ ( .A1(\arbiter._io_axi_araddr_T_6 ), .A2(\io_master_rdata [25] ), .ZN(_12489_ ) );
AND4_X1 _19340_ ( .A1(_11949_ ), .A2(_11982_ ), .A3(_11976_ ), .A4(_12489_ ), .ZN(_12490_ ) );
AOI21_X1 _19341_ ( .A(_12490_ ), .B1(_11952_ ), .B2(\ifu.inst [25] ), .ZN(_12491_ ) );
NAND3_X1 _19342_ ( .A1(_11940_ ), .A2(_12489_ ), .A3(_11895_ ), .ZN(_12492_ ) );
AND4_X1 _19343_ ( .A1(\icache.icache_reg_1_3 [25] ), .A2(_12036_ ), .A3(_10839_ ), .A4(_11996_ ), .ZN(_12493_ ) );
MUX2_X1 _19344_ ( .A(\icache.icache_reg_0_0 [25] ), .B(\icache.icache_reg_0_1 [25] ), .S(_11911_ ), .Z(_12494_ ) );
MUX2_X1 _19345_ ( .A(\icache.icache_reg_0_2 [25] ), .B(_12494_ ), .S(_12001_ ), .Z(_12495_ ) );
MUX2_X1 _19346_ ( .A(\icache.icache_reg_0_3 [25] ), .B(_12495_ ), .S(_12006_ ), .Z(_12496_ ) );
MUX2_X1 _19347_ ( .A(\icache.icache_reg_1_0 [25] ), .B(_12496_ ), .S(_11919_ ), .Z(_12497_ ) );
MUX2_X1 _19348_ ( .A(\icache.icache_reg_1_1 [25] ), .B(_12497_ ), .S(_12054_ ), .Z(_12498_ ) );
MUX2_X1 _19349_ ( .A(\icache.icache_reg_1_2 [25] ), .B(_12498_ ), .S(_11927_ ), .Z(_12499_ ) );
AOI21_X1 _19350_ ( .A(_12493_ ), .B1(_12499_ ), .B2(_12012_ ), .ZN(_12500_ ) );
OR2_X1 _19351_ ( .A1(_12500_ ), .A2(_12014_ ), .ZN(_12501_ ) );
AOI22_X1 _19352_ ( .A1(_11991_ ), .A2(\icache._io_out_arvalid_T ), .B1(_12492_ ), .B2(_12501_ ), .ZN(_12502_ ) );
NOR4_X1 _19353_ ( .A1(_12017_ ), .A2(_12019_ ), .A3(_12020_ ), .A4(_12500_ ), .ZN(_12503_ ) );
OAI21_X1 _19354_ ( .A(_12358_ ), .B1(_12502_ ), .B2(_12503_ ), .ZN(_12504_ ) );
NAND2_X1 _19355_ ( .A1(_12491_ ), .A2(_12504_ ), .ZN(\ifu.io_out_bits_inst [25] ) );
AOI21_X1 _19356_ ( .A(fanout_net_22 ), .B1(_12491_ ), .B2(_12504_ ), .ZN(_00259_ ) );
AND2_X1 _19357_ ( .A1(\arbiter._io_axi_araddr_T_6 ), .A2(\io_master_rdata [24] ), .ZN(_12505_ ) );
AND4_X1 _19358_ ( .A1(_11949_ ), .A2(_11982_ ), .A3(_11976_ ), .A4(_12505_ ), .ZN(_12506_ ) );
AOI21_X1 _19359_ ( .A(_12506_ ), .B1(_11952_ ), .B2(\ifu.inst [24] ), .ZN(_12507_ ) );
MUX2_X1 _19360_ ( .A(\icache.icache_reg_0_0 [24] ), .B(\icache.icache_reg_0_1 [24] ), .S(_11911_ ), .Z(_12508_ ) );
MUX2_X1 _19361_ ( .A(\icache.icache_reg_0_2 [24] ), .B(_12508_ ), .S(_12000_ ), .Z(_12509_ ) );
MUX2_X1 _19362_ ( .A(\icache.icache_reg_0_3 [24] ), .B(_12509_ ), .S(_12005_ ), .Z(_12510_ ) );
MUX2_X1 _19363_ ( .A(\icache.icache_reg_1_0 [24] ), .B(_12510_ ), .S(_12052_ ), .Z(_12511_ ) );
MUX2_X1 _19364_ ( .A(\icache.icache_reg_1_1 [24] ), .B(_12511_ ), .S(_12054_ ), .Z(_12512_ ) );
MUX2_X1 _19365_ ( .A(\icache.icache_reg_1_2 [24] ), .B(_12512_ ), .S(_12056_ ), .Z(_12513_ ) );
MUX2_X1 _19366_ ( .A(\icache.icache_reg_1_3 [24] ), .B(_12513_ ), .S(_12143_ ), .Z(_12514_ ) );
AND4_X1 _19367_ ( .A1(\icache._io_out_arvalid_T ), .A2(_11901_ ), .A3(_11903_ ), .A4(_12514_ ), .ZN(_12515_ ) );
AOI22_X1 _19368_ ( .A1(_12514_ ), .A2(_11945_ ), .B1(_12505_ ), .B2(_11942_ ), .ZN(_12516_ ) );
AOI21_X1 _19369_ ( .A(_12516_ ), .B1(_12092_ ), .B2(\icache._io_out_arvalid_T ), .ZN(_12517_ ) );
OAI21_X1 _19370_ ( .A(_12358_ ), .B1(_12515_ ), .B2(_12517_ ), .ZN(_12518_ ) );
NAND2_X1 _19371_ ( .A1(_12507_ ), .A2(_12518_ ), .ZN(\ifu.io_out_bits_inst [24] ) );
AOI21_X1 _19372_ ( .A(fanout_net_22 ), .B1(_12507_ ), .B2(_12518_ ), .ZN(_00260_ ) );
AND2_X1 _19373_ ( .A1(\arbiter._io_axi_araddr_T_6 ), .A2(\io_master_rdata [23] ), .ZN(_12519_ ) );
AND4_X1 _19374_ ( .A1(_11949_ ), .A2(_11982_ ), .A3(_11976_ ), .A4(_12519_ ), .ZN(_12520_ ) );
AOI21_X1 _19375_ ( .A(_12520_ ), .B1(_11952_ ), .B2(\ifu.inst [23] ), .ZN(_12521_ ) );
MUX2_X1 _19376_ ( .A(\icache.icache_reg_0_0 [23] ), .B(\icache.icache_reg_0_1 [23] ), .S(_11910_ ), .Z(_12522_ ) );
MUX2_X1 _19377_ ( .A(\icache.icache_reg_0_2 [23] ), .B(_12522_ ), .S(_12000_ ), .Z(_12523_ ) );
MUX2_X1 _19378_ ( .A(\icache.icache_reg_0_3 [23] ), .B(_12523_ ), .S(_12005_ ), .Z(_12524_ ) );
MUX2_X1 _19379_ ( .A(\icache.icache_reg_1_0 [23] ), .B(_12524_ ), .S(_12052_ ), .Z(_12525_ ) );
MUX2_X1 _19380_ ( .A(\icache.icache_reg_1_1 [23] ), .B(_12525_ ), .S(_12054_ ), .Z(_12526_ ) );
MUX2_X1 _19381_ ( .A(\icache.icache_reg_1_2 [23] ), .B(_12526_ ), .S(_12056_ ), .Z(_12527_ ) );
MUX2_X1 _19382_ ( .A(\icache.icache_reg_1_3 [23] ), .B(_12527_ ), .S(_12143_ ), .Z(_12528_ ) );
AND4_X1 _19383_ ( .A1(\icache._io_out_arvalid_T ), .A2(_11901_ ), .A3(_11903_ ), .A4(_12528_ ), .ZN(_12529_ ) );
AOI22_X1 _19384_ ( .A1(_12528_ ), .A2(_11945_ ), .B1(_12519_ ), .B2(_11942_ ), .ZN(_12530_ ) );
AOI21_X1 _19385_ ( .A(_12530_ ), .B1(_12092_ ), .B2(\icache._io_out_arvalid_T ), .ZN(_12531_ ) );
OAI21_X1 _19386_ ( .A(_12358_ ), .B1(_12529_ ), .B2(_12531_ ), .ZN(_12532_ ) );
NAND2_X1 _19387_ ( .A1(_12521_ ), .A2(_12532_ ), .ZN(\ifu.io_out_bits_inst [23] ) );
AOI21_X1 _19388_ ( .A(fanout_net_22 ), .B1(_12521_ ), .B2(_12532_ ), .ZN(_00261_ ) );
AND2_X1 _19389_ ( .A1(\arbiter._io_axi_araddr_T_6 ), .A2(\io_master_rdata [22] ), .ZN(_12533_ ) );
AND4_X1 _19390_ ( .A1(_11949_ ), .A2(_11982_ ), .A3(_11976_ ), .A4(_12533_ ), .ZN(_12534_ ) );
AOI21_X1 _19391_ ( .A(_12534_ ), .B1(_11952_ ), .B2(\ifu.inst [22] ), .ZN(_12535_ ) );
NAND3_X1 _19392_ ( .A1(_11940_ ), .A2(_12533_ ), .A3(_11895_ ), .ZN(_12536_ ) );
AND4_X1 _19393_ ( .A1(\icache.icache_reg_1_3 [22] ), .A2(_12036_ ), .A3(_10839_ ), .A4(_11996_ ), .ZN(_12537_ ) );
MUX2_X1 _19394_ ( .A(\icache.icache_reg_0_0 [22] ), .B(\icache.icache_reg_0_1 [22] ), .S(_11911_ ), .Z(_12538_ ) );
MUX2_X1 _19395_ ( .A(\icache.icache_reg_0_2 [22] ), .B(_12538_ ), .S(_12001_ ), .Z(_12539_ ) );
MUX2_X1 _19396_ ( .A(\icache.icache_reg_0_3 [22] ), .B(_12539_ ), .S(_12006_ ), .Z(_12540_ ) );
MUX2_X1 _19397_ ( .A(\icache.icache_reg_1_0 [22] ), .B(_12540_ ), .S(_12052_ ), .Z(_12541_ ) );
MUX2_X1 _19398_ ( .A(\icache.icache_reg_1_1 [22] ), .B(_12541_ ), .S(_12054_ ), .Z(_12542_ ) );
MUX2_X1 _19399_ ( .A(\icache.icache_reg_1_2 [22] ), .B(_12542_ ), .S(_11927_ ), .Z(_12543_ ) );
AOI21_X1 _19400_ ( .A(_12537_ ), .B1(_12543_ ), .B2(_12012_ ), .ZN(_12544_ ) );
OR2_X1 _19401_ ( .A1(_12544_ ), .A2(_12014_ ), .ZN(_12545_ ) );
AOI22_X1 _19402_ ( .A1(_11991_ ), .A2(\icache._io_out_arvalid_T ), .B1(_12536_ ), .B2(_12545_ ), .ZN(_12546_ ) );
NOR4_X1 _19403_ ( .A1(_12017_ ), .A2(_12019_ ), .A3(_12020_ ), .A4(_12544_ ), .ZN(_12547_ ) );
OAI21_X1 _19404_ ( .A(_11989_ ), .B1(_12546_ ), .B2(_12547_ ), .ZN(_12548_ ) );
NAND2_X1 _19405_ ( .A1(_12535_ ), .A2(_12548_ ), .ZN(\ifu.io_out_bits_inst [22] ) );
AOI21_X1 _19406_ ( .A(fanout_net_22 ), .B1(_12535_ ), .B2(_12548_ ), .ZN(_00262_ ) );
AND2_X1 _19407_ ( .A1(_11401_ ), .A2(_11402_ ), .ZN(_12549_ ) );
AOI211_X1 _19408_ ( .A(fanout_net_22 ), .B(_12549_ ), .C1(_idu_io_in_bits_T ), .C2(_11899_ ), .ZN(_00263_ ) );
NOR2_X1 _19409_ ( .A1(_10701_ ), .A2(fanout_net_22 ), .ZN(_00264_ ) );
AND2_X1 _19410_ ( .A1(_10833_ ), .A2(_09775_ ), .ZN(_12550_ ) );
NAND2_X1 _19411_ ( .A1(_11429_ ), .A2(_11432_ ), .ZN(_12551_ ) );
INV_X1 _19412_ ( .A(_12551_ ), .ZN(_12552_ ) );
AND2_X1 _19413_ ( .A1(_11468_ ), .A2(_11474_ ), .ZN(_12553_ ) );
AND2_X1 _19414_ ( .A1(_12552_ ), .A2(_12553_ ), .ZN(_12554_ ) );
AND2_X1 _19415_ ( .A1(_09236_ ), .A2(_09239_ ), .ZN(_12555_ ) );
AND2_X1 _19416_ ( .A1(_12554_ ), .A2(_12555_ ), .ZN(_12556_ ) );
AND2_X1 _19417_ ( .A1(_10466_ ), .A2(_10470_ ), .ZN(_12557_ ) );
AND2_X1 _19418_ ( .A1(_12556_ ), .A2(_12557_ ), .ZN(_12558_ ) );
AND2_X1 _19419_ ( .A1(_10424_ ), .A2(_10427_ ), .ZN(_12559_ ) );
INV_X1 _19420_ ( .A(_12559_ ), .ZN(_12560_ ) );
NOR3_X1 _19421_ ( .A1(_10511_ ), .A2(_12560_ ), .A3(_10515_ ), .ZN(_12561_ ) );
AND2_X1 _19422_ ( .A1(_12558_ ), .A2(_12561_ ), .ZN(_12562_ ) );
NOR2_X1 _19423_ ( .A1(_10553_ ), .A2(_10556_ ), .ZN(_12563_ ) );
AND2_X1 _19424_ ( .A1(_12562_ ), .A2(_12563_ ), .ZN(_12564_ ) );
AND2_X1 _19425_ ( .A1(_10285_ ), .A2(_10290_ ), .ZN(_12565_ ) );
NOR2_X1 _19426_ ( .A1(_10238_ ), .A2(_10244_ ), .ZN(_12566_ ) );
AND3_X1 _19427_ ( .A1(_12564_ ), .A2(_12565_ ), .A3(_12566_ ), .ZN(_12567_ ) );
NOR2_X1 _19428_ ( .A1(_10383_ ), .A2(_10385_ ), .ZN(_12568_ ) );
NOR2_X1 _19429_ ( .A1(_10339_ ), .A2(_10344_ ), .ZN(_12569_ ) );
AND3_X1 _19430_ ( .A1(_12567_ ), .A2(_12568_ ), .A3(_12569_ ), .ZN(_12570_ ) );
NOR2_X1 _19431_ ( .A1(_10143_ ), .A2(_10147_ ), .ZN(_12571_ ) );
AND2_X1 _19432_ ( .A1(_10192_ ), .A2(_10196_ ), .ZN(_12572_ ) );
AND3_X1 _19433_ ( .A1(_12570_ ), .A2(_12571_ ), .A3(_12572_ ), .ZN(_12573_ ) );
NOR2_X1 _19434_ ( .A1(_09857_ ), .A2(_09864_ ), .ZN(_12574_ ) );
NOR2_X1 _19435_ ( .A1(_09907_ ), .A2(_09912_ ), .ZN(_12575_ ) );
AND3_X1 _19436_ ( .A1(_12573_ ), .A2(_12574_ ), .A3(_12575_ ), .ZN(_12576_ ) );
NOR2_X1 _19437_ ( .A1(_10092_ ), .A2(_10097_ ), .ZN(_12577_ ) );
NAND3_X1 _19438_ ( .A1(_12576_ ), .A2(_10007_ ), .A3(_12577_ ), .ZN(_12578_ ) );
NOR3_X1 _19439_ ( .A1(_12578_ ), .A2(_09956_ ), .A3(_09964_ ), .ZN(_12579_ ) );
NOR2_X1 _19440_ ( .A1(_10047_ ), .A2(_10051_ ), .ZN(_12580_ ) );
AND2_X1 _19441_ ( .A1(_12579_ ), .A2(_12580_ ), .ZN(_12581_ ) );
NOR2_X1 _19442_ ( .A1(_09599_ ), .A2(_09604_ ), .ZN(_12582_ ) );
AND2_X1 _19443_ ( .A1(_12581_ ), .A2(_12582_ ), .ZN(_12583_ ) );
NOR2_X1 _19444_ ( .A1(_09552_ ), .A2(_09556_ ), .ZN(_12584_ ) );
AND2_X1 _19445_ ( .A1(_12583_ ), .A2(_12584_ ), .ZN(_12585_ ) );
NOR2_X1 _19446_ ( .A1(_09512_ ), .A2(_09518_ ), .ZN(_12586_ ) );
AND2_X1 _19447_ ( .A1(_12585_ ), .A2(_12586_ ), .ZN(_12587_ ) );
NOR2_X1 _19448_ ( .A1(_09642_ ), .A2(_09644_ ), .ZN(_12588_ ) );
AND2_X1 _19449_ ( .A1(_12587_ ), .A2(_12588_ ), .ZN(_12589_ ) );
NOR2_X1 _19450_ ( .A1(_09320_ ), .A2(_09326_ ), .ZN(_12590_ ) );
AND2_X1 _19451_ ( .A1(_12589_ ), .A2(_12590_ ), .ZN(_12591_ ) );
NOR2_X1 _19452_ ( .A1(_08992_ ), .A2(_09178_ ), .ZN(_12592_ ) );
AND2_X1 _19453_ ( .A1(_12591_ ), .A2(_12592_ ), .ZN(_12593_ ) );
NOR2_X1 _19454_ ( .A1(_09381_ ), .A2(_09398_ ), .ZN(_12594_ ) );
AND2_X1 _19455_ ( .A1(_09457_ ), .A2(_09464_ ), .ZN(_12595_ ) );
AND3_X1 _19456_ ( .A1(_12593_ ), .A2(_12594_ ), .A3(_12595_ ), .ZN(_12596_ ) );
AND2_X1 _19457_ ( .A1(_09698_ ), .A2(_09711_ ), .ZN(_12597_ ) );
INV_X1 _19458_ ( .A(_12597_ ), .ZN(_12598_ ) );
OR2_X1 _19459_ ( .A1(_09812_ ), .A2(\exu.io_in_bits_jalr ), .ZN(_12599_ ) );
AND2_X1 _19460_ ( .A1(_12599_ ), .A2(_09779_ ), .ZN(_12600_ ) );
INV_X1 _19461_ ( .A(_12600_ ), .ZN(_12601_ ) );
AND3_X1 _19462_ ( .A1(_12596_ ), .A2(_12598_ ), .A3(_12601_ ), .ZN(_12602_ ) );
NOR2_X1 _19463_ ( .A1(_09763_ ), .A2(_09768_ ), .ZN(_12603_ ) );
NOR2_X1 _19464_ ( .A1(_12602_ ), .A2(_12603_ ), .ZN(_12604_ ) );
AND4_X1 _19465_ ( .A1(_12603_ ), .A2(_12596_ ), .A3(_12598_ ), .A4(_12601_ ), .ZN(_12605_ ) );
OAI21_X1 _19466_ ( .A(_12550_ ), .B1(_12604_ ), .B2(_12605_ ), .ZN(_12606_ ) );
AND3_X1 _19467_ ( .A1(\ifu.pc [5] ), .A2(\ifu.pc [3] ), .A3(\ifu.pc [2] ), .ZN(_12607_ ) );
AND2_X2 _19468_ ( .A1(_12607_ ), .A2(\ifu.pc [4] ), .ZN(_12608_ ) );
AND2_X1 _19469_ ( .A1(\ifu.pc [7] ), .A2(\ifu.pc [6] ), .ZN(_12609_ ) );
AND2_X1 _19470_ ( .A1(_12608_ ), .A2(_12609_ ), .ZN(_12610_ ) );
AND4_X1 _19471_ ( .A1(\ifu.pc [11] ), .A2(_12610_ ), .A3(\ifu.pc [9] ), .A4(\ifu.pc [8] ), .ZN(_12611_ ) );
AND3_X1 _19472_ ( .A1(_12611_ ), .A2(\ifu.pc [13] ), .A3(\ifu.pc [10] ), .ZN(_12612_ ) );
AND3_X1 _19473_ ( .A1(_12612_ ), .A2(\ifu.pc [14] ), .A3(\ifu.pc [12] ), .ZN(_12613_ ) );
NAND3_X1 _19474_ ( .A1(_12613_ ), .A2(\ifu.pc [16] ), .A3(\ifu.pc [15] ), .ZN(_12614_ ) );
NOR3_X1 _19475_ ( .A1(_12614_ ), .A2(_10011_ ), .A3(_10099_ ), .ZN(_12615_ ) );
NAND3_X1 _19476_ ( .A1(_12615_ ), .A2(\ifu.pc [20] ), .A3(\ifu.pc [19] ), .ZN(_12616_ ) );
NOR2_X1 _19477_ ( .A1(_12616_ ), .A2(_09606_ ), .ZN(_12617_ ) );
AND4_X1 _19478_ ( .A1(\ifu.pc [22] ), .A2(_12617_ ), .A3(\ifu.pc [25] ), .A4(\ifu.pc [23] ), .ZN(_12618_ ) );
AND3_X1 _19479_ ( .A1(_12618_ ), .A2(\ifu.pc [27] ), .A3(\ifu.pc [24] ), .ZN(_12619_ ) );
NAND3_X1 _19480_ ( .A1(_12619_ ), .A2(\ifu.pc [28] ), .A3(\ifu.pc [26] ), .ZN(_12620_ ) );
NOR3_X1 _19481_ ( .A1(_12620_ ), .A2(_09713_ ), .A3(_09814_ ), .ZN(_12621_ ) );
XNOR2_X1 _19482_ ( .A(_12621_ ), .B(\ifu.pc [31] ), .ZN(_12622_ ) );
OAI221_X1 _19483_ ( .A(_10831_ ), .B1(_09775_ ), .B2(_12622_ ), .C1(_10711_ ), .C2(\ifu.state [2] ), .ZN(_12623_ ) );
AND2_X2 _19484_ ( .A1(_10833_ ), .A2(_09040_ ), .ZN(_12624_ ) );
BUF_X4 _19485_ ( .A(_12624_ ), .Z(_12625_ ) );
INV_X1 _19486_ ( .A(_11973_ ), .ZN(\ifu.io_out_bits_pc [31] ) );
OAI21_X1 _19487_ ( .A(_12623_ ), .B1(_12625_ ), .B2(\ifu.io_out_bits_pc [31] ), .ZN(_12626_ ) );
AOI21_X1 _19488_ ( .A(fanout_net_22 ), .B1(_12606_ ), .B2(_12626_ ), .ZN(_00265_ ) );
BUF_X4 _19489_ ( .A(_09775_ ), .Z(_12627_ ) );
NOR2_X1 _19490_ ( .A1(_12620_ ), .A2(_09814_ ), .ZN(_12628_ ) );
XNOR2_X1 _19491_ ( .A(_12628_ ), .B(\ifu.pc [30] ), .ZN(_12629_ ) );
OAI221_X1 _19492_ ( .A(_10831_ ), .B1(_12627_ ), .B2(_12629_ ), .C1(_10711_ ), .C2(\ifu.state [2] ), .ZN(_12630_ ) );
BUF_X4 _19493_ ( .A(_12624_ ), .Z(_12631_ ) );
INV_X1 _19494_ ( .A(_11970_ ), .ZN(\ifu.io_out_bits_pc [30] ) );
OAI21_X1 _19495_ ( .A(_12630_ ), .B1(_12631_ ), .B2(\ifu.io_out_bits_pc [30] ), .ZN(_12632_ ) );
INV_X1 _19496_ ( .A(_12602_ ), .ZN(_12633_ ) );
NAND2_X1 _19497_ ( .A1(_12596_ ), .A2(_12601_ ), .ZN(_12634_ ) );
NAND2_X1 _19498_ ( .A1(_12634_ ), .A2(_12597_ ), .ZN(_12635_ ) );
NAND3_X1 _19499_ ( .A1(_12633_ ), .A2(_12550_ ), .A3(_12635_ ), .ZN(_12636_ ) );
AOI21_X1 _19500_ ( .A(fanout_net_22 ), .B1(_12632_ ), .B2(_12636_ ), .ZN(_00266_ ) );
AND4_X1 _19501_ ( .A1(\ifu.pc [9] ), .A2(\ifu.pc [8] ), .A3(\ifu.pc [7] ), .A4(\ifu.pc [6] ), .ZN(_12637_ ) );
AND2_X2 _19502_ ( .A1(_12608_ ), .A2(_12637_ ), .ZN(_12638_ ) );
AND4_X1 _19503_ ( .A1(\ifu.pc [14] ), .A2(\ifu.pc [16] ), .A3(\ifu.pc [15] ), .A4(\ifu.pc [17] ), .ZN(_12639_ ) );
AND2_X1 _19504_ ( .A1(\ifu.pc [11] ), .A2(\ifu.pc [10] ), .ZN(_12640_ ) );
AND4_X1 _19505_ ( .A1(\ifu.pc [13] ), .A2(_12639_ ), .A3(\ifu.pc [12] ), .A4(_12640_ ), .ZN(_12641_ ) );
NAND3_X1 _19506_ ( .A1(_12638_ ), .A2(\ifu.pc [18] ), .A3(_12641_ ), .ZN(_12642_ ) );
XNOR2_X1 _19507_ ( .A(_12642_ ), .B(\ifu.pc [19] ), .ZN(_12643_ ) );
AND2_X1 _19508_ ( .A1(_09965_ ), .A2(_09966_ ), .ZN(_12644_ ) );
INV_X1 _19509_ ( .A(_12644_ ), .ZN(\ifu.io_out_bits_pc [19] ) );
INV_X2 _19510_ ( .A(_10833_ ), .ZN(_12645_ ) );
BUF_X4 _19511_ ( .A(_12645_ ), .Z(_12646_ ) );
AOI22_X1 _19512_ ( .A1(_12631_ ), .A2(_12643_ ), .B1(\ifu.io_out_bits_pc [19] ), .B2(_12646_ ), .ZN(_12647_ ) );
BUF_X4 _19513_ ( .A(_12627_ ), .Z(_12648_ ) );
INV_X1 _19514_ ( .A(_12579_ ), .ZN(_12649_ ) );
OAI21_X1 _19515_ ( .A(_12578_ ), .B1(_09956_ ), .B2(_09964_ ), .ZN(_12650_ ) );
NAND4_X1 _19516_ ( .A1(_idu_io_in_bits_T ), .A2(_12648_ ), .A3(_12649_ ), .A4(_12650_ ), .ZN(_12651_ ) );
AOI21_X1 _19517_ ( .A(fanout_net_22 ), .B1(_12647_ ), .B2(_12651_ ), .ZN(_00267_ ) );
AND2_X1 _19518_ ( .A1(_12638_ ), .A2(_12641_ ), .ZN(_12652_ ) );
XNOR2_X1 _19519_ ( .A(_12652_ ), .B(_10011_ ), .ZN(_12653_ ) );
AND2_X1 _19520_ ( .A1(_10008_ ), .A2(_10009_ ), .ZN(_12654_ ) );
INV_X1 _19521_ ( .A(_12654_ ), .ZN(\ifu.io_out_bits_pc [18] ) );
AOI22_X1 _19522_ ( .A1(_12631_ ), .A2(_12653_ ), .B1(\ifu.io_out_bits_pc [18] ), .B2(_12646_ ), .ZN(_12655_ ) );
INV_X1 _19523_ ( .A(_10712_ ), .ZN(_12656_ ) );
BUF_X4 _19524_ ( .A(_12656_ ), .Z(_12657_ ) );
BUF_X4 _19525_ ( .A(_10831_ ), .Z(_12658_ ) );
NAND2_X1 _19526_ ( .A1(_12576_ ), .A2(_12577_ ), .ZN(_12659_ ) );
XNOR2_X1 _19527_ ( .A(_12659_ ), .B(_10007_ ), .ZN(_12660_ ) );
NAND4_X1 _19528_ ( .A1(_12657_ ), .A2(_12658_ ), .A3(_12648_ ), .A4(_12660_ ), .ZN(_12661_ ) );
AOI21_X1 _19529_ ( .A(fanout_net_22 ), .B1(_12655_ ), .B2(_12661_ ), .ZN(_00268_ ) );
AND3_X1 _19530_ ( .A1(_12640_ ), .A2(\ifu.pc [13] ), .A3(\ifu.pc [12] ), .ZN(_12662_ ) );
AND2_X1 _19531_ ( .A1(_12638_ ), .A2(_12662_ ), .ZN(_12663_ ) );
NAND3_X1 _19532_ ( .A1(_12663_ ), .A2(\ifu.pc [14] ), .A3(\ifu.pc [15] ), .ZN(_12664_ ) );
NOR2_X1 _19533_ ( .A1(_12664_ ), .A2(_09916_ ), .ZN(_12665_ ) );
XNOR2_X1 _19534_ ( .A(_12665_ ), .B(_10099_ ), .ZN(_12666_ ) );
INV_X1 _19535_ ( .A(_10101_ ), .ZN(\ifu.io_out_bits_pc [17] ) );
AOI22_X1 _19536_ ( .A1(_12631_ ), .A2(_12666_ ), .B1(\ifu.io_out_bits_pc [17] ), .B2(_12646_ ), .ZN(_12667_ ) );
AND4_X1 _19537_ ( .A1(_12563_ ), .A2(_10285_ ), .A3(_10290_ ), .A4(_12561_ ), .ZN(_12668_ ) );
AND2_X1 _19538_ ( .A1(_12558_ ), .A2(_12668_ ), .ZN(_12669_ ) );
AND2_X1 _19539_ ( .A1(_12569_ ), .A2(_12566_ ), .ZN(_12670_ ) );
AND3_X1 _19540_ ( .A1(_12670_ ), .A2(_12568_ ), .A3(_12572_ ), .ZN(_12671_ ) );
AND2_X1 _19541_ ( .A1(_12669_ ), .A2(_12671_ ), .ZN(_12672_ ) );
AND3_X1 _19542_ ( .A1(_12574_ ), .A2(_12672_ ), .A3(_12571_ ), .ZN(_12673_ ) );
NAND2_X1 _19543_ ( .A1(_12673_ ), .A2(_12575_ ), .ZN(_12674_ ) );
XNOR2_X1 _19544_ ( .A(_12674_ ), .B(_12577_ ), .ZN(_12675_ ) );
NAND4_X1 _19545_ ( .A1(_12657_ ), .A2(_12658_ ), .A3(_12648_ ), .A4(_12675_ ), .ZN(_12676_ ) );
AOI21_X1 _19546_ ( .A(fanout_net_22 ), .B1(_12667_ ), .B2(_12676_ ), .ZN(_00269_ ) );
XNOR2_X1 _19547_ ( .A(_12664_ ), .B(\ifu.pc [16] ), .ZN(_12677_ ) );
AND2_X1 _19548_ ( .A1(_09913_ ), .A2(_09914_ ), .ZN(_12678_ ) );
INV_X1 _19549_ ( .A(_12678_ ), .ZN(\ifu.io_out_bits_pc [16] ) );
AOI22_X1 _19550_ ( .A1(_12631_ ), .A2(_12677_ ), .B1(\ifu.io_out_bits_pc [16] ), .B2(_12646_ ), .ZN(_12679_ ) );
NAND3_X1 _19551_ ( .A1(_12574_ ), .A2(_12672_ ), .A3(_12571_ ), .ZN(_12680_ ) );
XNOR2_X1 _19552_ ( .A(_12680_ ), .B(_12575_ ), .ZN(_12681_ ) );
NAND4_X1 _19553_ ( .A1(_12657_ ), .A2(_12658_ ), .A3(_12648_ ), .A4(_12681_ ), .ZN(_12682_ ) );
AOI21_X1 _19554_ ( .A(fanout_net_22 ), .B1(_12679_ ), .B2(_12682_ ), .ZN(_00270_ ) );
NAND3_X1 _19555_ ( .A1(_12638_ ), .A2(\ifu.pc [14] ), .A3(_12662_ ), .ZN(_12683_ ) );
XNOR2_X1 _19556_ ( .A(_12683_ ), .B(\ifu.pc [15] ), .ZN(_12684_ ) );
AND2_X1 _19557_ ( .A1(_09865_ ), .A2(_09866_ ), .ZN(_12685_ ) );
INV_X1 _19558_ ( .A(_12685_ ), .ZN(\ifu.io_out_bits_pc [15] ) );
AOI22_X1 _19559_ ( .A1(_12631_ ), .A2(_12684_ ), .B1(\ifu.io_out_bits_pc [15] ), .B2(_12646_ ), .ZN(_12686_ ) );
NAND3_X1 _19560_ ( .A1(_12669_ ), .A2(_12571_ ), .A3(_12671_ ), .ZN(_12687_ ) );
XNOR2_X1 _19561_ ( .A(_12574_ ), .B(_12687_ ), .ZN(_12688_ ) );
NAND4_X1 _19562_ ( .A1(_12657_ ), .A2(_12658_ ), .A3(_12648_ ), .A4(_12688_ ), .ZN(_12689_ ) );
AOI21_X1 _19563_ ( .A(fanout_net_22 ), .B1(_12686_ ), .B2(_12689_ ), .ZN(_00271_ ) );
XNOR2_X1 _19564_ ( .A(_12663_ ), .B(_10151_ ), .ZN(_12690_ ) );
AND2_X1 _19565_ ( .A1(_10148_ ), .A2(_10149_ ), .ZN(_12691_ ) );
INV_X1 _19566_ ( .A(_12691_ ), .ZN(\ifu.io_out_bits_pc [14] ) );
AOI22_X1 _19567_ ( .A1(_12631_ ), .A2(_12690_ ), .B1(\ifu.io_out_bits_pc [14] ), .B2(_12646_ ), .ZN(_12692_ ) );
XOR2_X1 _19568_ ( .A(_12672_ ), .B(_12571_ ), .Z(_12693_ ) );
NAND4_X1 _19569_ ( .A1(_12657_ ), .A2(_12658_ ), .A3(_12648_ ), .A4(_12693_ ), .ZN(_12694_ ) );
AOI21_X1 _19570_ ( .A(fanout_net_22 ), .B1(_12692_ ), .B2(_12694_ ), .ZN(_00272_ ) );
NAND3_X1 _19571_ ( .A1(_12608_ ), .A2(_12640_ ), .A3(_12637_ ), .ZN(_12695_ ) );
NOR2_X1 _19572_ ( .A1(_12695_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_5_A_$_MUX__Y_B ), .ZN(_12696_ ) );
XNOR2_X1 _19573_ ( .A(_12696_ ), .B(_10200_ ), .ZN(_12697_ ) );
AND2_X1 _19574_ ( .A1(_10197_ ), .A2(_10198_ ), .ZN(_12698_ ) );
INV_X1 _19575_ ( .A(_12698_ ), .ZN(\ifu.io_out_bits_pc [13] ) );
BUF_X4 _19576_ ( .A(_12645_ ), .Z(_12699_ ) );
AOI22_X1 _19577_ ( .A1(_12631_ ), .A2(_12697_ ), .B1(\ifu.io_out_bits_pc [13] ), .B2(_12699_ ), .ZN(_12700_ ) );
NAND3_X1 _19578_ ( .A1(_12669_ ), .A2(_12568_ ), .A3(_12670_ ), .ZN(_12701_ ) );
XNOR2_X1 _19579_ ( .A(_12701_ ), .B(_12572_ ), .ZN(_12702_ ) );
NAND4_X1 _19580_ ( .A1(_12657_ ), .A2(_12658_ ), .A3(_12648_ ), .A4(_12702_ ), .ZN(_12703_ ) );
AOI21_X1 _19581_ ( .A(fanout_net_22 ), .B1(_12700_ ), .B2(_12703_ ), .ZN(_00273_ ) );
AOI21_X1 _19582_ ( .A(_12568_ ), .B1(_12567_ ), .B2(_12569_ ), .ZN(_12704_ ) );
OR4_X1 _19583_ ( .A1(_11899_ ), .A2(_12645_ ), .A3(_12570_ ), .A4(_12704_ ), .ZN(_12705_ ) );
XNOR2_X1 _19584_ ( .A(_12695_ ), .B(\ifu.pc [12] ), .ZN(_12706_ ) );
NAND2_X1 _19585_ ( .A1(_10386_ ), .A2(_10387_ ), .ZN(\ifu.io_out_bits_pc [12] ) );
AOI22_X1 _19586_ ( .A1(_12625_ ), .A2(_12706_ ), .B1(\ifu.io_out_bits_pc [12] ), .B2(_12699_ ), .ZN(_12707_ ) );
AOI21_X1 _19587_ ( .A(fanout_net_22 ), .B1(_12705_ ), .B2(_12707_ ), .ZN(_00274_ ) );
NAND3_X1 _19588_ ( .A1(_12608_ ), .A2(_10246_ ), .A3(_12637_ ), .ZN(_12708_ ) );
XNOR2_X1 _19589_ ( .A(_12708_ ), .B(\ifu.pc [11] ), .ZN(_12709_ ) );
NAND2_X1 _19590_ ( .A1(_10345_ ), .A2(_10346_ ), .ZN(\ifu.io_out_bits_pc [11] ) );
AOI22_X1 _19591_ ( .A1(_12625_ ), .A2(_12709_ ), .B1(\ifu.io_out_bits_pc [11] ), .B2(_12699_ ), .ZN(_12710_ ) );
XOR2_X1 _19592_ ( .A(_12567_ ), .B(_12569_ ), .Z(_12711_ ) );
NAND4_X1 _19593_ ( .A1(_12657_ ), .A2(_12658_ ), .A3(_12627_ ), .A4(_12711_ ), .ZN(_12712_ ) );
AOI21_X1 _19594_ ( .A(fanout_net_22 ), .B1(_12710_ ), .B2(_12712_ ), .ZN(_00275_ ) );
XOR2_X1 _19595_ ( .A(_12638_ ), .B(\ifu.pc [10] ), .Z(_12713_ ) );
NAND2_X1 _19596_ ( .A1(_10245_ ), .A2(_10247_ ), .ZN(\ifu.io_out_bits_pc [10] ) );
AOI22_X1 _19597_ ( .A1(_12625_ ), .A2(_12713_ ), .B1(\ifu.io_out_bits_pc [10] ), .B2(_12699_ ), .ZN(_12714_ ) );
XOR2_X1 _19598_ ( .A(_12669_ ), .B(_12566_ ), .Z(_12715_ ) );
NAND4_X1 _19599_ ( .A1(_12657_ ), .A2(_12658_ ), .A3(_12627_ ), .A4(_12715_ ), .ZN(_12716_ ) );
AOI21_X1 _19600_ ( .A(fanout_net_22 ), .B1(_12714_ ), .B2(_12716_ ), .ZN(_00276_ ) );
INV_X1 _19601_ ( .A(_12652_ ), .ZN(_12717_ ) );
AND4_X1 _19602_ ( .A1(\ifu.pc [22] ), .A2(\ifu.pc [25] ), .A3(\ifu.pc [24] ), .A4(\ifu.pc [23] ), .ZN(_12718_ ) );
AND2_X1 _19603_ ( .A1(\ifu.pc [19] ), .A2(\ifu.pc [18] ), .ZN(_12719_ ) );
NAND4_X1 _19604_ ( .A1(_12718_ ), .A2(\ifu.pc [21] ), .A3(\ifu.pc [20] ), .A4(_12719_ ), .ZN(_12720_ ) );
OR3_X1 _19605_ ( .A1(_12717_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_1_A_$_MUX__Y_B ), .A3(_12720_ ), .ZN(_12721_ ) );
XNOR2_X1 _19606_ ( .A(_12721_ ), .B(\ifu.pc [27] ), .ZN(_12722_ ) );
NAND2_X1 _19607_ ( .A1(_09465_ ), .A2(_09467_ ), .ZN(\ifu.io_out_bits_pc [27] ) );
AOI22_X1 _19608_ ( .A1(_12625_ ), .A2(_12722_ ), .B1(\ifu.io_out_bits_pc [27] ), .B2(_12699_ ), .ZN(_12723_ ) );
AND2_X1 _19609_ ( .A1(_12593_ ), .A2(_12595_ ), .ZN(_12724_ ) );
NOR4_X1 _19610_ ( .A1(_10712_ ), .A2(_12724_ ), .A3(_10832_ ), .A4(_11899_ ), .ZN(_12725_ ) );
OAI21_X1 _19611_ ( .A(_12725_ ), .B1(_12595_ ), .B2(_12593_ ), .ZN(_12726_ ) );
AOI21_X1 _19612_ ( .A(fanout_net_22 ), .B1(_12723_ ), .B2(_12726_ ), .ZN(_00277_ ) );
AOI211_X1 _19613_ ( .A(_11899_ ), .B(_12645_ ), .C1(_12565_ ), .C2(_12564_ ), .ZN(_12727_ ) );
OAI21_X1 _19614_ ( .A(_12727_ ), .B1(_12565_ ), .B2(_12564_ ), .ZN(_12728_ ) );
INV_X1 _19615_ ( .A(_12610_ ), .ZN(_12729_ ) );
OR2_X1 _19616_ ( .A1(_12729_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_9_A_$_MUX__Y_B ), .ZN(_12730_ ) );
XNOR2_X1 _19617_ ( .A(_12730_ ), .B(\ifu.pc [9] ), .ZN(_12731_ ) );
OR2_X1 _19618_ ( .A1(_10291_ ), .A2(_10292_ ), .ZN(\ifu.io_out_bits_pc [9] ) );
AOI22_X1 _19619_ ( .A1(_12625_ ), .A2(_12731_ ), .B1(\ifu.io_out_bits_pc [9] ), .B2(_12699_ ), .ZN(_12732_ ) );
AOI21_X1 _19620_ ( .A(fanout_net_22 ), .B1(_12728_ ), .B2(_12732_ ), .ZN(_00278_ ) );
BUF_X2 _19621_ ( .A(_10833_ ), .Z(_12733_ ) );
OAI211_X1 _19622_ ( .A(_12733_ ), .B(_12627_ ), .C1(_12563_ ), .C2(_12562_ ), .ZN(_12734_ ) );
OR2_X1 _19623_ ( .A1(_12734_ ), .A2(_12564_ ), .ZN(_12735_ ) );
XOR2_X1 _19624_ ( .A(_12610_ ), .B(\ifu.pc [8] ), .Z(_12736_ ) );
NAND2_X1 _19625_ ( .A1(_10557_ ), .A2(_10558_ ), .ZN(\ifu.io_out_bits_pc [8] ) );
AOI22_X1 _19626_ ( .A1(_12625_ ), .A2(_12736_ ), .B1(\ifu.io_out_bits_pc [8] ), .B2(_12699_ ), .ZN(_12737_ ) );
AOI21_X1 _19627_ ( .A(fanout_net_22 ), .B1(_12735_ ), .B2(_12737_ ), .ZN(_00279_ ) );
NAND2_X1 _19628_ ( .A1(_12608_ ), .A2(_10429_ ), .ZN(_12738_ ) );
XNOR2_X1 _19629_ ( .A(_12738_ ), .B(\ifu.pc [7] ), .ZN(_12739_ ) );
NAND2_X1 _19630_ ( .A1(_10516_ ), .A2(_10517_ ), .ZN(\ifu.io_out_bits_pc [7] ) );
AOI22_X1 _19631_ ( .A1(_12625_ ), .A2(_12739_ ), .B1(\ifu.io_out_bits_pc [7] ), .B2(_12699_ ), .ZN(_12740_ ) );
NAND2_X1 _19632_ ( .A1(_12558_ ), .A2(_12559_ ), .ZN(_12741_ ) );
OAI21_X1 _19633_ ( .A(_12741_ ), .B1(_10515_ ), .B2(_10511_ ), .ZN(_12742_ ) );
NAND4_X1 _19634_ ( .A1(_12656_ ), .A2(_10831_ ), .A3(_09775_ ), .A4(_12742_ ), .ZN(_12743_ ) );
OR2_X1 _19635_ ( .A1(_12743_ ), .A2(_12562_ ), .ZN(_12744_ ) );
AOI21_X1 _19636_ ( .A(fanout_net_22 ), .B1(_12740_ ), .B2(_12744_ ), .ZN(_00280_ ) );
XNOR2_X1 _19637_ ( .A(_12608_ ), .B(\ifu.pc [6] ), .ZN(_12745_ ) );
OAI221_X1 _19638_ ( .A(_10831_ ), .B1(_12627_ ), .B2(_12745_ ), .C1(_10711_ ), .C2(\ifu.state [2] ), .ZN(_12746_ ) );
NAND2_X1 _19639_ ( .A1(_10428_ ), .A2(_10430_ ), .ZN(\ifu.io_out_bits_pc [6] ) );
OAI21_X1 _19640_ ( .A(_12746_ ), .B1(_12631_ ), .B2(\ifu.io_out_bits_pc [6] ), .ZN(_12747_ ) );
XNOR2_X1 _19641_ ( .A(_12558_ ), .B(_12560_ ), .ZN(_12748_ ) );
NAND4_X1 _19642_ ( .A1(_12657_ ), .A2(_12658_ ), .A3(_12627_ ), .A4(_12748_ ), .ZN(_12749_ ) );
AOI21_X1 _19643_ ( .A(fanout_net_22 ), .B1(_12747_ ), .B2(_12749_ ), .ZN(_00281_ ) );
OAI211_X1 _19644_ ( .A(_12733_ ), .B(_12627_ ), .C1(_12557_ ), .C2(_12556_ ), .ZN(_12750_ ) );
OR2_X1 _19645_ ( .A1(_12750_ ), .A2(_12558_ ), .ZN(_12751_ ) );
AND2_X1 _19646_ ( .A1(\ifu.pc [3] ), .A2(\ifu.pc [2] ), .ZN(_12752_ ) );
NAND2_X1 _19647_ ( .A1(_12752_ ), .A2(_09241_ ), .ZN(_12753_ ) );
XNOR2_X1 _19648_ ( .A(_12753_ ), .B(\ifu.pc [5] ), .ZN(_12754_ ) );
OR2_X1 _19649_ ( .A1(_10471_ ), .A2(_10472_ ), .ZN(\ifu.io_out_bits_pc [5] ) );
AOI22_X1 _19650_ ( .A1(_12625_ ), .A2(_12754_ ), .B1(\ifu.io_out_bits_pc [5] ), .B2(_12699_ ), .ZN(_12755_ ) );
AOI21_X1 _19651_ ( .A(fanout_net_22 ), .B1(_12751_ ), .B2(_12755_ ), .ZN(_00282_ ) );
OAI211_X1 _19652_ ( .A(_12733_ ), .B(_12627_ ), .C1(_12555_ ), .C2(_12554_ ), .ZN(_12756_ ) );
OR2_X1 _19653_ ( .A1(_12756_ ), .A2(_12556_ ), .ZN(_12757_ ) );
XOR2_X1 _19654_ ( .A(_12752_ ), .B(\ifu.pc [4] ), .Z(_12758_ ) );
AOI22_X1 _19655_ ( .A1(_12625_ ), .A2(_12758_ ), .B1(\ifu.io_out_bits_pc [4] ), .B2(_12645_ ), .ZN(_12759_ ) );
AOI21_X1 _19656_ ( .A(fanout_net_22 ), .B1(_12757_ ), .B2(_12759_ ), .ZN(_00283_ ) );
AOI21_X1 _19657_ ( .A(_12553_ ), .B1(_11429_ ), .B2(_11432_ ), .ZN(_12760_ ) );
OR4_X1 _19658_ ( .A1(_11899_ ), .A2(_12645_ ), .A3(_12554_ ), .A4(_12760_ ), .ZN(_12761_ ) );
XOR2_X1 _19659_ ( .A(\ifu.pc [3] ), .B(\ifu.pc [2] ), .Z(_12762_ ) );
NAND2_X1 _19660_ ( .A1(_11475_ ), .A2(_11476_ ), .ZN(\ifu.io_out_bits_pc [3] ) );
AOI22_X1 _19661_ ( .A1(_12624_ ), .A2(_12762_ ), .B1(_12699_ ), .B2(\ifu.io_out_bits_pc [3] ), .ZN(_12763_ ) );
AOI21_X1 _19662_ ( .A(fanout_net_22 ), .B1(_12761_ ), .B2(_12763_ ), .ZN(_00284_ ) );
NAND2_X1 _19663_ ( .A1(_11433_ ), .A2(_11434_ ), .ZN(\ifu.io_out_bits_pc [2] ) );
OAI21_X1 _19664_ ( .A(_10922_ ), .B1(_idu_io_in_bits_T ), .B2(\ifu.io_out_bits_pc [2] ), .ZN(_12764_ ) );
AOI21_X1 _19665_ ( .A(_12764_ ), .B1(_idu_io_in_bits_T ), .B2(\ifu.io_out_bits_pc [2] ), .ZN(_00285_ ) );
OAI211_X1 _19666_ ( .A(_12733_ ), .B(_12627_ ), .C1(_12592_ ), .C2(_12591_ ), .ZN(_12765_ ) );
OR2_X1 _19667_ ( .A1(_12765_ ), .A2(_12593_ ), .ZN(_12766_ ) );
OR2_X1 _19668_ ( .A1(_12717_ ), .A2(_12720_ ), .ZN(_12767_ ) );
XNOR2_X1 _19669_ ( .A(_12767_ ), .B(\ifu.pc [26] ), .ZN(_12768_ ) );
NAND2_X1 _19670_ ( .A1(_09179_ ), .A2(_09186_ ), .ZN(\ifu.io_out_bits_pc [26] ) );
AOI22_X1 _19671_ ( .A1(_12624_ ), .A2(_12768_ ), .B1(\ifu.io_out_bits_pc [26] ), .B2(_12645_ ), .ZN(_12769_ ) );
AOI21_X1 _19672_ ( .A(fanout_net_22 ), .B1(_12766_ ), .B2(_12769_ ), .ZN(_00286_ ) );
AND3_X1 _19673_ ( .A1(_12719_ ), .A2(\ifu.pc [21] ), .A3(\ifu.pc [20] ), .ZN(_12770_ ) );
AND2_X1 _19674_ ( .A1(_12652_ ), .A2(_12770_ ), .ZN(_12771_ ) );
AND3_X1 _19675_ ( .A1(_12771_ ), .A2(\ifu.pc [22] ), .A3(\ifu.pc [23] ), .ZN(_12772_ ) );
NAND2_X1 _19676_ ( .A1(_12772_ ), .A2(_09648_ ), .ZN(_12773_ ) );
XNOR2_X1 _19677_ ( .A(_12773_ ), .B(\ifu.pc [25] ), .ZN(_12774_ ) );
AND3_X1 _19678_ ( .A1(_12733_ ), .A2(_11899_ ), .A3(_12774_ ), .ZN(_12775_ ) );
NAND2_X1 _19679_ ( .A1(_09327_ ), .A2(_09329_ ), .ZN(\ifu.io_out_bits_pc [25] ) );
AOI21_X1 _19680_ ( .A(_12775_ ), .B1(\ifu.io_out_bits_pc [25] ), .B2(_12646_ ), .ZN(_12776_ ) );
OAI211_X1 _19681_ ( .A(_12733_ ), .B(_09775_ ), .C1(_12590_ ), .C2(_12589_ ), .ZN(_12777_ ) );
OR2_X1 _19682_ ( .A1(_12777_ ), .A2(_12591_ ), .ZN(_12778_ ) );
AOI21_X1 _19683_ ( .A(fanout_net_22 ), .B1(_12776_ ), .B2(_12778_ ), .ZN(_00287_ ) );
OAI211_X1 _19684_ ( .A(_12733_ ), .B(_09775_ ), .C1(_12588_ ), .C2(_12587_ ), .ZN(_12779_ ) );
OR2_X1 _19685_ ( .A1(_12779_ ), .A2(_12589_ ), .ZN(_12780_ ) );
XOR2_X1 _19686_ ( .A(_12772_ ), .B(\ifu.pc [24] ), .Z(_12781_ ) );
AND2_X1 _19687_ ( .A1(_09645_ ), .A2(_09646_ ), .ZN(\ifu.io_out_bits_pc [24] ) );
AOI22_X1 _19688_ ( .A1(_12624_ ), .A2(_12781_ ), .B1(\ifu.io_out_bits_pc [24] ), .B2(_12645_ ), .ZN(_12782_ ) );
AOI21_X1 _19689_ ( .A(fanout_net_22 ), .B1(_12780_ ), .B2(_12782_ ), .ZN(_00288_ ) );
OAI211_X1 _19690_ ( .A(_12733_ ), .B(_09775_ ), .C1(_12586_ ), .C2(_12585_ ), .ZN(_12783_ ) );
OR2_X1 _19691_ ( .A1(_12783_ ), .A2(_12587_ ), .ZN(_12784_ ) );
NAND3_X1 _19692_ ( .A1(_12652_ ), .A2(\ifu.pc [22] ), .A3(_12770_ ), .ZN(_12785_ ) );
XNOR2_X1 _19693_ ( .A(_12785_ ), .B(\ifu.pc [23] ), .ZN(_12786_ ) );
NAND2_X1 _19694_ ( .A1(_09519_ ), .A2(_09520_ ), .ZN(\ifu.io_out_bits_pc [23] ) );
AOI22_X1 _19695_ ( .A1(_12624_ ), .A2(_12786_ ), .B1(\ifu.io_out_bits_pc [23] ), .B2(_12645_ ), .ZN(_12787_ ) );
AOI21_X1 _19696_ ( .A(fanout_net_23 ), .B1(_12784_ ), .B2(_12787_ ), .ZN(_00289_ ) );
XNOR2_X1 _19697_ ( .A(_12771_ ), .B(_09558_ ), .ZN(_12788_ ) );
AND3_X1 _19698_ ( .A1(_12733_ ), .A2(_11899_ ), .A3(_12788_ ), .ZN(_12789_ ) );
INV_X1 _19699_ ( .A(_09560_ ), .ZN(\ifu.io_out_bits_pc [22] ) );
AOI21_X1 _19700_ ( .A(_12789_ ), .B1(\ifu.io_out_bits_pc [22] ), .B2(_12646_ ), .ZN(_12790_ ) );
INV_X1 _19701_ ( .A(_12585_ ), .ZN(_12791_ ) );
OR2_X1 _19702_ ( .A1(_12583_ ), .A2(_12584_ ), .ZN(_12792_ ) );
NAND4_X1 _19703_ ( .A1(_idu_io_in_bits_T ), .A2(_12648_ ), .A3(_12791_ ), .A4(_12792_ ), .ZN(_12793_ ) );
AOI21_X1 _19704_ ( .A(fanout_net_23 ), .B1(_12790_ ), .B2(_12793_ ), .ZN(_00290_ ) );
NAND3_X1 _19705_ ( .A1(_12638_ ), .A2(_12641_ ), .A3(_12719_ ), .ZN(_12794_ ) );
NOR2_X1 _19706_ ( .A1(_12794_ ), .A2(_10055_ ), .ZN(_12795_ ) );
XNOR2_X1 _19707_ ( .A(_12795_ ), .B(_09606_ ), .ZN(_12796_ ) );
AND3_X1 _19708_ ( .A1(_12733_ ), .A2(_11899_ ), .A3(_12796_ ), .ZN(_12797_ ) );
INV_X1 _19709_ ( .A(_09608_ ), .ZN(\ifu.io_out_bits_pc [21] ) );
AOI21_X1 _19710_ ( .A(_12797_ ), .B1(\ifu.io_out_bits_pc [21] ), .B2(_12646_ ), .ZN(_12798_ ) );
INV_X1 _19711_ ( .A(_12583_ ), .ZN(_12799_ ) );
OR2_X1 _19712_ ( .A1(_12581_ ), .A2(_12582_ ), .ZN(_12800_ ) );
NAND4_X1 _19713_ ( .A1(_idu_io_in_bits_T ), .A2(_12648_ ), .A3(_12799_ ), .A4(_12800_ ), .ZN(_12801_ ) );
AOI21_X1 _19714_ ( .A(fanout_net_23 ), .B1(_12798_ ), .B2(_12801_ ), .ZN(_00291_ ) );
XNOR2_X1 _19715_ ( .A(_12794_ ), .B(\ifu.pc [20] ), .ZN(_12802_ ) );
AND3_X1 _19716_ ( .A1(_10833_ ), .A2(_11899_ ), .A3(_12802_ ), .ZN(_12803_ ) );
AND2_X1 _19717_ ( .A1(_10052_ ), .A2(_10053_ ), .ZN(_12804_ ) );
INV_X1 _19718_ ( .A(_12804_ ), .ZN(\ifu.io_out_bits_pc [20] ) );
AOI21_X1 _19719_ ( .A(_12803_ ), .B1(\ifu.io_out_bits_pc [20] ), .B2(_12646_ ), .ZN(_12805_ ) );
INV_X1 _19720_ ( .A(_12581_ ), .ZN(_12806_ ) );
OR2_X1 _19721_ ( .A1(_12579_ ), .A2(_12580_ ), .ZN(_12807_ ) );
NAND4_X1 _19722_ ( .A1(_idu_io_in_bits_T ), .A2(_12648_ ), .A3(_12806_ ), .A4(_12807_ ), .ZN(_12808_ ) );
AOI21_X1 _19723_ ( .A(fanout_net_23 ), .B1(_12805_ ), .B2(_12808_ ), .ZN(_00292_ ) );
INV_X1 _19724_ ( .A(_11974_ ), .ZN(\ifu.io_out_bits_pc [29] ) );
NOR2_X1 _19725_ ( .A1(_12717_ ), .A2(_12720_ ), .ZN(_12809_ ) );
AND2_X1 _19726_ ( .A1(\ifu.pc [27] ), .A2(\ifu.pc [26] ), .ZN(_12810_ ) );
NAND3_X1 _19727_ ( .A1(_12809_ ), .A2(\ifu.pc [28] ), .A3(_12810_ ), .ZN(_12811_ ) );
XNOR2_X1 _19728_ ( .A(_12811_ ), .B(\ifu.pc [29] ), .ZN(_12812_ ) );
AOI221_X1 _19729_ ( .A(fanout_net_23 ), .B1(_12645_ ), .B2(\ifu.io_out_bits_pc [29] ), .C1(_12624_ ), .C2(_12812_ ), .ZN(_12813_ ) );
XNOR2_X1 _19730_ ( .A(_12596_ ), .B(_12600_ ), .ZN(_12814_ ) );
NAND2_X1 _19731_ ( .A1(_12814_ ), .A2(_12550_ ), .ZN(_12815_ ) );
NAND2_X1 _19732_ ( .A1(_12813_ ), .A2(_12815_ ), .ZN(_00293_ ) );
INV_X1 _19733_ ( .A(_12596_ ), .ZN(_12816_ ) );
OR2_X1 _19734_ ( .A1(_12724_ ), .A2(_12594_ ), .ZN(_12817_ ) );
NAND3_X1 _19735_ ( .A1(_12550_ ), .A2(_12816_ ), .A3(_12817_ ), .ZN(_12818_ ) );
AOI21_X1 _19736_ ( .A(fanout_net_23 ), .B1(_09399_ ), .B2(_09403_ ), .ZN(_12819_ ) );
INV_X1 _19737_ ( .A(_12631_ ), .ZN(\ifu.pc_$_SDFFE_PP0P__Q_E ) );
NAND2_X1 _19738_ ( .A1(_12809_ ), .A2(_12810_ ), .ZN(_12820_ ) );
XNOR2_X1 _19739_ ( .A(_12820_ ), .B(_09400_ ), .ZN(_12821_ ) );
OAI221_X1 _19740_ ( .A(_12818_ ), .B1(_00230_ ), .B2(_12819_ ), .C1(\ifu.pc_$_SDFFE_PP0P__Q_E ), .C2(_12821_ ), .ZN(_00294_ ) );
NAND2_X1 _19741_ ( .A1(\ifu.start [0] ), .A2(\ifu.start [1] ), .ZN(_12822_ ) );
NAND3_X1 _19742_ ( .A1(\ifu._start_T ), .A2(\ifu.ren_REG_$_DFF_P__Q_D_$_NAND__Y_B ), .A3(_12822_ ), .ZN(_00295_ ) );
BUF_X2 _19743_ ( .A(_11358_ ), .Z(\exu._io_out_bits_wdata_T_1 [4] ) );
BUF_X4 _19744_ ( .A(_11397_ ), .Z(_12823_ ) );
MUX2_X1 _19745_ ( .A(\exu._GEN_0 [15] ), .B(\exu._GEN_0 [7] ), .S(_12823_ ), .Z(_12824_ ) );
INV_X1 _19746_ ( .A(_11358_ ), .ZN(_12825_ ) );
AND2_X1 _19747_ ( .A1(_12824_ ), .A2(_12825_ ), .ZN(_00296_ ) );
MUX2_X1 _19748_ ( .A(\exu._GEN_0 [14] ), .B(\exu._GEN_0 [6] ), .S(_12823_ ), .Z(_12826_ ) );
AND2_X1 _19749_ ( .A1(_12826_ ), .A2(_12825_ ), .ZN(_00297_ ) );
INV_X1 _19750_ ( .A(_11397_ ), .ZN(_12827_ ) );
BUF_X2 _19751_ ( .A(_12827_ ), .Z(_12828_ ) );
AND4_X1 _19752_ ( .A1(\exu._GEN_0 [5] ), .A2(_11356_ ), .A3(_11357_ ), .A4(_12828_ ), .ZN(_00298_ ) );
INV_X1 _19753_ ( .A(_11396_ ), .ZN(_12829_ ) );
AOI21_X1 _19754_ ( .A(\exu.io_out_bits_wdata_$_MUX__Y_11_B_$_ANDNOT__Y_B ), .B1(_09054_ ), .B2(_12829_ ), .ZN(_12830_ ) );
AND3_X1 _19755_ ( .A1(_12830_ ), .A2(_11356_ ), .A3(_11357_ ), .ZN(_00299_ ) );
INV_X1 _19756_ ( .A(\exu.io_out_bits_wdata_$_MUX__Y_12_B_$_ANDNOT__Y_B ), .ZN(_12831_ ) );
AND4_X1 _19757_ ( .A1(_12831_ ), .A2(_11356_ ), .A3(_11357_ ), .A4(_12828_ ), .ZN(_00300_ ) );
INV_X1 _19758_ ( .A(\exu.io_out_bits_wdata_$_MUX__Y_13_B_$_ANDNOT__Y_B ), .ZN(_12832_ ) );
AND4_X1 _19759_ ( .A1(_12832_ ), .A2(_11356_ ), .A3(_11357_ ), .A4(_12828_ ), .ZN(_00301_ ) );
INV_X1 _19760_ ( .A(\exu.io_out_bits_wdata_$_MUX__Y_14_B_$_ANDNOT__Y_B ), .ZN(_12833_ ) );
AND4_X1 _19761_ ( .A1(_12833_ ), .A2(_11356_ ), .A3(_11357_ ), .A4(_12828_ ), .ZN(_00302_ ) );
AND4_X1 _19762_ ( .A1(\exu._GEN_0 [0] ), .A2(_11356_ ), .A3(_11357_ ), .A4(_12828_ ), .ZN(_00303_ ) );
MUX2_X1 _19763_ ( .A(\exu._GEN_0 [13] ), .B(\exu._GEN_0 [5] ), .S(_12823_ ), .Z(_12834_ ) );
AND2_X1 _19764_ ( .A1(_12834_ ), .A2(_12825_ ), .ZN(_00304_ ) );
MUX2_X1 _19765_ ( .A(\exu._GEN_0 [12] ), .B(\exu._GEN_0 [4] ), .S(_11397_ ), .Z(_12835_ ) );
AND2_X1 _19766_ ( .A1(_12835_ ), .A2(_12825_ ), .ZN(_00305_ ) );
MUX2_X1 _19767_ ( .A(\exu._GEN_0 [11] ), .B(\exu._GEN_0 [3] ), .S(_11397_ ), .Z(_12836_ ) );
AND2_X1 _19768_ ( .A1(_12836_ ), .A2(_12825_ ), .ZN(_00306_ ) );
MUX2_X1 _19769_ ( .A(\exu._GEN_0 [10] ), .B(\exu._GEN_0 [2] ), .S(_11397_ ), .Z(_12837_ ) );
AND2_X1 _19770_ ( .A1(_12837_ ), .A2(_12825_ ), .ZN(_00307_ ) );
MUX2_X1 _19771_ ( .A(\exu._GEN_0 [9] ), .B(\exu._GEN_0 [1] ), .S(_11397_ ), .Z(_12838_ ) );
AND2_X1 _19772_ ( .A1(_12838_ ), .A2(_12825_ ), .ZN(_00308_ ) );
MUX2_X1 _19773_ ( .A(\exu._GEN_0 [8] ), .B(\exu._GEN_0 [0] ), .S(_11397_ ), .Z(_12839_ ) );
AND2_X1 _19774_ ( .A1(_12839_ ), .A2(_12825_ ), .ZN(_00309_ ) );
AOI21_X1 _19775_ ( .A(_08833_ ), .B1(_09054_ ), .B2(_12829_ ), .ZN(_12840_ ) );
AND3_X1 _19776_ ( .A1(_12840_ ), .A2(_11356_ ), .A3(_11357_ ), .ZN(_00310_ ) );
INV_X1 _19777_ ( .A(\exu._GEN_0 [6] ), .ZN(_12841_ ) );
AOI21_X1 _19778_ ( .A(_12841_ ), .B1(_09054_ ), .B2(_12829_ ), .ZN(_12842_ ) );
AND3_X1 _19779_ ( .A1(_12842_ ), .A2(_11356_ ), .A3(_11357_ ), .ZN(_00311_ ) );
INV_X1 _19780_ ( .A(\exu.io_in_valid ), .ZN(_12843_ ) );
AOI21_X1 _19781_ ( .A(_10991_ ), .B1(_12843_ ), .B2(_10827_ ), .ZN(_lsu_io_in_bits_T ) );
AOI211_X1 _19782_ ( .A(fanout_net_23 ), .B(_10991_ ), .C1(_12843_ ), .C2(_10827_ ), .ZN(_00312_ ) );
AND2_X2 _19783_ ( .A1(\wbu.io_in_bits_wen_csr ), .A2(\ifu.io_valid ), .ZN(_12844_ ) );
INV_X1 _19784_ ( .A(_12844_ ), .ZN(_12845_ ) );
NOR2_X1 _19785_ ( .A1(_12845_ ), .A2(\wbu.io_in_bits_csr_wdata [31] ), .ZN(_12846_ ) );
INV_X1 _19786_ ( .A(fanout_net_28 ), .ZN(_12847_ ) );
AND2_X2 _19787_ ( .A1(fanout_net_28 ), .A2(\wbu.io_in_bits_csr_waddr [0] ), .ZN(_12848_ ) );
AOI221_X4 _19788_ ( .A(_12844_ ), .B1(\wbu._GEN_135 [31] ), .B2(_12847_ ), .C1(\wbu.csr_3 [31] ), .C2(_12848_ ), .ZN(_12849_ ) );
AND3_X1 _19789_ ( .A1(_08577_ ), .A2(\wbu.csr_2 [31] ), .A3(fanout_net_28 ), .ZN(_12850_ ) );
INV_X1 _19790_ ( .A(_12850_ ), .ZN(_12851_ ) );
AOI211_X1 _19791_ ( .A(fanout_net_23 ), .B(_12846_ ), .C1(_12849_ ), .C2(_12851_ ), .ZN(_00313_ ) );
BUF_X4 _19792_ ( .A(_12845_ ), .Z(_12852_ ) );
NOR2_X1 _19793_ ( .A1(_12852_ ), .A2(\wbu.io_in_bits_csr_wdata [30] ), .ZN(_12853_ ) );
BUF_X4 _19794_ ( .A(_12844_ ), .Z(_12854_ ) );
BUF_X4 _19795_ ( .A(_12847_ ), .Z(_12855_ ) );
BUF_X2 _19796_ ( .A(_12848_ ), .Z(wbu_io_in_bits_csr_waddr_$_AND__A_Y ) );
AOI221_X4 _19797_ ( .A(_12854_ ), .B1(\wbu._GEN_135 [30] ), .B2(_12855_ ), .C1(\wbu.csr_3 [30] ), .C2(wbu_io_in_bits_csr_waddr_$_AND__A_Y ), .ZN(_12856_ ) );
NAND3_X1 _19798_ ( .A1(_08578_ ), .A2(\wbu.csr_2 [30] ), .A3(fanout_net_28 ), .ZN(_12857_ ) );
AOI211_X1 _19799_ ( .A(fanout_net_23 ), .B(_12853_ ), .C1(_12856_ ), .C2(_12857_ ), .ZN(_00314_ ) );
NOR2_X1 _19800_ ( .A1(_12852_ ), .A2(\wbu.io_in_bits_csr_wdata [21] ), .ZN(_12858_ ) );
AOI221_X4 _19801_ ( .A(_12854_ ), .B1(\wbu._GEN_135 [21] ), .B2(_12855_ ), .C1(\wbu.csr_3 [21] ), .C2(wbu_io_in_bits_csr_waddr_$_AND__A_Y ), .ZN(_12859_ ) );
NAND3_X1 _19802_ ( .A1(_08578_ ), .A2(\wbu.csr_2 [21] ), .A3(fanout_net_28 ), .ZN(_12860_ ) );
AOI211_X1 _19803_ ( .A(fanout_net_23 ), .B(_12858_ ), .C1(_12859_ ), .C2(_12860_ ), .ZN(_00315_ ) );
NOR2_X1 _19804_ ( .A1(_12852_ ), .A2(\wbu.io_in_bits_csr_wdata [20] ), .ZN(_12861_ ) );
AOI221_X4 _19805_ ( .A(_12854_ ), .B1(\wbu._GEN_135 [20] ), .B2(_12855_ ), .C1(\wbu.csr_3 [20] ), .C2(wbu_io_in_bits_csr_waddr_$_AND__A_Y ), .ZN(_12862_ ) );
NAND3_X1 _19806_ ( .A1(_08578_ ), .A2(\wbu.csr_2 [20] ), .A3(fanout_net_28 ), .ZN(_12863_ ) );
AOI211_X1 _19807_ ( .A(fanout_net_23 ), .B(_12861_ ), .C1(_12862_ ), .C2(_12863_ ), .ZN(_00316_ ) );
NOR2_X1 _19808_ ( .A1(_12852_ ), .A2(\wbu.io_in_bits_csr_wdata [19] ), .ZN(_12864_ ) );
AOI221_X4 _19809_ ( .A(_12854_ ), .B1(\wbu._GEN_135 [19] ), .B2(_12855_ ), .C1(\wbu.csr_3 [19] ), .C2(wbu_io_in_bits_csr_waddr_$_AND__A_Y ), .ZN(_12865_ ) );
NAND3_X1 _19810_ ( .A1(_08578_ ), .A2(\wbu.csr_2 [19] ), .A3(fanout_net_28 ), .ZN(_12866_ ) );
AOI211_X1 _19811_ ( .A(fanout_net_23 ), .B(_12864_ ), .C1(_12865_ ), .C2(_12866_ ), .ZN(_00317_ ) );
NOR2_X1 _19812_ ( .A1(_12852_ ), .A2(\wbu.io_in_bits_csr_wdata [18] ), .ZN(_12867_ ) );
AOI221_X4 _19813_ ( .A(_12854_ ), .B1(\wbu._GEN_135 [18] ), .B2(_12855_ ), .C1(\wbu.csr_3 [18] ), .C2(wbu_io_in_bits_csr_waddr_$_AND__A_Y ), .ZN(_12868_ ) );
NAND3_X1 _19814_ ( .A1(_08578_ ), .A2(\wbu.csr_2 [18] ), .A3(fanout_net_28 ), .ZN(_12869_ ) );
AOI211_X1 _19815_ ( .A(fanout_net_23 ), .B(_12867_ ), .C1(_12868_ ), .C2(_12869_ ), .ZN(_00318_ ) );
NOR2_X1 _19816_ ( .A1(_12852_ ), .A2(\wbu.io_in_bits_csr_wdata [17] ), .ZN(_12870_ ) );
AOI221_X4 _19817_ ( .A(_12854_ ), .B1(\wbu._GEN_135 [17] ), .B2(_12855_ ), .C1(\wbu.csr_3 [17] ), .C2(wbu_io_in_bits_csr_waddr_$_AND__A_Y ), .ZN(_12871_ ) );
NAND3_X1 _19818_ ( .A1(_08578_ ), .A2(\wbu.csr_2 [17] ), .A3(fanout_net_28 ), .ZN(_12872_ ) );
AOI211_X1 _19819_ ( .A(fanout_net_23 ), .B(_12870_ ), .C1(_12871_ ), .C2(_12872_ ), .ZN(_00319_ ) );
NOR2_X1 _19820_ ( .A1(_12852_ ), .A2(\wbu.io_in_bits_csr_wdata [16] ), .ZN(_12873_ ) );
AOI221_X4 _19821_ ( .A(_12854_ ), .B1(\wbu._GEN_135 [16] ), .B2(_12855_ ), .C1(\wbu.csr_3 [16] ), .C2(wbu_io_in_bits_csr_waddr_$_AND__A_Y ), .ZN(_12874_ ) );
NAND3_X1 _19822_ ( .A1(_08578_ ), .A2(\wbu.csr_2 [16] ), .A3(fanout_net_28 ), .ZN(_12875_ ) );
AOI211_X1 _19823_ ( .A(fanout_net_23 ), .B(_12873_ ), .C1(_12874_ ), .C2(_12875_ ), .ZN(_00320_ ) );
NOR2_X1 _19824_ ( .A1(_12852_ ), .A2(\wbu.io_in_bits_csr_wdata [15] ), .ZN(_12876_ ) );
AOI221_X4 _19825_ ( .A(_12854_ ), .B1(\wbu._GEN_135 [15] ), .B2(_12855_ ), .C1(\wbu.csr_3 [15] ), .C2(wbu_io_in_bits_csr_waddr_$_AND__A_Y ), .ZN(_12877_ ) );
NAND3_X1 _19826_ ( .A1(_08578_ ), .A2(\wbu.csr_2 [15] ), .A3(fanout_net_28 ), .ZN(_12878_ ) );
AOI211_X1 _19827_ ( .A(fanout_net_23 ), .B(_12876_ ), .C1(_12877_ ), .C2(_12878_ ), .ZN(_00321_ ) );
NOR2_X1 _19828_ ( .A1(_12852_ ), .A2(\wbu.io_in_bits_csr_wdata [14] ), .ZN(_12879_ ) );
AOI221_X4 _19829_ ( .A(_12854_ ), .B1(\wbu._GEN_135 [14] ), .B2(_12855_ ), .C1(\wbu.csr_3 [14] ), .C2(wbu_io_in_bits_csr_waddr_$_AND__A_Y ), .ZN(_12880_ ) );
NAND3_X1 _19830_ ( .A1(_08578_ ), .A2(\wbu.csr_2 [14] ), .A3(fanout_net_28 ), .ZN(_12881_ ) );
AOI211_X1 _19831_ ( .A(fanout_net_23 ), .B(_12879_ ), .C1(_12880_ ), .C2(_12881_ ), .ZN(_00322_ ) );
NOR2_X1 _19832_ ( .A1(_12852_ ), .A2(\wbu.io_in_bits_csr_wdata [13] ), .ZN(_12882_ ) );
BUF_X4 _19833_ ( .A(_12847_ ), .Z(_12883_ ) );
BUF_X4 _19834_ ( .A(_12848_ ), .Z(_12884_ ) );
AOI221_X4 _19835_ ( .A(_12854_ ), .B1(\wbu._GEN_135 [13] ), .B2(_12883_ ), .C1(\wbu.csr_3 [13] ), .C2(_12884_ ), .ZN(_12885_ ) );
BUF_X4 _19836_ ( .A(_08577_ ), .Z(_12886_ ) );
NAND3_X1 _19837_ ( .A1(_12886_ ), .A2(\wbu.csr_2 [13] ), .A3(fanout_net_28 ), .ZN(_12887_ ) );
AOI211_X1 _19838_ ( .A(fanout_net_23 ), .B(_12882_ ), .C1(_12885_ ), .C2(_12887_ ), .ZN(_00323_ ) );
BUF_X4 _19839_ ( .A(_12845_ ), .Z(_12888_ ) );
NOR2_X1 _19840_ ( .A1(_12888_ ), .A2(\wbu.io_in_bits_csr_wdata [12] ), .ZN(_12889_ ) );
BUF_X4 _19841_ ( .A(_12844_ ), .Z(_12890_ ) );
AOI221_X4 _19842_ ( .A(_12890_ ), .B1(\wbu._GEN_135 [12] ), .B2(_12883_ ), .C1(\wbu.csr_3 [12] ), .C2(_12884_ ), .ZN(_12891_ ) );
NAND3_X1 _19843_ ( .A1(_12886_ ), .A2(\wbu.csr_2 [12] ), .A3(fanout_net_28 ), .ZN(_12892_ ) );
AOI211_X1 _19844_ ( .A(fanout_net_23 ), .B(_12889_ ), .C1(_12891_ ), .C2(_12892_ ), .ZN(_00324_ ) );
NOR2_X1 _19845_ ( .A1(_12888_ ), .A2(\wbu.io_in_bits_csr_wdata [29] ), .ZN(_12893_ ) );
AOI221_X4 _19846_ ( .A(_12890_ ), .B1(\wbu._GEN_135 [29] ), .B2(_12883_ ), .C1(\wbu.csr_3 [29] ), .C2(_12884_ ), .ZN(_12894_ ) );
NAND3_X1 _19847_ ( .A1(_12886_ ), .A2(\wbu.csr_2 [29] ), .A3(fanout_net_28 ), .ZN(_12895_ ) );
AOI211_X1 _19848_ ( .A(fanout_net_23 ), .B(_12893_ ), .C1(_12894_ ), .C2(_12895_ ), .ZN(_00325_ ) );
NOR2_X1 _19849_ ( .A1(_12888_ ), .A2(\wbu.io_in_bits_csr_wdata [11] ), .ZN(_12896_ ) );
AOI221_X4 _19850_ ( .A(_12890_ ), .B1(\wbu._GEN_135 [11] ), .B2(_12883_ ), .C1(\wbu.csr_3 [11] ), .C2(_12884_ ), .ZN(_12897_ ) );
NAND3_X1 _19851_ ( .A1(_12886_ ), .A2(\wbu.csr_2 [11] ), .A3(fanout_net_28 ), .ZN(_12898_ ) );
AOI211_X1 _19852_ ( .A(fanout_net_23 ), .B(_12896_ ), .C1(_12897_ ), .C2(_12898_ ), .ZN(_00326_ ) );
NOR2_X1 _19853_ ( .A1(_12888_ ), .A2(\wbu.io_in_bits_csr_wdata [10] ), .ZN(_12899_ ) );
AOI221_X4 _19854_ ( .A(_12890_ ), .B1(\wbu._GEN_135 [10] ), .B2(_12883_ ), .C1(\wbu.csr_3 [10] ), .C2(_12884_ ), .ZN(_12900_ ) );
NAND3_X1 _19855_ ( .A1(_12886_ ), .A2(\wbu.csr_2 [10] ), .A3(fanout_net_28 ), .ZN(_12901_ ) );
AOI211_X1 _19856_ ( .A(fanout_net_23 ), .B(_12899_ ), .C1(_12900_ ), .C2(_12901_ ), .ZN(_00327_ ) );
NOR2_X1 _19857_ ( .A1(_12888_ ), .A2(\wbu.io_in_bits_csr_wdata [9] ), .ZN(_12902_ ) );
AOI221_X4 _19858_ ( .A(_12890_ ), .B1(\wbu._GEN_135 [9] ), .B2(_12883_ ), .C1(\wbu.csr_3 [9] ), .C2(_12884_ ), .ZN(_12903_ ) );
NAND3_X1 _19859_ ( .A1(_12886_ ), .A2(\wbu.csr_2 [9] ), .A3(fanout_net_28 ), .ZN(_12904_ ) );
AOI211_X1 _19860_ ( .A(fanout_net_23 ), .B(_12902_ ), .C1(_12903_ ), .C2(_12904_ ), .ZN(_00328_ ) );
NOR2_X1 _19861_ ( .A1(_12888_ ), .A2(\wbu.io_in_bits_csr_wdata [8] ), .ZN(_12905_ ) );
AOI221_X4 _19862_ ( .A(_12890_ ), .B1(\wbu._GEN_135 [8] ), .B2(_12883_ ), .C1(\wbu.csr_3 [8] ), .C2(_12884_ ), .ZN(_12906_ ) );
NAND3_X1 _19863_ ( .A1(_12886_ ), .A2(\wbu.csr_2 [8] ), .A3(fanout_net_28 ), .ZN(_12907_ ) );
AOI211_X1 _19864_ ( .A(fanout_net_23 ), .B(_12905_ ), .C1(_12906_ ), .C2(_12907_ ), .ZN(_00329_ ) );
NOR2_X1 _19865_ ( .A1(_12888_ ), .A2(\wbu.io_in_bits_csr_wdata [7] ), .ZN(_12908_ ) );
AOI221_X4 _19866_ ( .A(_12890_ ), .B1(\wbu._GEN_135 [7] ), .B2(_12883_ ), .C1(\wbu.csr_3 [7] ), .C2(_12884_ ), .ZN(_12909_ ) );
NAND3_X1 _19867_ ( .A1(_12886_ ), .A2(\wbu.csr_2 [7] ), .A3(fanout_net_28 ), .ZN(_12910_ ) );
AOI211_X1 _19868_ ( .A(fanout_net_23 ), .B(_12908_ ), .C1(_12909_ ), .C2(_12910_ ), .ZN(_00330_ ) );
NOR2_X1 _19869_ ( .A1(_12888_ ), .A2(\wbu.io_in_bits_csr_wdata [6] ), .ZN(_12911_ ) );
AOI221_X4 _19870_ ( .A(_12890_ ), .B1(\wbu._GEN_135 [6] ), .B2(_12883_ ), .C1(\wbu.csr_3 [6] ), .C2(_12884_ ), .ZN(_12912_ ) );
NAND3_X1 _19871_ ( .A1(_12886_ ), .A2(\wbu.csr_2 [6] ), .A3(fanout_net_28 ), .ZN(_12913_ ) );
AOI211_X1 _19872_ ( .A(fanout_net_23 ), .B(_12911_ ), .C1(_12912_ ), .C2(_12913_ ), .ZN(_00331_ ) );
NOR2_X1 _19873_ ( .A1(_12888_ ), .A2(\wbu.io_in_bits_csr_wdata [5] ), .ZN(_12914_ ) );
AOI221_X4 _19874_ ( .A(_12890_ ), .B1(\wbu._GEN_135 [5] ), .B2(_12883_ ), .C1(\wbu.csr_3 [5] ), .C2(_12884_ ), .ZN(_12915_ ) );
NAND3_X1 _19875_ ( .A1(_12886_ ), .A2(\wbu.csr_2 [5] ), .A3(fanout_net_28 ), .ZN(_12916_ ) );
AOI211_X1 _19876_ ( .A(fanout_net_23 ), .B(_12914_ ), .C1(_12915_ ), .C2(_12916_ ), .ZN(_00332_ ) );
NOR2_X1 _19877_ ( .A1(_12888_ ), .A2(\wbu.io_in_bits_csr_wdata [4] ), .ZN(_12917_ ) );
BUF_X4 _19878_ ( .A(_12847_ ), .Z(_12918_ ) );
BUF_X4 _19879_ ( .A(_12848_ ), .Z(_12919_ ) );
AOI221_X4 _19880_ ( .A(_12890_ ), .B1(\wbu._GEN_135 [4] ), .B2(_12918_ ), .C1(\wbu.csr_3 [4] ), .C2(_12919_ ), .ZN(_12920_ ) );
BUF_X4 _19881_ ( .A(_08577_ ), .Z(_12921_ ) );
NAND3_X1 _19882_ ( .A1(_12921_ ), .A2(\wbu.csr_2 [4] ), .A3(fanout_net_28 ), .ZN(_12922_ ) );
AOI211_X1 _19883_ ( .A(fanout_net_23 ), .B(_12917_ ), .C1(_12920_ ), .C2(_12922_ ), .ZN(_00333_ ) );
BUF_X4 _19884_ ( .A(_12845_ ), .Z(_12923_ ) );
NOR2_X1 _19885_ ( .A1(_12923_ ), .A2(\wbu.io_in_bits_csr_wdata [3] ), .ZN(_12924_ ) );
BUF_X4 _19886_ ( .A(_12844_ ), .Z(_12925_ ) );
AOI221_X4 _19887_ ( .A(_12925_ ), .B1(\wbu._GEN_135 [3] ), .B2(_12918_ ), .C1(\wbu.csr_3 [3] ), .C2(_12919_ ), .ZN(_12926_ ) );
NAND3_X1 _19888_ ( .A1(_12921_ ), .A2(\wbu.csr_2 [3] ), .A3(fanout_net_28 ), .ZN(_12927_ ) );
AOI211_X1 _19889_ ( .A(fanout_net_23 ), .B(_12924_ ), .C1(_12926_ ), .C2(_12927_ ), .ZN(_00334_ ) );
NOR2_X1 _19890_ ( .A1(_12923_ ), .A2(\wbu.io_in_bits_csr_wdata [2] ), .ZN(_12928_ ) );
AOI221_X4 _19891_ ( .A(_12925_ ), .B1(\wbu._GEN_135 [2] ), .B2(_12918_ ), .C1(\wbu.csr_3 [2] ), .C2(_12919_ ), .ZN(_12929_ ) );
NAND3_X1 _19892_ ( .A1(_12921_ ), .A2(\wbu.csr_2 [2] ), .A3(fanout_net_28 ), .ZN(_12930_ ) );
AOI211_X1 _19893_ ( .A(fanout_net_23 ), .B(_12928_ ), .C1(_12929_ ), .C2(_12930_ ), .ZN(_00335_ ) );
NOR2_X1 _19894_ ( .A1(_12923_ ), .A2(\wbu.io_in_bits_csr_wdata [28] ), .ZN(_12931_ ) );
AOI221_X4 _19895_ ( .A(_12925_ ), .B1(\wbu._GEN_135 [28] ), .B2(_12918_ ), .C1(\wbu.csr_3 [28] ), .C2(_12919_ ), .ZN(_12932_ ) );
NAND3_X1 _19896_ ( .A1(_12921_ ), .A2(\wbu.csr_2 [28] ), .A3(fanout_net_28 ), .ZN(_12933_ ) );
AOI211_X1 _19897_ ( .A(fanout_net_24 ), .B(_12931_ ), .C1(_12932_ ), .C2(_12933_ ), .ZN(_00336_ ) );
NOR2_X1 _19898_ ( .A1(_12923_ ), .A2(\wbu.io_in_bits_csr_wdata [1] ), .ZN(_12934_ ) );
AOI221_X4 _19899_ ( .A(_12925_ ), .B1(\wbu._GEN_135 [1] ), .B2(_12918_ ), .C1(\wbu.csr_3 [1] ), .C2(_12919_ ), .ZN(_12935_ ) );
NAND3_X1 _19900_ ( .A1(_12921_ ), .A2(\wbu.csr_2 [1] ), .A3(fanout_net_28 ), .ZN(_12936_ ) );
AOI211_X1 _19901_ ( .A(fanout_net_24 ), .B(_12934_ ), .C1(_12935_ ), .C2(_12936_ ), .ZN(_00337_ ) );
NOR2_X1 _19902_ ( .A1(_12923_ ), .A2(\wbu.io_in_bits_csr_wdata [0] ), .ZN(_12937_ ) );
AOI221_X4 _19903_ ( .A(_12925_ ), .B1(\wbu._GEN_135 [0] ), .B2(_12918_ ), .C1(\wbu.csr_3 [0] ), .C2(_12919_ ), .ZN(_12938_ ) );
NAND3_X1 _19904_ ( .A1(_12921_ ), .A2(\wbu.csr_2 [0] ), .A3(fanout_net_28 ), .ZN(_12939_ ) );
AOI211_X1 _19905_ ( .A(fanout_net_24 ), .B(_12937_ ), .C1(_12938_ ), .C2(_12939_ ), .ZN(_00338_ ) );
NOR2_X1 _19906_ ( .A1(_12923_ ), .A2(\wbu.io_in_bits_csr_wdata [27] ), .ZN(_12940_ ) );
AOI221_X4 _19907_ ( .A(_12925_ ), .B1(\wbu._GEN_135 [27] ), .B2(_12918_ ), .C1(\wbu.csr_3 [27] ), .C2(_12919_ ), .ZN(_12941_ ) );
NAND3_X1 _19908_ ( .A1(_12921_ ), .A2(\wbu.csr_2 [27] ), .A3(fanout_net_28 ), .ZN(_12942_ ) );
AOI211_X1 _19909_ ( .A(fanout_net_24 ), .B(_12940_ ), .C1(_12941_ ), .C2(_12942_ ), .ZN(_00339_ ) );
NOR2_X1 _19910_ ( .A1(_12923_ ), .A2(\wbu.io_in_bits_csr_wdata [26] ), .ZN(_12943_ ) );
AOI221_X4 _19911_ ( .A(_12925_ ), .B1(\wbu._GEN_135 [26] ), .B2(_12918_ ), .C1(\wbu.csr_3 [26] ), .C2(_12919_ ), .ZN(_12944_ ) );
NAND3_X1 _19912_ ( .A1(_12921_ ), .A2(\wbu.csr_2 [26] ), .A3(\wbu.io_in_bits_csr_waddr [1] ), .ZN(_12945_ ) );
AOI211_X1 _19913_ ( .A(fanout_net_24 ), .B(_12943_ ), .C1(_12944_ ), .C2(_12945_ ), .ZN(_00340_ ) );
NOR2_X1 _19914_ ( .A1(_12923_ ), .A2(\wbu.io_in_bits_csr_wdata [25] ), .ZN(_12946_ ) );
AOI221_X4 _19915_ ( .A(_12925_ ), .B1(\wbu._GEN_135 [25] ), .B2(_12918_ ), .C1(\wbu.csr_3 [25] ), .C2(_12919_ ), .ZN(_12947_ ) );
NAND3_X1 _19916_ ( .A1(_12921_ ), .A2(\wbu.csr_2 [25] ), .A3(\wbu.io_in_bits_csr_waddr [1] ), .ZN(_12948_ ) );
AOI211_X1 _19917_ ( .A(fanout_net_24 ), .B(_12946_ ), .C1(_12947_ ), .C2(_12948_ ), .ZN(_00341_ ) );
NOR2_X1 _19918_ ( .A1(_12923_ ), .A2(\wbu.io_in_bits_csr_wdata [24] ), .ZN(_12949_ ) );
AOI221_X4 _19919_ ( .A(_12925_ ), .B1(\wbu._GEN_135 [24] ), .B2(_12918_ ), .C1(\wbu.csr_3 [24] ), .C2(_12919_ ), .ZN(_12950_ ) );
NAND3_X1 _19920_ ( .A1(_12921_ ), .A2(\wbu.csr_2 [24] ), .A3(\wbu.io_in_bits_csr_waddr [1] ), .ZN(_12951_ ) );
AOI211_X1 _19921_ ( .A(fanout_net_24 ), .B(_12949_ ), .C1(_12950_ ), .C2(_12951_ ), .ZN(_00342_ ) );
NOR2_X1 _19922_ ( .A1(_12923_ ), .A2(\wbu.io_in_bits_csr_wdata [23] ), .ZN(_12952_ ) );
AOI221_X4 _19923_ ( .A(_12925_ ), .B1(\wbu._GEN_135 [23] ), .B2(_12847_ ), .C1(\wbu.csr_3 [23] ), .C2(_12848_ ), .ZN(_12953_ ) );
NAND3_X1 _19924_ ( .A1(_08577_ ), .A2(\wbu.csr_2 [23] ), .A3(\wbu.io_in_bits_csr_waddr [1] ), .ZN(_12954_ ) );
AOI211_X1 _19925_ ( .A(fanout_net_24 ), .B(_12952_ ), .C1(_12953_ ), .C2(_12954_ ), .ZN(_00343_ ) );
NOR2_X1 _19926_ ( .A1(_12845_ ), .A2(\wbu.io_in_bits_csr_wdata [22] ), .ZN(_12955_ ) );
AOI221_X4 _19927_ ( .A(_12844_ ), .B1(\wbu._GEN_135 [22] ), .B2(_12847_ ), .C1(\wbu.csr_3 [22] ), .C2(_12848_ ), .ZN(_12956_ ) );
NAND3_X1 _19928_ ( .A1(_08577_ ), .A2(\wbu.csr_2 [22] ), .A3(\wbu.io_in_bits_csr_waddr [1] ), .ZN(_12957_ ) );
AOI211_X1 _19929_ ( .A(fanout_net_24 ), .B(_12955_ ), .C1(_12956_ ), .C2(_12957_ ), .ZN(_00344_ ) );
OR2_X1 _19930_ ( .A1(_00313_ ), .A2(fanout_net_24 ), .ZN(_00345_ ) );
INV_X1 _19931_ ( .A(\wbu.io_in_bits_rd_wdata [31] ), .ZN(_12958_ ) );
NOR2_X1 _19932_ ( .A1(\wbu.io_in_bits_rd [0] ), .A2(\wbu.io_in_bits_rd [1] ), .ZN(_12959_ ) );
CLKBUF_X2 _19933_ ( .A(_12959_ ), .Z(_12960_ ) );
AND2_X1 _19934_ ( .A1(_08572_ ), .A2(_12960_ ), .ZN(_12961_ ) );
NAND2_X1 _19935_ ( .A1(_12961_ ), .A2(fanout_net_37 ), .ZN(_12962_ ) );
AND2_X1 _19936_ ( .A1(\ifu.io_valid ), .A2(\wbu.io_in_bits_wen_rd ), .ZN(_12963_ ) );
AND2_X2 _19937_ ( .A1(_12962_ ), .A2(_12963_ ), .ZN(_12964_ ) );
BUF_X4 _19938_ ( .A(_12964_ ), .Z(_12965_ ) );
AND2_X2 _19939_ ( .A1(\wbu.io_in_bits_rd [0] ), .A2(\wbu.io_in_bits_rd [1] ), .ZN(_12966_ ) );
AND2_X1 _19940_ ( .A1(\wbu.io_in_bits_rd [3] ), .A2(\wbu.io_in_bits_rd [2] ), .ZN(_12967_ ) );
AND2_X1 _19941_ ( .A1(_12966_ ), .A2(_12967_ ), .ZN(_12968_ ) );
AND2_X2 _19942_ ( .A1(_12968_ ), .A2(fanout_net_29 ), .ZN(_12969_ ) );
INV_X1 _19943_ ( .A(_12969_ ), .ZN(_12970_ ) );
BUF_X2 _19944_ ( .A(_12970_ ), .Z(_12971_ ) );
INV_X1 _19945_ ( .A(\wbu.io_in_bits_rd [0] ), .ZN(_12972_ ) );
AND3_X1 _19946_ ( .A1(_12967_ ), .A2(_12972_ ), .A3(\wbu.io_in_bits_rd [1] ), .ZN(_12973_ ) );
AND2_X1 _19947_ ( .A1(_12973_ ), .A2(fanout_net_29 ), .ZN(_12974_ ) );
BUF_X4 _19948_ ( .A(_12974_ ), .Z(_12975_ ) );
BUF_X2 _19949_ ( .A(_12975_ ), .Z(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ) );
NOR2_X1 _19950_ ( .A1(_08576_ ), .A2(\wbu.io_in_bits_rd [0] ), .ZN(_12976_ ) );
CLKBUF_X2 _19951_ ( .A(_12976_ ), .Z(_12977_ ) );
INV_X1 _19952_ ( .A(\wbu.io_in_bits_rd [3] ), .ZN(_12978_ ) );
NOR2_X1 _19953_ ( .A1(_12978_ ), .A2(\wbu.io_in_bits_rd [2] ), .ZN(_12979_ ) );
AND2_X1 _19954_ ( .A1(_12977_ ), .A2(_12979_ ), .ZN(_12980_ ) );
AND2_X1 _19955_ ( .A1(_12980_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _19956_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_12981_ ) );
BUF_X4 _19957_ ( .A(_12981_ ), .Z(_12982_ ) );
BUF_X4 _19958_ ( .A(_12982_ ), .Z(_12983_ ) );
BUF_X4 _19959_ ( .A(_12983_ ), .Z(_12984_ ) );
NOR2_X2 _19960_ ( .A1(_12972_ ), .A2(\wbu.io_in_bits_rd [1] ), .ZN(_12985_ ) );
BUF_X2 _19961_ ( .A(_12979_ ), .Z(_12986_ ) );
NAND4_X1 _19962_ ( .A1(_12985_ ), .A2(_12986_ ), .A3(fanout_net_37 ), .A4(\wbu.rf_9 [31] ), .ZN(_12987_ ) );
AND4_X1 _19963_ ( .A1(fanout_net_37 ), .A2(_12986_ ), .A3(\wbu.rf_8 [31] ), .A4(_12960_ ), .ZN(_12988_ ) );
AND3_X1 _19964_ ( .A1(_08572_ ), .A2(_12972_ ), .A3(\wbu.io_in_bits_rd [1] ), .ZN(_12989_ ) );
AND2_X2 _19965_ ( .A1(_12989_ ), .A2(fanout_net_37 ), .ZN(_12990_ ) );
BUF_X4 _19966_ ( .A(_12990_ ), .Z(_12991_ ) );
BUF_X4 _19967_ ( .A(_12991_ ), .Z(_12992_ ) );
BUF_X4 _19968_ ( .A(_12992_ ), .Z(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ) );
MUX2_X1 _19969_ ( .A(\wbu._GEN_71 [31] ), .B(\wbu.rf_2 [31] ), .S(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .Z(_12993_ ) );
AND2_X1 _19970_ ( .A1(_12966_ ), .A2(_08572_ ), .ZN(_12994_ ) );
AND2_X1 _19971_ ( .A1(_12994_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_Y ) );
INV_X1 _19972_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_Y ), .ZN(_12995_ ) );
BUF_X4 _19973_ ( .A(_12995_ ), .Z(_12996_ ) );
BUF_X4 _19974_ ( .A(_12996_ ), .Z(_12997_ ) );
BUF_X4 _19975_ ( .A(_12997_ ), .Z(_12998_ ) );
MUX2_X1 _19976_ ( .A(\wbu.rf_3 [31] ), .B(_12993_ ), .S(_12998_ ), .Z(_12999_ ) );
AND3_X1 _19977_ ( .A1(_12959_ ), .A2(_12978_ ), .A3(\wbu.io_in_bits_rd [2] ), .ZN(_13000_ ) );
AND2_X1 _19978_ ( .A1(_13000_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ) );
INV_X1 _19979_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ), .ZN(_13001_ ) );
BUF_X4 _19980_ ( .A(_13001_ ), .Z(_13002_ ) );
BUF_X4 _19981_ ( .A(_13002_ ), .Z(_13003_ ) );
BUF_X4 _19982_ ( .A(_13003_ ), .Z(_13004_ ) );
MUX2_X1 _19983_ ( .A(\wbu.rf_4 [31] ), .B(_12999_ ), .S(_13004_ ), .Z(_13005_ ) );
INV_X1 _19984_ ( .A(\wbu.io_in_bits_rd [2] ), .ZN(_13006_ ) );
NOR2_X2 _19985_ ( .A1(_13006_ ), .A2(\wbu.io_in_bits_rd [3] ), .ZN(_13007_ ) );
AND2_X2 _19986_ ( .A1(_12985_ ), .A2(_13007_ ), .ZN(_13008_ ) );
AND2_X1 _19987_ ( .A1(_13008_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _19988_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_13009_ ) );
BUF_X4 _19989_ ( .A(_13009_ ), .Z(_13010_ ) );
BUF_X4 _19990_ ( .A(_13010_ ), .Z(_13011_ ) );
BUF_X4 _19991_ ( .A(_13011_ ), .Z(_13012_ ) );
MUX2_X1 _19992_ ( .A(\wbu.rf_5 [31] ), .B(_13005_ ), .S(_13012_ ), .Z(_13013_ ) );
AND2_X1 _19993_ ( .A1(_12976_ ), .A2(_13007_ ), .ZN(_13014_ ) );
AND2_X1 _19994_ ( .A1(_13014_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_1_Y_$_ANDNOT__B_Y ) );
INV_X1 _19995_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .ZN(_13015_ ) );
BUF_X4 _19996_ ( .A(_13015_ ), .Z(_13016_ ) );
BUF_X4 _19997_ ( .A(_13016_ ), .Z(_13017_ ) );
BUF_X4 _19998_ ( .A(_13017_ ), .Z(_13018_ ) );
MUX2_X1 _19999_ ( .A(\wbu.rf_6 [31] ), .B(_13013_ ), .S(_13018_ ), .Z(_13019_ ) );
AND3_X1 _20000_ ( .A1(_12966_ ), .A2(_12978_ ), .A3(\wbu.io_in_bits_rd [2] ), .ZN(_13020_ ) );
AND2_X1 _20001_ ( .A1(_13020_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_Y ) );
INV_X1 _20002_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_Y ), .ZN(_13021_ ) );
BUF_X4 _20003_ ( .A(_13021_ ), .Z(_13022_ ) );
BUF_X4 _20004_ ( .A(_13022_ ), .Z(_13023_ ) );
BUF_X4 _20005_ ( .A(_13023_ ), .Z(_13024_ ) );
MUX2_X1 _20006_ ( .A(\wbu.rf_7 [31] ), .B(_13019_ ), .S(_13024_ ), .Z(_13025_ ) );
AND3_X1 _20007_ ( .A1(_12959_ ), .A2(\wbu.io_in_bits_rd [3] ), .A3(_13006_ ), .ZN(_13026_ ) );
AND2_X1 _20008_ ( .A1(_13026_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_Y ) );
INV_X1 _20009_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_Y ), .ZN(_13027_ ) );
BUF_X4 _20010_ ( .A(_13027_ ), .Z(_13028_ ) );
BUF_X4 _20011_ ( .A(_13028_ ), .Z(_13029_ ) );
BUF_X2 _20012_ ( .A(_13029_ ), .Z(_13030_ ) );
AOI21_X1 _20013_ ( .A(_12988_ ), .B1(_13025_ ), .B2(_13030_ ), .ZN(_13031_ ) );
AND2_X1 _20014_ ( .A1(_12985_ ), .A2(_12979_ ), .ZN(_13032_ ) );
AND2_X2 _20015_ ( .A1(_13032_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_Y ) );
OAI211_X1 _20016_ ( .A(_12984_ ), .B(_12987_ ), .C1(_13031_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_Y ), .ZN(_13033_ ) );
AND3_X1 _20017_ ( .A1(_12966_ ), .A2(\wbu.io_in_bits_rd [3] ), .A3(_13006_ ), .ZN(_13034_ ) );
AND2_X1 _20018_ ( .A1(_13034_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_1_Y_$_ANDNOT__B_Y ) );
INV_X1 _20019_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .ZN(_13035_ ) );
BUF_X4 _20020_ ( .A(_13035_ ), .Z(_13036_ ) );
BUF_X4 _20021_ ( .A(_13036_ ), .Z(_13037_ ) );
BUF_X4 _20022_ ( .A(_13037_ ), .Z(_13038_ ) );
BUF_X4 _20023_ ( .A(_12984_ ), .Z(_13039_ ) );
OAI211_X1 _20024_ ( .A(_13033_ ), .B(_13038_ ), .C1(\wbu.rf_10 [31] ), .C2(_13039_ ), .ZN(_13040_ ) );
AND2_X1 _20025_ ( .A1(_12967_ ), .A2(_12960_ ), .ZN(_13041_ ) );
AND2_X1 _20026_ ( .A1(_13041_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _20027_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_13042_ ) );
BUF_X4 _20028_ ( .A(_13042_ ), .Z(_13043_ ) );
BUF_X4 _20029_ ( .A(_13043_ ), .Z(_13044_ ) );
BUF_X4 _20030_ ( .A(_13044_ ), .Z(_13045_ ) );
BUF_X4 _20031_ ( .A(_12986_ ), .Z(_13046_ ) );
BUF_X4 _20032_ ( .A(_12966_ ), .Z(_13047_ ) );
NAND4_X1 _20033_ ( .A1(_13046_ ), .A2(fanout_net_37 ), .A3(_13047_ ), .A4(\wbu.rf_11 [31] ), .ZN(_13048_ ) );
NAND3_X1 _20034_ ( .A1(_13040_ ), .A2(_13045_ ), .A3(_13048_ ), .ZN(_13049_ ) );
AND3_X1 _20035_ ( .A1(_12967_ ), .A2(\wbu.io_in_bits_rd [0] ), .A3(_08576_ ), .ZN(_13050_ ) );
AND2_X1 _20036_ ( .A1(_13050_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _20037_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_13051_ ) );
BUF_X4 _20038_ ( .A(_13051_ ), .Z(_13052_ ) );
BUF_X4 _20039_ ( .A(_13052_ ), .Z(_13053_ ) );
BUF_X2 _20040_ ( .A(_13053_ ), .Z(_13054_ ) );
BUF_X4 _20041_ ( .A(_13045_ ), .Z(_13055_ ) );
OAI211_X1 _20042_ ( .A(_13049_ ), .B(_13054_ ), .C1(\wbu.rf_12 [31] ), .C2(_13055_ ), .ZN(_13056_ ) );
AND2_X1 _20043_ ( .A1(_12973_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _20044_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_13057_ ) );
BUF_X4 _20045_ ( .A(_13057_ ), .Z(_13058_ ) );
BUF_X4 _20046_ ( .A(_13058_ ), .Z(_13059_ ) );
BUF_X4 _20047_ ( .A(_13059_ ), .Z(_13060_ ) );
BUF_X4 _20048_ ( .A(_12985_ ), .Z(_13061_ ) );
BUF_X4 _20049_ ( .A(_13061_ ), .Z(_13062_ ) );
BUF_X2 _20050_ ( .A(_12967_ ), .Z(_13063_ ) );
BUF_X2 _20051_ ( .A(_13063_ ), .Z(_13064_ ) );
NAND4_X1 _20052_ ( .A1(_13062_ ), .A2(fanout_net_37 ), .A3(_13064_ ), .A4(\wbu.rf_13 [31] ), .ZN(_13065_ ) );
NAND3_X1 _20053_ ( .A1(_13056_ ), .A2(_13060_ ), .A3(_13065_ ), .ZN(_13066_ ) );
AND2_X2 _20054_ ( .A1(_12968_ ), .A2(fanout_net_37 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ) );
INV_X1 _20055_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .ZN(_13067_ ) );
BUF_X4 _20056_ ( .A(_13067_ ), .Z(_13068_ ) );
BUF_X4 _20057_ ( .A(_13068_ ), .Z(_13069_ ) );
BUF_X4 _20058_ ( .A(_13069_ ), .Z(_13070_ ) );
BUF_X4 _20059_ ( .A(_13059_ ), .Z(_13071_ ) );
OAI211_X1 _20060_ ( .A(_13066_ ), .B(_13070_ ), .C1(\wbu.rf_14 [31] ), .C2(_13071_ ), .ZN(_13072_ ) );
AND2_X1 _20061_ ( .A1(_12961_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__B_Y ) );
INV_X1 _20062_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__B_Y ), .ZN(_13073_ ) );
BUF_X4 _20063_ ( .A(_13073_ ), .Z(_13074_ ) );
BUF_X4 _20064_ ( .A(_13074_ ), .Z(_13075_ ) );
BUF_X4 _20065_ ( .A(_13075_ ), .Z(_13076_ ) );
BUF_X4 _20066_ ( .A(_13047_ ), .Z(_13077_ ) );
BUF_X4 _20067_ ( .A(_13063_ ), .Z(_13078_ ) );
BUF_X4 _20068_ ( .A(_13078_ ), .Z(_13079_ ) );
NAND4_X1 _20069_ ( .A1(_13077_ ), .A2(_13079_ ), .A3(fanout_net_37 ), .A4(\wbu.rf_15 [31] ), .ZN(_13080_ ) );
NAND3_X1 _20070_ ( .A1(_13072_ ), .A2(_13076_ ), .A3(_13080_ ), .ZN(_13081_ ) );
AND3_X1 _20071_ ( .A1(_08572_ ), .A2(\wbu.io_in_bits_rd [0] ), .A3(_08576_ ), .ZN(_13082_ ) );
AND2_X1 _20072_ ( .A1(_13082_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _20073_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_13083_ ) );
BUF_X4 _20074_ ( .A(_13083_ ), .Z(_13084_ ) );
BUF_X4 _20075_ ( .A(_13084_ ), .Z(_13085_ ) );
BUF_X4 _20076_ ( .A(_13085_ ), .Z(_13086_ ) );
BUF_X4 _20077_ ( .A(_13075_ ), .Z(_13087_ ) );
OAI211_X1 _20078_ ( .A(_13081_ ), .B(_13086_ ), .C1(\wbu.rf_16 [31] ), .C2(_13087_ ), .ZN(_13088_ ) );
AND2_X1 _20079_ ( .A1(_12989_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ) );
INV_X1 _20080_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .ZN(_13089_ ) );
BUF_X4 _20081_ ( .A(_13089_ ), .Z(_13090_ ) );
BUF_X4 _20082_ ( .A(_13090_ ), .Z(_13091_ ) );
BUF_X4 _20083_ ( .A(_13062_ ), .Z(_13092_ ) );
NAND4_X1 _20084_ ( .A1(_13092_ ), .A2(fanout_net_29 ), .A3(\wbu.rf_17 [31] ), .A4(_08574_ ), .ZN(_13093_ ) );
NAND3_X1 _20085_ ( .A1(_13088_ ), .A2(_13091_ ), .A3(_13093_ ), .ZN(_13094_ ) );
AND2_X1 _20086_ ( .A1(_12994_ ), .A2(fanout_net_29 ), .ZN(_13095_ ) );
INV_X2 _20087_ ( .A(_13095_ ), .ZN(_13096_ ) );
BUF_X4 _20088_ ( .A(_13096_ ), .Z(_13097_ ) );
BUF_X2 _20089_ ( .A(_13097_ ), .Z(_13098_ ) );
BUF_X4 _20090_ ( .A(_13091_ ), .Z(_13099_ ) );
OAI211_X1 _20091_ ( .A(_13094_ ), .B(_13098_ ), .C1(\wbu.rf_18 [31] ), .C2(_13099_ ), .ZN(_13100_ ) );
AND2_X1 _20092_ ( .A1(_13000_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_1_Y ) );
INV_X1 _20093_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .ZN(_13101_ ) );
BUF_X4 _20094_ ( .A(_13101_ ), .Z(_13102_ ) );
BUF_X4 _20095_ ( .A(_13102_ ), .Z(_13103_ ) );
BUF_X4 _20096_ ( .A(_13103_ ), .Z(_13104_ ) );
BUF_X4 _20097_ ( .A(_13077_ ), .Z(_13105_ ) );
BUF_X4 _20098_ ( .A(_13105_ ), .Z(_13106_ ) );
NAND4_X1 _20099_ ( .A1(_13106_ ), .A2(_08575_ ), .A3(fanout_net_29 ), .A4(\wbu.rf_19 [31] ), .ZN(_13107_ ) );
NAND3_X1 _20100_ ( .A1(_13100_ ), .A2(_13104_ ), .A3(_13107_ ), .ZN(_13108_ ) );
AND2_X1 _20101_ ( .A1(_13008_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_1_Y ) );
INV_X1 _20102_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_13109_ ) );
BUF_X4 _20103_ ( .A(_13109_ ), .Z(_13110_ ) );
BUF_X4 _20104_ ( .A(_13110_ ), .Z(_13111_ ) );
BUF_X4 _20105_ ( .A(_13111_ ), .Z(_13112_ ) );
BUF_X4 _20106_ ( .A(_13103_ ), .Z(_13113_ ) );
OAI211_X1 _20107_ ( .A(_13108_ ), .B(_13112_ ), .C1(\wbu.rf_20 [31] ), .C2(_13113_ ), .ZN(_13114_ ) );
AND2_X1 _20108_ ( .A1(_13014_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ) );
INV_X1 _20109_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .ZN(_13115_ ) );
BUF_X4 _20110_ ( .A(_13115_ ), .Z(_13116_ ) );
BUF_X4 _20111_ ( .A(_13116_ ), .Z(_13117_ ) );
BUF_X4 _20112_ ( .A(_13117_ ), .Z(_13118_ ) );
BUF_X4 _20113_ ( .A(_13062_ ), .Z(_13119_ ) );
BUF_X4 _20114_ ( .A(_13119_ ), .Z(_13120_ ) );
BUF_X4 _20115_ ( .A(_13007_ ), .Z(_13121_ ) );
BUF_X4 _20116_ ( .A(_13121_ ), .Z(_13122_ ) );
NAND4_X1 _20117_ ( .A1(_13120_ ), .A2(_13122_ ), .A3(fanout_net_29 ), .A4(\wbu.rf_21 [31] ), .ZN(_13123_ ) );
NAND3_X1 _20118_ ( .A1(_13114_ ), .A2(_13118_ ), .A3(_13123_ ), .ZN(_13124_ ) );
AND2_X1 _20119_ ( .A1(_13020_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ) );
INV_X1 _20120_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .ZN(_13125_ ) );
BUF_X4 _20121_ ( .A(_13125_ ), .Z(_13126_ ) );
BUF_X4 _20122_ ( .A(_13126_ ), .Z(_13127_ ) );
BUF_X4 _20123_ ( .A(_13117_ ), .Z(_13128_ ) );
OAI211_X1 _20124_ ( .A(_13124_ ), .B(_13127_ ), .C1(\wbu.rf_22 [31] ), .C2(_13128_ ), .ZN(_13129_ ) );
AND2_X2 _20125_ ( .A1(_13026_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_1_Y ) );
INV_X2 _20126_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_1_Y ), .ZN(_13130_ ) );
BUF_X4 _20127_ ( .A(_13130_ ), .Z(_13131_ ) );
BUF_X4 _20128_ ( .A(_13131_ ), .Z(_13132_ ) );
BUF_X4 _20129_ ( .A(_13122_ ), .Z(_13133_ ) );
BUF_X4 _20130_ ( .A(_13105_ ), .Z(_13134_ ) );
BUF_X4 _20131_ ( .A(_13134_ ), .Z(_13135_ ) );
NAND4_X1 _20132_ ( .A1(_13133_ ), .A2(fanout_net_29 ), .A3(_13135_ ), .A4(\wbu.rf_23 [31] ), .ZN(_13136_ ) );
NAND3_X1 _20133_ ( .A1(_13129_ ), .A2(_13132_ ), .A3(_13136_ ), .ZN(_13137_ ) );
AND2_X2 _20134_ ( .A1(_13032_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ) );
INV_X1 _20135_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .ZN(_13138_ ) );
BUF_X4 _20136_ ( .A(_13138_ ), .Z(_13139_ ) );
BUF_X4 _20137_ ( .A(_13139_ ), .Z(_13140_ ) );
BUF_X4 _20138_ ( .A(_13131_ ), .Z(_13141_ ) );
OAI211_X1 _20139_ ( .A(_13137_ ), .B(_13140_ ), .C1(\wbu.rf_24 [31] ), .C2(_13141_ ), .ZN(_13142_ ) );
AND2_X1 _20140_ ( .A1(_12980_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_Y_$_ANDNOT__B_1_Y ) );
INV_X2 _20141_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_13143_ ) );
BUF_X4 _20142_ ( .A(_13143_ ), .Z(_13144_ ) );
BUF_X4 _20143_ ( .A(_13144_ ), .Z(_13145_ ) );
BUF_X2 _20144_ ( .A(_13119_ ), .Z(_13146_ ) );
BUF_X2 _20145_ ( .A(_13146_ ), .Z(_13147_ ) );
BUF_X4 _20146_ ( .A(_13046_ ), .Z(_13148_ ) );
BUF_X4 _20147_ ( .A(_13148_ ), .Z(_13149_ ) );
NAND4_X1 _20148_ ( .A1(_13147_ ), .A2(_13149_ ), .A3(fanout_net_29 ), .A4(\wbu.rf_25 [31] ), .ZN(_13150_ ) );
NAND3_X1 _20149_ ( .A1(_13142_ ), .A2(_13145_ ), .A3(_13150_ ), .ZN(_13151_ ) );
AND2_X1 _20150_ ( .A1(_13034_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ) );
INV_X2 _20151_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .ZN(_13152_ ) );
BUF_X2 _20152_ ( .A(_13152_ ), .Z(_13153_ ) );
BUF_X4 _20153_ ( .A(_13144_ ), .Z(_13154_ ) );
OAI211_X1 _20154_ ( .A(_13151_ ), .B(_13153_ ), .C1(\wbu.rf_26 [31] ), .C2(_13154_ ), .ZN(_13155_ ) );
AND2_X2 _20155_ ( .A1(_13041_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_1_Y ) );
INV_X2 _20156_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_13156_ ) );
BUF_X4 _20157_ ( .A(_13156_ ), .Z(_13157_ ) );
BUF_X4 _20158_ ( .A(_13148_ ), .Z(_13158_ ) );
BUF_X4 _20159_ ( .A(_13158_ ), .Z(_13159_ ) );
BUF_X4 _20160_ ( .A(_13135_ ), .Z(_13160_ ) );
BUF_X4 _20161_ ( .A(_13160_ ), .Z(_13161_ ) );
NAND4_X1 _20162_ ( .A1(_13159_ ), .A2(fanout_net_29 ), .A3(_13161_ ), .A4(\wbu.rf_27 [31] ), .ZN(_13162_ ) );
NAND3_X1 _20163_ ( .A1(_13155_ ), .A2(_13157_ ), .A3(_13162_ ), .ZN(_13163_ ) );
AND2_X1 _20164_ ( .A1(_13050_ ), .A2(fanout_net_29 ), .ZN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ) );
INV_X2 _20165_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_13164_ ) );
BUF_X4 _20166_ ( .A(_13164_ ), .Z(_13165_ ) );
BUF_X4 _20167_ ( .A(_13156_ ), .Z(_13166_ ) );
BUF_X4 _20168_ ( .A(_13166_ ), .Z(_13167_ ) );
OAI211_X1 _20169_ ( .A(_13163_ ), .B(_13165_ ), .C1(\wbu.rf_28 [31] ), .C2(_13167_ ), .ZN(_13168_ ) );
BUF_X4 _20170_ ( .A(_13147_ ), .Z(_13169_ ) );
BUF_X4 _20171_ ( .A(_13079_ ), .Z(_13170_ ) );
NAND4_X1 _20172_ ( .A1(_13169_ ), .A2(fanout_net_29 ), .A3(_13170_ ), .A4(\wbu.rf_29 [31] ), .ZN(_13171_ ) );
AOI21_X1 _20173_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .B1(_13168_ ), .B2(_13171_ ), .ZN(_13172_ ) );
BUF_X2 _20174_ ( .A(_12977_ ), .Z(_13173_ ) );
BUF_X2 _20175_ ( .A(_13173_ ), .Z(_13174_ ) );
CLKBUF_X2 _20176_ ( .A(_13174_ ), .Z(_13175_ ) );
BUF_X2 _20177_ ( .A(_13079_ ), .Z(_13176_ ) );
AND4_X1 _20178_ ( .A1(fanout_net_29 ), .A2(_13175_ ), .A3(\wbu.rf_30 [31] ), .A4(_13176_ ), .ZN(_13177_ ) );
OAI21_X1 _20179_ ( .A(_12971_ ), .B1(_13172_ ), .B2(_13177_ ), .ZN(_13178_ ) );
BUF_X4 _20180_ ( .A(_12969_ ), .Z(_13179_ ) );
BUF_X2 _20181_ ( .A(_12962_ ), .Z(_13180_ ) );
BUF_X2 _20182_ ( .A(_13180_ ), .Z(_13181_ ) );
BUF_X2 _20183_ ( .A(_12963_ ), .Z(_13182_ ) );
BUF_X2 _20184_ ( .A(_13182_ ), .Z(_13183_ ) );
AOI22_X1 _20185_ ( .A1(_13179_ ), .A2(\wbu.rf_31 [31] ), .B1(_13181_ ), .B2(_13183_ ), .ZN(_13184_ ) );
AOI221_X4 _20186_ ( .A(fanout_net_24 ), .B1(_12958_ ), .B2(_12965_ ), .C1(_13178_ ), .C2(_13184_ ), .ZN(_00346_ ) );
INV_X1 _20187_ ( .A(\wbu.io_in_bits_rd_wdata [30] ), .ZN(_13185_ ) );
BUF_X4 _20188_ ( .A(_13122_ ), .Z(_13186_ ) );
NAND4_X1 _20189_ ( .A1(_13186_ ), .A2(fanout_net_29 ), .A3(_13134_ ), .A4(\wbu.rf_23 [30] ), .ZN(_13187_ ) );
BUF_X2 _20190_ ( .A(_13121_ ), .Z(_13188_ ) );
AND4_X1 _20191_ ( .A1(fanout_net_29 ), .A2(_13174_ ), .A3(_13188_ ), .A4(\wbu.rf_22 [30] ), .ZN(_13189_ ) );
MUX2_X1 _20192_ ( .A(\wbu._GEN_71 [30] ), .B(\wbu.rf_2 [30] ), .S(_12991_ ), .Z(_13190_ ) );
MUX2_X1 _20193_ ( .A(\wbu.rf_3 [30] ), .B(_13190_ ), .S(_12996_ ), .Z(_13191_ ) );
MUX2_X1 _20194_ ( .A(\wbu.rf_4 [30] ), .B(_13191_ ), .S(_13002_ ), .Z(_13192_ ) );
MUX2_X1 _20195_ ( .A(\wbu.rf_5 [30] ), .B(_13192_ ), .S(_13010_ ), .Z(_13193_ ) );
MUX2_X1 _20196_ ( .A(\wbu.rf_6 [30] ), .B(_13193_ ), .S(_13016_ ), .Z(_13194_ ) );
MUX2_X1 _20197_ ( .A(\wbu.rf_7 [30] ), .B(_13194_ ), .S(_13022_ ), .Z(_13195_ ) );
MUX2_X1 _20198_ ( .A(\wbu.rf_8 [30] ), .B(_13195_ ), .S(_13028_ ), .Z(_13196_ ) );
INV_X2 _20199_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_Y ), .ZN(_13197_ ) );
BUF_X4 _20200_ ( .A(_13197_ ), .Z(_13198_ ) );
MUX2_X1 _20201_ ( .A(\wbu.rf_9 [30] ), .B(_13196_ ), .S(_13198_ ), .Z(_13199_ ) );
MUX2_X1 _20202_ ( .A(\wbu.rf_10 [30] ), .B(_13199_ ), .S(_12983_ ), .Z(_13200_ ) );
MUX2_X1 _20203_ ( .A(\wbu.rf_11 [30] ), .B(_13200_ ), .S(_13036_ ), .Z(_13201_ ) );
MUX2_X1 _20204_ ( .A(\wbu.rf_12 [30] ), .B(_13201_ ), .S(_13043_ ), .Z(_13202_ ) );
MUX2_X1 _20205_ ( .A(\wbu.rf_13 [30] ), .B(_13202_ ), .S(_13052_ ), .Z(_13203_ ) );
MUX2_X1 _20206_ ( .A(\wbu.rf_14 [30] ), .B(_13203_ ), .S(_13058_ ), .Z(_13204_ ) );
MUX2_X1 _20207_ ( .A(\wbu.rf_15 [30] ), .B(_13204_ ), .S(_13068_ ), .Z(_13205_ ) );
MUX2_X1 _20208_ ( .A(\wbu.rf_16 [30] ), .B(_13205_ ), .S(_13074_ ), .Z(_13206_ ) );
MUX2_X1 _20209_ ( .A(\wbu.rf_17 [30] ), .B(_13206_ ), .S(_13084_ ), .Z(_13207_ ) );
MUX2_X1 _20210_ ( .A(\wbu.rf_18 [30] ), .B(_13207_ ), .S(_13090_ ), .Z(_13208_ ) );
MUX2_X1 _20211_ ( .A(\wbu.rf_19 [30] ), .B(_13208_ ), .S(_13097_ ), .Z(_13209_ ) );
MUX2_X1 _20212_ ( .A(\wbu.rf_20 [30] ), .B(_13209_ ), .S(_13103_ ), .Z(_13210_ ) );
MUX2_X1 _20213_ ( .A(\wbu.rf_21 [30] ), .B(_13210_ ), .S(_13111_ ), .Z(_13211_ ) );
BUF_X4 _20214_ ( .A(_13117_ ), .Z(_13212_ ) );
AOI21_X1 _20215_ ( .A(_13189_ ), .B1(_13211_ ), .B2(_13212_ ), .ZN(_13213_ ) );
OAI211_X1 _20216_ ( .A(_13132_ ), .B(_13187_ ), .C1(_13213_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .ZN(_13214_ ) );
OAI211_X1 _20217_ ( .A(_13214_ ), .B(_13140_ ), .C1(\wbu.rf_24 [30] ), .C2(_13141_ ), .ZN(_13215_ ) );
NAND4_X1 _20218_ ( .A1(_13147_ ), .A2(_13149_ ), .A3(fanout_net_29 ), .A4(\wbu.rf_25 [30] ), .ZN(_13216_ ) );
NAND3_X1 _20219_ ( .A1(_13215_ ), .A2(_13145_ ), .A3(_13216_ ), .ZN(_13217_ ) );
BUF_X4 _20220_ ( .A(_13152_ ), .Z(_13218_ ) );
OAI211_X1 _20221_ ( .A(_13217_ ), .B(_13218_ ), .C1(\wbu.rf_26 [30] ), .C2(_13154_ ), .ZN(_13219_ ) );
NAND4_X1 _20222_ ( .A1(_13159_ ), .A2(fanout_net_29 ), .A3(_13161_ ), .A4(\wbu.rf_27 [30] ), .ZN(_13220_ ) );
NAND3_X1 _20223_ ( .A1(_13219_ ), .A2(_13157_ ), .A3(_13220_ ), .ZN(_13221_ ) );
OAI211_X1 _20224_ ( .A(_13221_ ), .B(_13165_ ), .C1(\wbu.rf_28 [30] ), .C2(_13167_ ), .ZN(_13222_ ) );
NAND4_X1 _20225_ ( .A1(_13169_ ), .A2(fanout_net_29 ), .A3(_13170_ ), .A4(\wbu.rf_29 [30] ), .ZN(_13223_ ) );
AOI21_X1 _20226_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .B1(_13222_ ), .B2(_13223_ ), .ZN(_13224_ ) );
AND4_X1 _20227_ ( .A1(fanout_net_30 ), .A2(_13175_ ), .A3(\wbu.rf_30 [30] ), .A4(_13176_ ), .ZN(_13225_ ) );
OAI21_X1 _20228_ ( .A(_12971_ ), .B1(_13224_ ), .B2(_13225_ ), .ZN(_13226_ ) );
AOI22_X1 _20229_ ( .A1(_13179_ ), .A2(\wbu.rf_31 [30] ), .B1(_13181_ ), .B2(_13183_ ), .ZN(_13227_ ) );
AOI221_X4 _20230_ ( .A(fanout_net_24 ), .B1(_13185_ ), .B2(_12965_ ), .C1(_13226_ ), .C2(_13227_ ), .ZN(_00347_ ) );
BUF_X2 _20231_ ( .A(_12960_ ), .Z(_13228_ ) );
BUF_X2 _20232_ ( .A(_13228_ ), .Z(_13229_ ) );
NAND4_X1 _20233_ ( .A1(_13170_ ), .A2(_13229_ ), .A3(fanout_net_30 ), .A4(\wbu.rf_28 [21] ), .ZN(_13230_ ) );
BUF_X4 _20234_ ( .A(_13126_ ), .Z(_13231_ ) );
NOR2_X1 _20235_ ( .A1(_13231_ ), .A2(\wbu.rf_23 [21] ), .ZN(_13232_ ) );
OR2_X1 _20236_ ( .A1(_13098_ ), .A2(\wbu.rf_19 [21] ), .ZN(_13233_ ) );
MUX2_X1 _20237_ ( .A(\wbu._GEN_71 [21] ), .B(\wbu.rf_2 [21] ), .S(_12991_ ), .Z(_13234_ ) );
MUX2_X1 _20238_ ( .A(\wbu.rf_3 [21] ), .B(_13234_ ), .S(_12997_ ), .Z(_13235_ ) );
MUX2_X1 _20239_ ( .A(\wbu.rf_4 [21] ), .B(_13235_ ), .S(_13003_ ), .Z(_13236_ ) );
MUX2_X1 _20240_ ( .A(\wbu.rf_5 [21] ), .B(_13236_ ), .S(_13011_ ), .Z(_13237_ ) );
MUX2_X1 _20241_ ( .A(\wbu.rf_6 [21] ), .B(_13237_ ), .S(_13016_ ), .Z(_13238_ ) );
MUX2_X1 _20242_ ( .A(\wbu.rf_7 [21] ), .B(_13238_ ), .S(_13023_ ), .Z(_13239_ ) );
MUX2_X1 _20243_ ( .A(\wbu.rf_8 [21] ), .B(_13239_ ), .S(_13029_ ), .Z(_13240_ ) );
MUX2_X1 _20244_ ( .A(\wbu.rf_9 [21] ), .B(_13240_ ), .S(_13198_ ), .Z(_13241_ ) );
MUX2_X1 _20245_ ( .A(\wbu.rf_10 [21] ), .B(_13241_ ), .S(_12983_ ), .Z(_13242_ ) );
MUX2_X1 _20246_ ( .A(\wbu.rf_11 [21] ), .B(_13242_ ), .S(_13037_ ), .Z(_13243_ ) );
MUX2_X1 _20247_ ( .A(\wbu.rf_12 [21] ), .B(_13243_ ), .S(_13044_ ), .Z(_13244_ ) );
MUX2_X1 _20248_ ( .A(\wbu.rf_13 [21] ), .B(_13244_ ), .S(_13053_ ), .Z(_13245_ ) );
MUX2_X1 _20249_ ( .A(\wbu.rf_14 [21] ), .B(_13245_ ), .S(_13059_ ), .Z(_13246_ ) );
MUX2_X1 _20250_ ( .A(\wbu.rf_15 [21] ), .B(_13246_ ), .S(_13069_ ), .Z(_13247_ ) );
MUX2_X1 _20251_ ( .A(\wbu.rf_16 [21] ), .B(_13247_ ), .S(_13075_ ), .Z(_13248_ ) );
MUX2_X1 _20252_ ( .A(\wbu.rf_17 [21] ), .B(_13248_ ), .S(_13085_ ), .Z(_13249_ ) );
MUX2_X1 _20253_ ( .A(\wbu.rf_18 [21] ), .B(_13249_ ), .S(_13099_ ), .Z(_13250_ ) );
BUF_X2 _20254_ ( .A(_13095_ ), .Z(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ) );
OAI211_X1 _20255_ ( .A(_13113_ ), .B(_13233_ ), .C1(_13250_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .ZN(_13251_ ) );
NAND4_X1 _20256_ ( .A1(_13122_ ), .A2(fanout_net_30 ), .A3(\wbu.rf_20 [21] ), .A4(_13228_ ), .ZN(_13252_ ) );
AOI21_X1 _20257_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_1_Y ), .B1(_13251_ ), .B2(_13252_ ), .ZN(_13253_ ) );
AND3_X1 _20258_ ( .A1(_13008_ ), .A2(fanout_net_30 ), .A3(\wbu.rf_21 [21] ), .ZN(_13254_ ) );
OAI21_X1 _20259_ ( .A(_13128_ ), .B1(_13253_ ), .B2(_13254_ ), .ZN(_13255_ ) );
AOI21_X1 _20260_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .B1(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .B2(\wbu.rf_22 [21] ), .ZN(_13256_ ) );
AOI211_X1 _20261_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_1_Y ), .B(_13232_ ), .C1(_13255_ ), .C2(_13256_ ), .ZN(_13257_ ) );
AND4_X1 _20262_ ( .A1(fanout_net_30 ), .A2(_13148_ ), .A3(\wbu.rf_24 [21] ), .A4(_13229_ ), .ZN(_13258_ ) );
OAI21_X1 _20263_ ( .A(_13140_ ), .B1(_13257_ ), .B2(_13258_ ), .ZN(_13259_ ) );
BUF_X2 _20264_ ( .A(_13144_ ), .Z(_13260_ ) );
NAND3_X1 _20265_ ( .A1(_13032_ ), .A2(fanout_net_30 ), .A3(\wbu.rf_25 [21] ), .ZN(_13261_ ) );
AND3_X1 _20266_ ( .A1(_13259_ ), .A2(_13260_ ), .A3(_13261_ ), .ZN(_13262_ ) );
NOR2_X1 _20267_ ( .A1(_13154_ ), .A2(\wbu.rf_26 [21] ), .ZN(_13263_ ) );
OAI21_X1 _20268_ ( .A(_13153_ ), .B1(_13262_ ), .B2(_13263_ ), .ZN(_13264_ ) );
OAI21_X1 _20269_ ( .A(_13264_ ), .B1(\wbu.rf_27 [21] ), .B2(_13153_ ), .ZN(_13265_ ) );
OAI211_X1 _20270_ ( .A(_13165_ ), .B(_13230_ ), .C1(_13265_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_13266_ ) );
INV_X1 _20271_ ( .A(_12975_ ), .ZN(_13267_ ) );
BUF_X4 _20272_ ( .A(_13267_ ), .Z(_13268_ ) );
BUF_X4 _20273_ ( .A(_13165_ ), .Z(_13269_ ) );
OAI211_X1 _20274_ ( .A(_13266_ ), .B(_13268_ ), .C1(\wbu.rf_29 [21] ), .C2(_13269_ ), .ZN(_13270_ ) );
BUF_X4 _20275_ ( .A(_12970_ ), .Z(_13271_ ) );
BUF_X4 _20276_ ( .A(_13175_ ), .Z(_13272_ ) );
BUF_X4 _20277_ ( .A(_13170_ ), .Z(_13273_ ) );
NAND4_X1 _20278_ ( .A1(_13272_ ), .A2(fanout_net_30 ), .A3(_13273_ ), .A4(\wbu.rf_30 [21] ), .ZN(_13274_ ) );
NAND3_X1 _20279_ ( .A1(_13270_ ), .A2(_13271_ ), .A3(_13274_ ), .ZN(_13275_ ) );
INV_X2 _20280_ ( .A(_12964_ ), .ZN(_13276_ ) );
OAI211_X1 _20281_ ( .A(_13275_ ), .B(_13276_ ), .C1(\wbu.rf_31 [21] ), .C2(_13271_ ), .ZN(_13277_ ) );
NAND3_X1 _20282_ ( .A1(_13181_ ), .A2(\wbu.io_in_bits_rd_wdata [21] ), .A3(_13183_ ), .ZN(_13278_ ) );
AOI21_X1 _20283_ ( .A(fanout_net_24 ), .B1(_13277_ ), .B2(_13278_ ), .ZN(_00348_ ) );
INV_X1 _20284_ ( .A(\wbu.io_in_bits_rd_wdata [20] ), .ZN(_13279_ ) );
NAND4_X1 _20285_ ( .A1(_12985_ ), .A2(_12986_ ), .A3(fanout_net_37 ), .A4(\wbu.rf_9 [20] ), .ZN(_13280_ ) );
AND4_X1 _20286_ ( .A1(fanout_net_37 ), .A2(_12986_ ), .A3(\wbu.rf_8 [20] ), .A4(_12960_ ), .ZN(_13281_ ) );
MUX2_X1 _20287_ ( .A(\wbu._GEN_71 [20] ), .B(\wbu.rf_2 [20] ), .S(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .Z(_13282_ ) );
MUX2_X1 _20288_ ( .A(\wbu.rf_3 [20] ), .B(_13282_ ), .S(_12998_ ), .Z(_13283_ ) );
MUX2_X1 _20289_ ( .A(\wbu.rf_4 [20] ), .B(_13283_ ), .S(_13004_ ), .Z(_13284_ ) );
MUX2_X1 _20290_ ( .A(\wbu.rf_5 [20] ), .B(_13284_ ), .S(_13012_ ), .Z(_13285_ ) );
MUX2_X1 _20291_ ( .A(\wbu.rf_6 [20] ), .B(_13285_ ), .S(_13018_ ), .Z(_13286_ ) );
MUX2_X1 _20292_ ( .A(\wbu.rf_7 [20] ), .B(_13286_ ), .S(_13024_ ), .Z(_13287_ ) );
AOI21_X1 _20293_ ( .A(_13281_ ), .B1(_13287_ ), .B2(_13030_ ), .ZN(_13288_ ) );
OAI211_X1 _20294_ ( .A(_12984_ ), .B(_13280_ ), .C1(_13288_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_Y ), .ZN(_13289_ ) );
OAI211_X1 _20295_ ( .A(_13289_ ), .B(_13038_ ), .C1(\wbu.rf_10 [20] ), .C2(_13039_ ), .ZN(_13290_ ) );
NAND4_X1 _20296_ ( .A1(_13046_ ), .A2(fanout_net_37 ), .A3(_13047_ ), .A4(\wbu.rf_11 [20] ), .ZN(_13291_ ) );
NAND3_X1 _20297_ ( .A1(_13290_ ), .A2(_13045_ ), .A3(_13291_ ), .ZN(_13292_ ) );
OAI211_X1 _20298_ ( .A(_13292_ ), .B(_13054_ ), .C1(\wbu.rf_12 [20] ), .C2(_13055_ ), .ZN(_13293_ ) );
NAND4_X1 _20299_ ( .A1(_13062_ ), .A2(fanout_net_37 ), .A3(_13064_ ), .A4(\wbu.rf_13 [20] ), .ZN(_13294_ ) );
NAND3_X1 _20300_ ( .A1(_13293_ ), .A2(_13060_ ), .A3(_13294_ ), .ZN(_13295_ ) );
OAI211_X1 _20301_ ( .A(_13295_ ), .B(_13070_ ), .C1(\wbu.rf_14 [20] ), .C2(_13071_ ), .ZN(_13296_ ) );
NAND4_X1 _20302_ ( .A1(_13077_ ), .A2(_13079_ ), .A3(fanout_net_37 ), .A4(\wbu.rf_15 [20] ), .ZN(_13297_ ) );
NAND3_X1 _20303_ ( .A1(_13296_ ), .A2(_13076_ ), .A3(_13297_ ), .ZN(_13298_ ) );
OAI211_X1 _20304_ ( .A(_13298_ ), .B(_13086_ ), .C1(\wbu.rf_16 [20] ), .C2(_13087_ ), .ZN(_13299_ ) );
NAND4_X1 _20305_ ( .A1(_13092_ ), .A2(fanout_net_30 ), .A3(\wbu.rf_17 [20] ), .A4(_08574_ ), .ZN(_13300_ ) );
NAND3_X1 _20306_ ( .A1(_13299_ ), .A2(_13091_ ), .A3(_13300_ ), .ZN(_13301_ ) );
OAI211_X1 _20307_ ( .A(_13301_ ), .B(_13098_ ), .C1(\wbu.rf_18 [20] ), .C2(_13099_ ), .ZN(_13302_ ) );
NAND4_X1 _20308_ ( .A1(_13106_ ), .A2(_08575_ ), .A3(fanout_net_30 ), .A4(\wbu.rf_19 [20] ), .ZN(_13303_ ) );
NAND3_X1 _20309_ ( .A1(_13302_ ), .A2(_13104_ ), .A3(_13303_ ), .ZN(_13304_ ) );
OAI211_X1 _20310_ ( .A(_13304_ ), .B(_13112_ ), .C1(\wbu.rf_20 [20] ), .C2(_13113_ ), .ZN(_13305_ ) );
NAND4_X1 _20311_ ( .A1(_13120_ ), .A2(_13122_ ), .A3(fanout_net_30 ), .A4(\wbu.rf_21 [20] ), .ZN(_13306_ ) );
NAND3_X1 _20312_ ( .A1(_13305_ ), .A2(_13118_ ), .A3(_13306_ ), .ZN(_13307_ ) );
OAI211_X1 _20313_ ( .A(_13307_ ), .B(_13127_ ), .C1(\wbu.rf_22 [20] ), .C2(_13212_ ), .ZN(_13308_ ) );
NAND4_X1 _20314_ ( .A1(_13133_ ), .A2(fanout_net_30 ), .A3(_13135_ ), .A4(\wbu.rf_23 [20] ), .ZN(_13309_ ) );
NAND3_X1 _20315_ ( .A1(_13308_ ), .A2(_13132_ ), .A3(_13309_ ), .ZN(_13310_ ) );
OAI211_X1 _20316_ ( .A(_13310_ ), .B(_13140_ ), .C1(\wbu.rf_24 [20] ), .C2(_13141_ ), .ZN(_13311_ ) );
BUF_X2 _20317_ ( .A(_13146_ ), .Z(_13312_ ) );
NAND4_X1 _20318_ ( .A1(_13312_ ), .A2(_13149_ ), .A3(fanout_net_30 ), .A4(\wbu.rf_25 [20] ), .ZN(_13313_ ) );
NAND3_X1 _20319_ ( .A1(_13311_ ), .A2(_13145_ ), .A3(_13313_ ), .ZN(_13314_ ) );
OAI211_X1 _20320_ ( .A(_13314_ ), .B(_13218_ ), .C1(\wbu.rf_26 [20] ), .C2(_13154_ ), .ZN(_13315_ ) );
NAND4_X1 _20321_ ( .A1(_13159_ ), .A2(fanout_net_30 ), .A3(_13161_ ), .A4(\wbu.rf_27 [20] ), .ZN(_13316_ ) );
NAND3_X1 _20322_ ( .A1(_13315_ ), .A2(_13157_ ), .A3(_13316_ ), .ZN(_13317_ ) );
OAI211_X1 _20323_ ( .A(_13317_ ), .B(_13165_ ), .C1(\wbu.rf_28 [20] ), .C2(_13167_ ), .ZN(_13318_ ) );
NAND4_X1 _20324_ ( .A1(_13169_ ), .A2(fanout_net_30 ), .A3(_13170_ ), .A4(\wbu.rf_29 [20] ), .ZN(_13319_ ) );
AOI21_X1 _20325_ ( .A(_12975_ ), .B1(_13318_ ), .B2(_13319_ ), .ZN(_13320_ ) );
AND4_X1 _20326_ ( .A1(fanout_net_30 ), .A2(_13175_ ), .A3(\wbu.rf_30 [20] ), .A4(_13176_ ), .ZN(_13321_ ) );
OAI21_X1 _20327_ ( .A(_12971_ ), .B1(_13320_ ), .B2(_13321_ ), .ZN(_13322_ ) );
AOI22_X1 _20328_ ( .A1(_13179_ ), .A2(\wbu.rf_31 [20] ), .B1(_13180_ ), .B2(_13182_ ), .ZN(_13323_ ) );
AOI221_X4 _20329_ ( .A(fanout_net_24 ), .B1(_13279_ ), .B2(_12965_ ), .C1(_13322_ ), .C2(_13323_ ), .ZN(_00349_ ) );
BUF_X4 _20330_ ( .A(_12964_ ), .Z(_13324_ ) );
NAND4_X1 _20331_ ( .A1(_13272_ ), .A2(fanout_net_30 ), .A3(_13273_ ), .A4(\wbu.rf_30 [19] ), .ZN(_13325_ ) );
BUF_X2 _20332_ ( .A(_13147_ ), .Z(_13326_ ) );
BUF_X2 _20333_ ( .A(_13079_ ), .Z(_13327_ ) );
AND4_X1 _20334_ ( .A1(fanout_net_30 ), .A2(_13326_ ), .A3(\wbu.rf_29 [19] ), .A4(_13327_ ), .ZN(_13328_ ) );
NAND4_X1 _20335_ ( .A1(_13146_ ), .A2(_13148_ ), .A3(fanout_net_30 ), .A4(\wbu.rf_25 [19] ), .ZN(_13329_ ) );
NAND4_X1 _20336_ ( .A1(_13121_ ), .A2(fanout_net_30 ), .A3(_13106_ ), .A4(\wbu.rf_23 [19] ), .ZN(_13330_ ) );
NAND4_X1 _20337_ ( .A1(_13173_ ), .A2(fanout_net_37 ), .A3(_13063_ ), .A4(\wbu.rf_14 [19] ), .ZN(_13331_ ) );
AND4_X1 _20338_ ( .A1(fanout_net_37 ), .A2(_12985_ ), .A3(\wbu.rf_13 [19] ), .A4(_13063_ ), .ZN(_13332_ ) );
MUX2_X1 _20339_ ( .A(\wbu._GEN_71 [19] ), .B(\wbu.rf_2 [19] ), .S(_12992_ ), .Z(_13333_ ) );
MUX2_X1 _20340_ ( .A(\wbu.rf_3 [19] ), .B(_13333_ ), .S(_12997_ ), .Z(_13334_ ) );
MUX2_X1 _20341_ ( .A(\wbu.rf_4 [19] ), .B(_13334_ ), .S(_13003_ ), .Z(_13335_ ) );
MUX2_X1 _20342_ ( .A(\wbu.rf_5 [19] ), .B(_13335_ ), .S(_13011_ ), .Z(_13336_ ) );
MUX2_X1 _20343_ ( .A(\wbu.rf_6 [19] ), .B(_13336_ ), .S(_13017_ ), .Z(_13337_ ) );
MUX2_X1 _20344_ ( .A(\wbu.rf_7 [19] ), .B(_13337_ ), .S(_13023_ ), .Z(_13338_ ) );
MUX2_X1 _20345_ ( .A(\wbu.rf_8 [19] ), .B(_13338_ ), .S(_13029_ ), .Z(_13339_ ) );
MUX2_X1 _20346_ ( .A(\wbu.rf_9 [19] ), .B(_13339_ ), .S(_13198_ ), .Z(_13340_ ) );
MUX2_X1 _20347_ ( .A(\wbu.rf_10 [19] ), .B(_13340_ ), .S(_12983_ ), .Z(_13341_ ) );
MUX2_X1 _20348_ ( .A(\wbu.rf_11 [19] ), .B(_13341_ ), .S(_13037_ ), .Z(_13342_ ) );
MUX2_X1 _20349_ ( .A(\wbu.rf_12 [19] ), .B(_13342_ ), .S(_13044_ ), .Z(_13343_ ) );
AOI21_X1 _20350_ ( .A(_13332_ ), .B1(_13343_ ), .B2(_13053_ ), .ZN(_13344_ ) );
OAI211_X1 _20351_ ( .A(_13069_ ), .B(_13331_ ), .C1(_13344_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_13345_ ) );
OAI211_X1 _20352_ ( .A(_13345_ ), .B(_13074_ ), .C1(\wbu.rf_15 [19] ), .C2(_13069_ ), .ZN(_13346_ ) );
NAND4_X1 _20353_ ( .A1(_08573_ ), .A2(_13228_ ), .A3(fanout_net_30 ), .A4(\wbu.rf_16 [19] ), .ZN(_13347_ ) );
NAND3_X1 _20354_ ( .A1(_13346_ ), .A2(_13084_ ), .A3(_13347_ ), .ZN(_13348_ ) );
OAI211_X1 _20355_ ( .A(_13348_ ), .B(_13090_ ), .C1(\wbu.rf_17 [19] ), .C2(_13085_ ), .ZN(_13349_ ) );
BUF_X2 _20356_ ( .A(_08573_ ), .Z(_13350_ ) );
NAND4_X1 _20357_ ( .A1(_13173_ ), .A2(fanout_net_30 ), .A3(\wbu.rf_18 [19] ), .A4(_13350_ ), .ZN(_13351_ ) );
AOI21_X1 _20358_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .B1(_13349_ ), .B2(_13351_ ), .ZN(_13352_ ) );
NAND3_X1 _20359_ ( .A1(_12994_ ), .A2(fanout_net_30 ), .A3(\wbu.rf_19 [19] ), .ZN(_13353_ ) );
NAND2_X1 _20360_ ( .A1(_13102_ ), .A2(_13353_ ), .ZN(_13354_ ) );
OAI221_X1 _20361_ ( .A(_13110_ ), .B1(\wbu.rf_20 [19] ), .B2(_13102_ ), .C1(_13352_ ), .C2(_13354_ ), .ZN(_13355_ ) );
NAND4_X1 _20362_ ( .A1(_13119_ ), .A2(_13121_ ), .A3(fanout_net_30 ), .A4(\wbu.rf_21 [19] ), .ZN(_13356_ ) );
AOI21_X1 _20363_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .B1(_13355_ ), .B2(_13356_ ), .ZN(_13357_ ) );
AOI21_X1 _20364_ ( .A(_13357_ ), .B1(\wbu.rf_22 [19] ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .ZN(_13358_ ) );
OAI211_X1 _20365_ ( .A(_13130_ ), .B(_13330_ ), .C1(_13358_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .ZN(_13359_ ) );
OAI21_X1 _20366_ ( .A(_13359_ ), .B1(\wbu.rf_24 [19] ), .B2(_13131_ ), .ZN(_13360_ ) );
OAI21_X1 _20367_ ( .A(_13329_ ), .B1(_13360_ ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .ZN(_13361_ ) );
MUX2_X1 _20368_ ( .A(\wbu.rf_26 [19] ), .B(_13361_ ), .S(_13143_ ), .Z(_13362_ ) );
BUF_X4 _20369_ ( .A(_13152_ ), .Z(_13363_ ) );
MUX2_X1 _20370_ ( .A(\wbu.rf_27 [19] ), .B(_13362_ ), .S(_13363_ ), .Z(_13364_ ) );
BUF_X4 _20371_ ( .A(_13156_ ), .Z(_13365_ ) );
MUX2_X1 _20372_ ( .A(\wbu.rf_28 [19] ), .B(_13364_ ), .S(_13365_ ), .Z(_13366_ ) );
AOI21_X1 _20373_ ( .A(_13328_ ), .B1(_13366_ ), .B2(_13269_ ), .ZN(_13367_ ) );
OAI211_X1 _20374_ ( .A(_12971_ ), .B(_13325_ ), .C1(_13367_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_13368_ ) );
BUF_X2 _20375_ ( .A(_12970_ ), .Z(_13369_ ) );
OR2_X1 _20376_ ( .A1(_13369_ ), .A2(\wbu.rf_31 [19] ), .ZN(_13370_ ) );
AOI21_X1 _20377_ ( .A(_13324_ ), .B1(_13368_ ), .B2(_13370_ ), .ZN(_13371_ ) );
INV_X1 _20378_ ( .A(\wbu.io_in_bits_rd_wdata [19] ), .ZN(_13372_ ) );
BUF_X4 _20379_ ( .A(_13324_ ), .Z(_13373_ ) );
AOI211_X1 _20380_ ( .A(fanout_net_24 ), .B(_13371_ ), .C1(_13372_ ), .C2(_13373_ ), .ZN(_00350_ ) );
BUF_X2 _20381_ ( .A(_12970_ ), .Z(_13374_ ) );
NAND4_X1 _20382_ ( .A1(_13272_ ), .A2(fanout_net_30 ), .A3(_13273_ ), .A4(\wbu.rf_30 [18] ), .ZN(_13375_ ) );
CLKBUF_X2 _20383_ ( .A(_13079_ ), .Z(_13376_ ) );
AND4_X1 _20384_ ( .A1(fanout_net_30 ), .A2(_13326_ ), .A3(\wbu.rf_29 [18] ), .A4(_13376_ ), .ZN(_13377_ ) );
BUF_X2 _20385_ ( .A(_13148_ ), .Z(_13378_ ) );
NAND4_X1 _20386_ ( .A1(_13174_ ), .A2(_13378_ ), .A3(fanout_net_30 ), .A4(\wbu.rf_26 [18] ), .ZN(_13379_ ) );
AND4_X1 _20387_ ( .A1(fanout_net_30 ), .A2(_13146_ ), .A3(_13148_ ), .A4(\wbu.rf_25 [18] ), .ZN(_13380_ ) );
BUF_X4 _20388_ ( .A(_13103_ ), .Z(_13381_ ) );
OR2_X1 _20389_ ( .A1(_13086_ ), .A2(\wbu.rf_17 [18] ), .ZN(_13382_ ) );
BUF_X4 _20390_ ( .A(_13198_ ), .Z(_13383_ ) );
OR2_X1 _20391_ ( .A1(_13030_ ), .A2(\wbu.rf_8 [18] ), .ZN(_13384_ ) );
MUX2_X1 _20392_ ( .A(\wbu._GEN_71 [18] ), .B(\wbu.rf_2 [18] ), .S(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .Z(_13385_ ) );
MUX2_X1 _20393_ ( .A(\wbu.rf_3 [18] ), .B(_13385_ ), .S(_12998_ ), .Z(_13386_ ) );
MUX2_X1 _20394_ ( .A(\wbu.rf_4 [18] ), .B(_13386_ ), .S(_13004_ ), .Z(_13387_ ) );
MUX2_X1 _20395_ ( .A(\wbu.rf_5 [18] ), .B(_13387_ ), .S(_13012_ ), .Z(_13388_ ) );
MUX2_X1 _20396_ ( .A(\wbu.rf_6 [18] ), .B(_13388_ ), .S(_13018_ ), .Z(_13389_ ) );
MUX2_X1 _20397_ ( .A(\wbu.rf_7 [18] ), .B(_13389_ ), .S(_13024_ ), .Z(_13390_ ) );
OAI211_X1 _20398_ ( .A(_13383_ ), .B(_13384_ ), .C1(_13390_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_Y ), .ZN(_13391_ ) );
NAND4_X1 _20399_ ( .A1(_12985_ ), .A2(_13046_ ), .A3(fanout_net_37 ), .A4(\wbu.rf_9 [18] ), .ZN(_13392_ ) );
NAND3_X1 _20400_ ( .A1(_13391_ ), .A2(_13039_ ), .A3(_13392_ ), .ZN(_13393_ ) );
OAI211_X1 _20401_ ( .A(_13393_ ), .B(_13038_ ), .C1(\wbu.rf_10 [18] ), .C2(_13039_ ), .ZN(_13394_ ) );
NAND4_X1 _20402_ ( .A1(_13148_ ), .A2(fanout_net_37 ), .A3(_13047_ ), .A4(\wbu.rf_11 [18] ), .ZN(_13395_ ) );
NAND3_X1 _20403_ ( .A1(_13394_ ), .A2(_13045_ ), .A3(_13395_ ), .ZN(_13396_ ) );
OAI211_X1 _20404_ ( .A(_13396_ ), .B(_13054_ ), .C1(\wbu.rf_12 [18] ), .C2(_13055_ ), .ZN(_13397_ ) );
NAND4_X1 _20405_ ( .A1(_13062_ ), .A2(fanout_net_37 ), .A3(_13078_ ), .A4(\wbu.rf_13 [18] ), .ZN(_13398_ ) );
NAND3_X1 _20406_ ( .A1(_13397_ ), .A2(_13060_ ), .A3(_13398_ ), .ZN(_13399_ ) );
OAI211_X1 _20407_ ( .A(_13399_ ), .B(_13070_ ), .C1(\wbu.rf_14 [18] ), .C2(_13071_ ), .ZN(_13400_ ) );
NAND4_X1 _20408_ ( .A1(_13077_ ), .A2(_13079_ ), .A3(fanout_net_38 ), .A4(\wbu.rf_15 [18] ), .ZN(_13401_ ) );
NAND2_X1 _20409_ ( .A1(_13400_ ), .A2(_13401_ ), .ZN(_13402_ ) );
MUX2_X1 _20410_ ( .A(\wbu.rf_16 [18] ), .B(_13402_ ), .S(_13076_ ), .Z(_13403_ ) );
OAI211_X1 _20411_ ( .A(_13099_ ), .B(_13382_ ), .C1(_13403_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_13404_ ) );
NAND4_X1 _20412_ ( .A1(_13174_ ), .A2(fanout_net_30 ), .A3(\wbu.rf_18 [18] ), .A4(_08575_ ), .ZN(_13405_ ) );
AOI21_X1 _20413_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .B1(_13404_ ), .B2(_13405_ ), .ZN(_13406_ ) );
NAND3_X1 _20414_ ( .A1(_12994_ ), .A2(fanout_net_30 ), .A3(\wbu.rf_19 [18] ), .ZN(_13407_ ) );
NAND2_X1 _20415_ ( .A1(_13381_ ), .A2(_13407_ ), .ZN(_13408_ ) );
OAI221_X1 _20416_ ( .A(_13112_ ), .B1(\wbu.rf_20 [18] ), .B2(_13381_ ), .C1(_13406_ ), .C2(_13408_ ), .ZN(_13409_ ) );
NAND4_X1 _20417_ ( .A1(_13120_ ), .A2(_13122_ ), .A3(fanout_net_30 ), .A4(\wbu.rf_21 [18] ), .ZN(_13410_ ) );
NAND3_X1 _20418_ ( .A1(_13409_ ), .A2(_13212_ ), .A3(_13410_ ), .ZN(_13411_ ) );
OR2_X1 _20419_ ( .A1(_13117_ ), .A2(\wbu.rf_22 [18] ), .ZN(_13412_ ) );
NAND3_X1 _20420_ ( .A1(_13411_ ), .A2(_13231_ ), .A3(_13412_ ), .ZN(_13413_ ) );
BUF_X4 _20421_ ( .A(_13131_ ), .Z(_13414_ ) );
NAND3_X1 _20422_ ( .A1(_13020_ ), .A2(fanout_net_31 ), .A3(\wbu.rf_23 [18] ), .ZN(_13415_ ) );
NAND3_X1 _20423_ ( .A1(_13413_ ), .A2(_13414_ ), .A3(_13415_ ), .ZN(_13416_ ) );
NOR2_X1 _20424_ ( .A1(_13131_ ), .A2(\wbu.rf_24 [18] ), .ZN(_13417_ ) );
NOR2_X1 _20425_ ( .A1(_13417_ ), .A2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .ZN(_13418_ ) );
AOI21_X1 _20426_ ( .A(_13380_ ), .B1(_13416_ ), .B2(_13418_ ), .ZN(_13419_ ) );
OAI21_X1 _20427_ ( .A(_13379_ ), .B1(_13419_ ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_13420_ ) );
MUX2_X1 _20428_ ( .A(\wbu.rf_27 [18] ), .B(_13420_ ), .S(_13218_ ), .Z(_13421_ ) );
MUX2_X1 _20429_ ( .A(\wbu.rf_28 [18] ), .B(_13421_ ), .S(_13365_ ), .Z(_13422_ ) );
AOI21_X1 _20430_ ( .A(_13377_ ), .B1(_13422_ ), .B2(_13269_ ), .ZN(_13423_ ) );
OAI211_X1 _20431_ ( .A(_13374_ ), .B(_13375_ ), .C1(_13423_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_13424_ ) );
OAI211_X1 _20432_ ( .A(_13424_ ), .B(_13276_ ), .C1(\wbu.rf_31 [18] ), .C2(_13271_ ), .ZN(_13425_ ) );
NAND3_X1 _20433_ ( .A1(_13181_ ), .A2(\wbu.io_in_bits_rd_wdata [18] ), .A3(_13183_ ), .ZN(_13426_ ) );
AOI21_X1 _20434_ ( .A(fanout_net_24 ), .B1(_13425_ ), .B2(_13426_ ), .ZN(_00351_ ) );
INV_X1 _20435_ ( .A(\wbu.io_in_bits_rd_wdata [17] ), .ZN(_13427_ ) );
NAND4_X1 _20436_ ( .A1(_12985_ ), .A2(_12986_ ), .A3(fanout_net_38 ), .A4(\wbu.rf_9 [17] ), .ZN(_13428_ ) );
AND4_X1 _20437_ ( .A1(fanout_net_38 ), .A2(_12986_ ), .A3(\wbu.rf_8 [17] ), .A4(_12960_ ), .ZN(_13429_ ) );
MUX2_X1 _20438_ ( .A(\wbu._GEN_71 [17] ), .B(\wbu.rf_2 [17] ), .S(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .Z(_13430_ ) );
MUX2_X1 _20439_ ( .A(\wbu.rf_3 [17] ), .B(_13430_ ), .S(_12998_ ), .Z(_13431_ ) );
MUX2_X1 _20440_ ( .A(\wbu.rf_4 [17] ), .B(_13431_ ), .S(_13004_ ), .Z(_13432_ ) );
MUX2_X1 _20441_ ( .A(\wbu.rf_5 [17] ), .B(_13432_ ), .S(_13012_ ), .Z(_13433_ ) );
MUX2_X1 _20442_ ( .A(\wbu.rf_6 [17] ), .B(_13433_ ), .S(_13018_ ), .Z(_13434_ ) );
MUX2_X1 _20443_ ( .A(\wbu.rf_7 [17] ), .B(_13434_ ), .S(_13024_ ), .Z(_13435_ ) );
AOI21_X1 _20444_ ( .A(_13429_ ), .B1(_13435_ ), .B2(_13030_ ), .ZN(_13436_ ) );
OAI211_X1 _20445_ ( .A(_12984_ ), .B(_13428_ ), .C1(_13436_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_Y ), .ZN(_13437_ ) );
OAI211_X1 _20446_ ( .A(_13437_ ), .B(_13038_ ), .C1(\wbu.rf_10 [17] ), .C2(_13039_ ), .ZN(_13438_ ) );
NAND4_X1 _20447_ ( .A1(_13046_ ), .A2(fanout_net_38 ), .A3(_13047_ ), .A4(\wbu.rf_11 [17] ), .ZN(_13439_ ) );
NAND3_X1 _20448_ ( .A1(_13438_ ), .A2(_13045_ ), .A3(_13439_ ), .ZN(_13440_ ) );
OAI211_X1 _20449_ ( .A(_13440_ ), .B(_13054_ ), .C1(\wbu.rf_12 [17] ), .C2(_13055_ ), .ZN(_13441_ ) );
NAND4_X1 _20450_ ( .A1(_13062_ ), .A2(fanout_net_38 ), .A3(_13064_ ), .A4(\wbu.rf_13 [17] ), .ZN(_13442_ ) );
NAND3_X1 _20451_ ( .A1(_13441_ ), .A2(_13060_ ), .A3(_13442_ ), .ZN(_13443_ ) );
OAI211_X1 _20452_ ( .A(_13443_ ), .B(_13070_ ), .C1(\wbu.rf_14 [17] ), .C2(_13071_ ), .ZN(_13444_ ) );
NAND4_X1 _20453_ ( .A1(_13077_ ), .A2(_13078_ ), .A3(fanout_net_38 ), .A4(\wbu.rf_15 [17] ), .ZN(_13445_ ) );
NAND3_X1 _20454_ ( .A1(_13444_ ), .A2(_13076_ ), .A3(_13445_ ), .ZN(_13446_ ) );
OAI211_X1 _20455_ ( .A(_13446_ ), .B(_13086_ ), .C1(\wbu.rf_16 [17] ), .C2(_13087_ ), .ZN(_13447_ ) );
NAND4_X1 _20456_ ( .A1(_13092_ ), .A2(fanout_net_31 ), .A3(\wbu.rf_17 [17] ), .A4(_08574_ ), .ZN(_13448_ ) );
NAND3_X1 _20457_ ( .A1(_13447_ ), .A2(_13091_ ), .A3(_13448_ ), .ZN(_13449_ ) );
BUF_X4 _20458_ ( .A(_13090_ ), .Z(_13450_ ) );
OAI211_X1 _20459_ ( .A(_13449_ ), .B(_13098_ ), .C1(\wbu.rf_18 [17] ), .C2(_13450_ ), .ZN(_13451_ ) );
NAND4_X1 _20460_ ( .A1(_13106_ ), .A2(_08575_ ), .A3(fanout_net_31 ), .A4(\wbu.rf_19 [17] ), .ZN(_13452_ ) );
NAND3_X1 _20461_ ( .A1(_13451_ ), .A2(_13104_ ), .A3(_13452_ ), .ZN(_13453_ ) );
OAI211_X1 _20462_ ( .A(_13453_ ), .B(_13112_ ), .C1(\wbu.rf_20 [17] ), .C2(_13381_ ), .ZN(_13454_ ) );
NAND4_X1 _20463_ ( .A1(_13120_ ), .A2(_13188_ ), .A3(fanout_net_31 ), .A4(\wbu.rf_21 [17] ), .ZN(_13455_ ) );
NAND3_X1 _20464_ ( .A1(_13454_ ), .A2(_13118_ ), .A3(_13455_ ), .ZN(_13456_ ) );
OAI211_X1 _20465_ ( .A(_13456_ ), .B(_13127_ ), .C1(\wbu.rf_22 [17] ), .C2(_13212_ ), .ZN(_13457_ ) );
NAND4_X1 _20466_ ( .A1(_13133_ ), .A2(fanout_net_31 ), .A3(_13135_ ), .A4(\wbu.rf_23 [17] ), .ZN(_13458_ ) );
NAND3_X1 _20467_ ( .A1(_13457_ ), .A2(_13132_ ), .A3(_13458_ ), .ZN(_13459_ ) );
BUF_X4 _20468_ ( .A(_13139_ ), .Z(_13460_ ) );
OAI211_X1 _20469_ ( .A(_13459_ ), .B(_13460_ ), .C1(\wbu.rf_24 [17] ), .C2(_13141_ ), .ZN(_13461_ ) );
NAND4_X1 _20470_ ( .A1(_13312_ ), .A2(_13149_ ), .A3(fanout_net_31 ), .A4(\wbu.rf_25 [17] ), .ZN(_13462_ ) );
NAND3_X1 _20471_ ( .A1(_13461_ ), .A2(_13145_ ), .A3(_13462_ ), .ZN(_13463_ ) );
OAI211_X1 _20472_ ( .A(_13463_ ), .B(_13218_ ), .C1(\wbu.rf_26 [17] ), .C2(_13154_ ), .ZN(_13464_ ) );
NAND4_X1 _20473_ ( .A1(_13159_ ), .A2(fanout_net_31 ), .A3(_13161_ ), .A4(\wbu.rf_27 [17] ), .ZN(_13465_ ) );
NAND3_X1 _20474_ ( .A1(_13464_ ), .A2(_13157_ ), .A3(_13465_ ), .ZN(_13466_ ) );
OAI211_X1 _20475_ ( .A(_13466_ ), .B(_13165_ ), .C1(\wbu.rf_28 [17] ), .C2(_13167_ ), .ZN(_13467_ ) );
NAND4_X1 _20476_ ( .A1(_13169_ ), .A2(fanout_net_31 ), .A3(_13170_ ), .A4(\wbu.rf_29 [17] ), .ZN(_13468_ ) );
AOI21_X1 _20477_ ( .A(_12975_ ), .B1(_13467_ ), .B2(_13468_ ), .ZN(_13469_ ) );
AND4_X1 _20478_ ( .A1(fanout_net_31 ), .A2(_13175_ ), .A3(\wbu.rf_30 [17] ), .A4(_13176_ ), .ZN(_13470_ ) );
OAI21_X1 _20479_ ( .A(_12971_ ), .B1(_13469_ ), .B2(_13470_ ), .ZN(_13471_ ) );
AOI22_X1 _20480_ ( .A1(_13179_ ), .A2(\wbu.rf_31 [17] ), .B1(_13180_ ), .B2(_13182_ ), .ZN(_13472_ ) );
AOI221_X4 _20481_ ( .A(fanout_net_24 ), .B1(_13427_ ), .B2(_12965_ ), .C1(_13471_ ), .C2(_13472_ ), .ZN(_00352_ ) );
BUF_X4 _20482_ ( .A(_12964_ ), .Z(_13473_ ) );
CLKBUF_X2 _20483_ ( .A(_12968_ ), .Z(_13474_ ) );
AND3_X1 _20484_ ( .A1(_13474_ ), .A2(fanout_net_31 ), .A3(\wbu.rf_31 [16] ), .ZN(_13475_ ) );
NAND4_X1 _20485_ ( .A1(_13061_ ), .A2(fanout_net_38 ), .A3(_13064_ ), .A4(\wbu.rf_13 [16] ), .ZN(_13476_ ) );
AND4_X1 _20486_ ( .A1(fanout_net_38 ), .A2(_13063_ ), .A3(\wbu.rf_12 [16] ), .A4(_12960_ ), .ZN(_13477_ ) );
MUX2_X1 _20487_ ( .A(\wbu._GEN_71 [16] ), .B(\wbu.rf_2 [16] ), .S(_12992_ ), .Z(_13478_ ) );
MUX2_X1 _20488_ ( .A(\wbu.rf_3 [16] ), .B(_13478_ ), .S(_12997_ ), .Z(_13479_ ) );
MUX2_X1 _20489_ ( .A(\wbu.rf_4 [16] ), .B(_13479_ ), .S(_13003_ ), .Z(_13480_ ) );
MUX2_X1 _20490_ ( .A(\wbu.rf_5 [16] ), .B(_13480_ ), .S(_13011_ ), .Z(_13481_ ) );
MUX2_X1 _20491_ ( .A(\wbu.rf_6 [16] ), .B(_13481_ ), .S(_13017_ ), .Z(_13482_ ) );
MUX2_X1 _20492_ ( .A(\wbu.rf_7 [16] ), .B(_13482_ ), .S(_13023_ ), .Z(_13483_ ) );
MUX2_X1 _20493_ ( .A(\wbu.rf_8 [16] ), .B(_13483_ ), .S(_13029_ ), .Z(_13484_ ) );
MUX2_X1 _20494_ ( .A(\wbu.rf_9 [16] ), .B(_13484_ ), .S(_13383_ ), .Z(_13485_ ) );
MUX2_X1 _20495_ ( .A(\wbu.rf_10 [16] ), .B(_13485_ ), .S(_12984_ ), .Z(_13486_ ) );
MUX2_X1 _20496_ ( .A(\wbu.rf_11 [16] ), .B(_13486_ ), .S(_13038_ ), .Z(_13487_ ) );
AOI21_X1 _20497_ ( .A(_13477_ ), .B1(_13487_ ), .B2(_13045_ ), .ZN(_13488_ ) );
OAI211_X1 _20498_ ( .A(_13059_ ), .B(_13476_ ), .C1(_13488_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_13489_ ) );
OAI211_X1 _20499_ ( .A(_13489_ ), .B(_13070_ ), .C1(\wbu.rf_14 [16] ), .C2(_13060_ ), .ZN(_13490_ ) );
NAND4_X1 _20500_ ( .A1(_13047_ ), .A2(_13078_ ), .A3(fanout_net_38 ), .A4(\wbu.rf_15 [16] ), .ZN(_13491_ ) );
NAND3_X1 _20501_ ( .A1(_13490_ ), .A2(_13075_ ), .A3(_13491_ ), .ZN(_13492_ ) );
OAI211_X1 _20502_ ( .A(_13492_ ), .B(_13085_ ), .C1(\wbu.rf_16 [16] ), .C2(_13076_ ), .ZN(_13493_ ) );
NAND4_X1 _20503_ ( .A1(_13092_ ), .A2(fanout_net_31 ), .A3(\wbu.rf_17 [16] ), .A4(_13350_ ), .ZN(_13494_ ) );
NAND3_X1 _20504_ ( .A1(_13493_ ), .A2(_13091_ ), .A3(_13494_ ), .ZN(_13495_ ) );
OAI211_X1 _20505_ ( .A(_13495_ ), .B(_13097_ ), .C1(\wbu.rf_18 [16] ), .C2(_13450_ ), .ZN(_13496_ ) );
BUF_X2 _20506_ ( .A(_13350_ ), .Z(_13497_ ) );
NAND4_X1 _20507_ ( .A1(_13105_ ), .A2(_13497_ ), .A3(fanout_net_31 ), .A4(\wbu.rf_19 [16] ), .ZN(_13498_ ) );
NAND3_X1 _20508_ ( .A1(_13496_ ), .A2(_13103_ ), .A3(_13498_ ), .ZN(_13499_ ) );
OAI211_X1 _20509_ ( .A(_13499_ ), .B(_13111_ ), .C1(\wbu.rf_20 [16] ), .C2(_13104_ ), .ZN(_13500_ ) );
NAND4_X1 _20510_ ( .A1(_13119_ ), .A2(_13121_ ), .A3(fanout_net_31 ), .A4(\wbu.rf_21 [16] ), .ZN(_13501_ ) );
NAND3_X1 _20511_ ( .A1(_13500_ ), .A2(_13117_ ), .A3(_13501_ ), .ZN(_13502_ ) );
OAI211_X1 _20512_ ( .A(_13502_ ), .B(_13127_ ), .C1(\wbu.rf_22 [16] ), .C2(_13118_ ), .ZN(_13503_ ) );
NAND4_X1 _20513_ ( .A1(_13186_ ), .A2(fanout_net_31 ), .A3(_13134_ ), .A4(\wbu.rf_23 [16] ), .ZN(_13504_ ) );
NAND3_X1 _20514_ ( .A1(_13503_ ), .A2(_13131_ ), .A3(_13504_ ), .ZN(_13505_ ) );
OAI211_X1 _20515_ ( .A(_13505_ ), .B(_13460_ ), .C1(\wbu.rf_24 [16] ), .C2(_13414_ ), .ZN(_13506_ ) );
NAND4_X1 _20516_ ( .A1(_13146_ ), .A2(_13378_ ), .A3(fanout_net_31 ), .A4(\wbu.rf_25 [16] ), .ZN(_13507_ ) );
NAND3_X1 _20517_ ( .A1(_13506_ ), .A2(_13144_ ), .A3(_13507_ ), .ZN(_13508_ ) );
OAI211_X1 _20518_ ( .A(_13508_ ), .B(_13363_ ), .C1(\wbu.rf_26 [16] ), .C2(_13260_ ), .ZN(_13509_ ) );
NAND4_X1 _20519_ ( .A1(_13158_ ), .A2(fanout_net_31 ), .A3(_13160_ ), .A4(\wbu.rf_27 [16] ), .ZN(_13510_ ) );
NAND3_X1 _20520_ ( .A1(_13509_ ), .A2(_13166_ ), .A3(_13510_ ), .ZN(_13511_ ) );
BUF_X4 _20521_ ( .A(_13164_ ), .Z(_13512_ ) );
OAI211_X1 _20522_ ( .A(_13511_ ), .B(_13512_ ), .C1(\wbu.rf_28 [16] ), .C2(_13365_ ), .ZN(_13513_ ) );
NAND4_X1 _20523_ ( .A1(_13326_ ), .A2(fanout_net_31 ), .A3(_13327_ ), .A4(\wbu.rf_29 [16] ), .ZN(_13514_ ) );
NAND2_X1 _20524_ ( .A1(_13513_ ), .A2(_13514_ ), .ZN(_13515_ ) );
MUX2_X1 _20525_ ( .A(\wbu.rf_30 [16] ), .B(_13515_ ), .S(_13268_ ), .Z(_13516_ ) );
AOI211_X1 _20526_ ( .A(_13473_ ), .B(_13475_ ), .C1(_13516_ ), .C2(_13271_ ), .ZN(_13517_ ) );
INV_X1 _20527_ ( .A(\wbu.io_in_bits_rd_wdata [16] ), .ZN(_13518_ ) );
AOI211_X1 _20528_ ( .A(fanout_net_24 ), .B(_13517_ ), .C1(_13518_ ), .C2(_13373_ ), .ZN(_00353_ ) );
INV_X1 _20529_ ( .A(\wbu.io_in_bits_rd_wdata [15] ), .ZN(_13519_ ) );
NAND4_X1 _20530_ ( .A1(_13312_ ), .A2(_13378_ ), .A3(fanout_net_31 ), .A4(\wbu.rf_25 [15] ), .ZN(_13520_ ) );
AND4_X1 _20531_ ( .A1(fanout_net_31 ), .A2(_13148_ ), .A3(\wbu.rf_24 [15] ), .A4(_13229_ ), .ZN(_13521_ ) );
MUX2_X1 _20532_ ( .A(\wbu._GEN_71 [15] ), .B(\wbu.rf_2 [15] ), .S(_12990_ ), .Z(_13522_ ) );
MUX2_X1 _20533_ ( .A(\wbu.rf_3 [15] ), .B(_13522_ ), .S(_12995_ ), .Z(_13523_ ) );
MUX2_X1 _20534_ ( .A(\wbu.rf_4 [15] ), .B(_13523_ ), .S(_13001_ ), .Z(_13524_ ) );
MUX2_X1 _20535_ ( .A(\wbu.rf_5 [15] ), .B(_13524_ ), .S(_13009_ ), .Z(_13525_ ) );
MUX2_X1 _20536_ ( .A(\wbu.rf_6 [15] ), .B(_13525_ ), .S(_13015_ ), .Z(_13526_ ) );
MUX2_X1 _20537_ ( .A(\wbu.rf_7 [15] ), .B(_13526_ ), .S(_13021_ ), .Z(_13527_ ) );
MUX2_X1 _20538_ ( .A(\wbu.rf_8 [15] ), .B(_13527_ ), .S(_13027_ ), .Z(_13528_ ) );
MUX2_X1 _20539_ ( .A(\wbu.rf_9 [15] ), .B(_13528_ ), .S(_13197_ ), .Z(_13529_ ) );
MUX2_X1 _20540_ ( .A(\wbu.rf_10 [15] ), .B(_13529_ ), .S(_12982_ ), .Z(_13530_ ) );
MUX2_X1 _20541_ ( .A(\wbu.rf_11 [15] ), .B(_13530_ ), .S(_13036_ ), .Z(_13531_ ) );
MUX2_X1 _20542_ ( .A(\wbu.rf_12 [15] ), .B(_13531_ ), .S(_13043_ ), .Z(_13532_ ) );
MUX2_X1 _20543_ ( .A(\wbu.rf_13 [15] ), .B(_13532_ ), .S(_13052_ ), .Z(_13533_ ) );
MUX2_X1 _20544_ ( .A(\wbu.rf_14 [15] ), .B(_13533_ ), .S(_13057_ ), .Z(_13534_ ) );
MUX2_X1 _20545_ ( .A(\wbu.rf_15 [15] ), .B(_13534_ ), .S(_13068_ ), .Z(_13535_ ) );
MUX2_X1 _20546_ ( .A(\wbu.rf_16 [15] ), .B(_13535_ ), .S(_13074_ ), .Z(_13536_ ) );
MUX2_X1 _20547_ ( .A(\wbu.rf_17 [15] ), .B(_13536_ ), .S(_13084_ ), .Z(_13537_ ) );
MUX2_X1 _20548_ ( .A(\wbu.rf_18 [15] ), .B(_13537_ ), .S(_13090_ ), .Z(_13538_ ) );
MUX2_X1 _20549_ ( .A(\wbu.rf_19 [15] ), .B(_13538_ ), .S(_13097_ ), .Z(_13539_ ) );
MUX2_X1 _20550_ ( .A(\wbu.rf_20 [15] ), .B(_13539_ ), .S(_13102_ ), .Z(_13540_ ) );
MUX2_X1 _20551_ ( .A(\wbu.rf_21 [15] ), .B(_13540_ ), .S(_13110_ ), .Z(_13541_ ) );
MUX2_X1 _20552_ ( .A(\wbu.rf_22 [15] ), .B(_13541_ ), .S(_13116_ ), .Z(_13542_ ) );
MUX2_X1 _20553_ ( .A(\wbu.rf_23 [15] ), .B(_13542_ ), .S(_13127_ ), .Z(_13543_ ) );
AOI21_X1 _20554_ ( .A(_13521_ ), .B1(_13543_ ), .B2(_13414_ ), .ZN(_13544_ ) );
OAI211_X1 _20555_ ( .A(_13144_ ), .B(_13520_ ), .C1(_13544_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .ZN(_13545_ ) );
OAI211_X1 _20556_ ( .A(_13545_ ), .B(_13218_ ), .C1(\wbu.rf_26 [15] ), .C2(_13154_ ), .ZN(_13546_ ) );
NAND4_X1 _20557_ ( .A1(_13159_ ), .A2(fanout_net_31 ), .A3(_13161_ ), .A4(\wbu.rf_27 [15] ), .ZN(_13547_ ) );
NAND3_X1 _20558_ ( .A1(_13546_ ), .A2(_13157_ ), .A3(_13547_ ), .ZN(_13548_ ) );
OAI211_X1 _20559_ ( .A(_13548_ ), .B(_13512_ ), .C1(\wbu.rf_28 [15] ), .C2(_13167_ ), .ZN(_13549_ ) );
NAND4_X1 _20560_ ( .A1(_13169_ ), .A2(fanout_net_31 ), .A3(_13176_ ), .A4(\wbu.rf_29 [15] ), .ZN(_13550_ ) );
AOI21_X1 _20561_ ( .A(_12975_ ), .B1(_13549_ ), .B2(_13550_ ), .ZN(_13551_ ) );
AND4_X1 _20562_ ( .A1(fanout_net_31 ), .A2(_13175_ ), .A3(\wbu.rf_30 [15] ), .A4(_13376_ ), .ZN(_13552_ ) );
OAI21_X1 _20563_ ( .A(_12971_ ), .B1(_13551_ ), .B2(_13552_ ), .ZN(_13553_ ) );
AOI22_X1 _20564_ ( .A1(_13179_ ), .A2(\wbu.rf_31 [15] ), .B1(_13180_ ), .B2(_13182_ ), .ZN(_13554_ ) );
AOI221_X4 _20565_ ( .A(fanout_net_24 ), .B1(_13519_ ), .B2(_12965_ ), .C1(_13553_ ), .C2(_13554_ ), .ZN(_00354_ ) );
NAND4_X1 _20566_ ( .A1(_13272_ ), .A2(fanout_net_31 ), .A3(_13273_ ), .A4(\wbu.rf_30 [14] ), .ZN(_13555_ ) );
AND4_X1 _20567_ ( .A1(fanout_net_31 ), .A2(_13147_ ), .A3(\wbu.rf_29 [14] ), .A4(_13327_ ), .ZN(_13556_ ) );
NAND3_X1 _20568_ ( .A1(_13000_ ), .A2(fanout_net_31 ), .A3(\wbu.rf_20 [14] ), .ZN(_13557_ ) );
NAND4_X1 _20569_ ( .A1(_13061_ ), .A2(fanout_net_31 ), .A3(\wbu.rf_17 [14] ), .A4(_08573_ ), .ZN(_13558_ ) );
AND4_X1 _20570_ ( .A1(fanout_net_31 ), .A2(_08573_ ), .A3(_12960_ ), .A4(\wbu.rf_16 [14] ), .ZN(_13559_ ) );
MUX2_X1 _20571_ ( .A(\wbu._GEN_71 [14] ), .B(\wbu.rf_2 [14] ), .S(_12991_ ), .Z(_13560_ ) );
MUX2_X1 _20572_ ( .A(\wbu.rf_3 [14] ), .B(_13560_ ), .S(_12996_ ), .Z(_13561_ ) );
MUX2_X1 _20573_ ( .A(\wbu.rf_4 [14] ), .B(_13561_ ), .S(_13002_ ), .Z(_13562_ ) );
MUX2_X1 _20574_ ( .A(\wbu.rf_5 [14] ), .B(_13562_ ), .S(_13010_ ), .Z(_13563_ ) );
MUX2_X1 _20575_ ( .A(\wbu.rf_6 [14] ), .B(_13563_ ), .S(_13016_ ), .Z(_13564_ ) );
MUX2_X1 _20576_ ( .A(\wbu.rf_7 [14] ), .B(_13564_ ), .S(_13022_ ), .Z(_13565_ ) );
MUX2_X1 _20577_ ( .A(\wbu.rf_8 [14] ), .B(_13565_ ), .S(_13028_ ), .Z(_13566_ ) );
MUX2_X1 _20578_ ( .A(\wbu.rf_9 [14] ), .B(_13566_ ), .S(_13197_ ), .Z(_13567_ ) );
MUX2_X1 _20579_ ( .A(\wbu.rf_10 [14] ), .B(_13567_ ), .S(_12982_ ), .Z(_13568_ ) );
MUX2_X1 _20580_ ( .A(\wbu.rf_11 [14] ), .B(_13568_ ), .S(_13036_ ), .Z(_13569_ ) );
MUX2_X1 _20581_ ( .A(\wbu.rf_12 [14] ), .B(_13569_ ), .S(_13043_ ), .Z(_13570_ ) );
MUX2_X1 _20582_ ( .A(\wbu.rf_13 [14] ), .B(_13570_ ), .S(_13052_ ), .Z(_13571_ ) );
MUX2_X1 _20583_ ( .A(\wbu.rf_14 [14] ), .B(_13571_ ), .S(_13058_ ), .Z(_13572_ ) );
MUX2_X1 _20584_ ( .A(\wbu.rf_15 [14] ), .B(_13572_ ), .S(_13068_ ), .Z(_13573_ ) );
AOI21_X1 _20585_ ( .A(_13559_ ), .B1(_13573_ ), .B2(_13074_ ), .ZN(_13574_ ) );
OAI211_X1 _20586_ ( .A(_13090_ ), .B(_13558_ ), .C1(_13574_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_13575_ ) );
OR2_X1 _20587_ ( .A1(_13089_ ), .A2(\wbu.rf_18 [14] ), .ZN(_13576_ ) );
AOI21_X1 _20588_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .B1(_13575_ ), .B2(_13576_ ), .ZN(_13577_ ) );
OAI21_X1 _20589_ ( .A(_13102_ ), .B1(_13096_ ), .B2(\wbu.rf_19 [14] ), .ZN(_13578_ ) );
OAI21_X1 _20590_ ( .A(_13557_ ), .B1(_13577_ ), .B2(_13578_ ), .ZN(_13579_ ) );
MUX2_X1 _20591_ ( .A(\wbu.rf_21 [14] ), .B(_13579_ ), .S(_13110_ ), .Z(_13580_ ) );
MUX2_X1 _20592_ ( .A(\wbu.rf_22 [14] ), .B(_13580_ ), .S(_13116_ ), .Z(_13581_ ) );
MUX2_X1 _20593_ ( .A(\wbu.rf_23 [14] ), .B(_13581_ ), .S(_13126_ ), .Z(_13582_ ) );
MUX2_X1 _20594_ ( .A(\wbu.rf_24 [14] ), .B(_13582_ ), .S(_13130_ ), .Z(_13583_ ) );
MUX2_X1 _20595_ ( .A(\wbu.rf_25 [14] ), .B(_13583_ ), .S(_13139_ ), .Z(_13584_ ) );
MUX2_X1 _20596_ ( .A(\wbu.rf_26 [14] ), .B(_13584_ ), .S(_13143_ ), .Z(_13585_ ) );
MUX2_X1 _20597_ ( .A(\wbu.rf_27 [14] ), .B(_13585_ ), .S(_13363_ ), .Z(_13586_ ) );
MUX2_X1 _20598_ ( .A(\wbu.rf_28 [14] ), .B(_13586_ ), .S(_13157_ ), .Z(_13587_ ) );
AOI21_X1 _20599_ ( .A(_13556_ ), .B1(_13587_ ), .B2(_13269_ ), .ZN(_13588_ ) );
OAI211_X1 _20600_ ( .A(_12971_ ), .B(_13555_ ), .C1(_13588_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_13589_ ) );
OR2_X1 _20601_ ( .A1(_13369_ ), .A2(\wbu.rf_31 [14] ), .ZN(_13590_ ) );
AOI21_X1 _20602_ ( .A(_13324_ ), .B1(_13589_ ), .B2(_13590_ ), .ZN(_13591_ ) );
INV_X1 _20603_ ( .A(\wbu.io_in_bits_rd_wdata [14] ), .ZN(_13592_ ) );
AOI211_X1 _20604_ ( .A(fanout_net_24 ), .B(_13591_ ), .C1(_13592_ ), .C2(_13373_ ), .ZN(_00355_ ) );
AND3_X1 _20605_ ( .A1(_13474_ ), .A2(fanout_net_31 ), .A3(\wbu.rf_31 [13] ), .ZN(_13593_ ) );
NAND4_X1 _20606_ ( .A1(_12966_ ), .A2(_13063_ ), .A3(fanout_net_38 ), .A4(\wbu.rf_15 [13] ), .ZN(_13594_ ) );
AND4_X1 _20607_ ( .A1(fanout_net_38 ), .A2(_12977_ ), .A3(\wbu.rf_14 [13] ), .A4(_13063_ ), .ZN(_13595_ ) );
MUX2_X1 _20608_ ( .A(\wbu._GEN_71 [13] ), .B(\wbu.rf_2 [13] ), .S(_12991_ ), .Z(_13596_ ) );
MUX2_X1 _20609_ ( .A(\wbu.rf_3 [13] ), .B(_13596_ ), .S(_12996_ ), .Z(_13597_ ) );
MUX2_X1 _20610_ ( .A(\wbu.rf_4 [13] ), .B(_13597_ ), .S(_13002_ ), .Z(_13598_ ) );
MUX2_X1 _20611_ ( .A(\wbu.rf_5 [13] ), .B(_13598_ ), .S(_13010_ ), .Z(_13599_ ) );
MUX2_X1 _20612_ ( .A(\wbu.rf_6 [13] ), .B(_13599_ ), .S(_13016_ ), .Z(_13600_ ) );
MUX2_X1 _20613_ ( .A(\wbu.rf_7 [13] ), .B(_13600_ ), .S(_13022_ ), .Z(_13601_ ) );
MUX2_X1 _20614_ ( .A(\wbu.rf_8 [13] ), .B(_13601_ ), .S(_13028_ ), .Z(_13602_ ) );
MUX2_X1 _20615_ ( .A(\wbu.rf_9 [13] ), .B(_13602_ ), .S(_13197_ ), .Z(_13603_ ) );
MUX2_X1 _20616_ ( .A(\wbu.rf_10 [13] ), .B(_13603_ ), .S(_12982_ ), .Z(_13604_ ) );
MUX2_X1 _20617_ ( .A(\wbu.rf_11 [13] ), .B(_13604_ ), .S(_13036_ ), .Z(_13605_ ) );
MUX2_X1 _20618_ ( .A(\wbu.rf_12 [13] ), .B(_13605_ ), .S(_13043_ ), .Z(_13606_ ) );
MUX2_X1 _20619_ ( .A(\wbu.rf_13 [13] ), .B(_13606_ ), .S(_13052_ ), .Z(_13607_ ) );
AOI21_X1 _20620_ ( .A(_13595_ ), .B1(_13607_ ), .B2(_13058_ ), .ZN(_13608_ ) );
OAI211_X1 _20621_ ( .A(_13073_ ), .B(_13594_ ), .C1(_13608_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .ZN(_13609_ ) );
OAI211_X1 _20622_ ( .A(_13609_ ), .B(_13083_ ), .C1(\wbu.rf_16 [13] ), .C2(_13073_ ), .ZN(_13610_ ) );
NAND4_X1 _20623_ ( .A1(_12985_ ), .A2(fanout_net_31 ), .A3(\wbu.rf_17 [13] ), .A4(_08572_ ), .ZN(_13611_ ) );
AOI21_X1 _20624_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .B1(_13610_ ), .B2(_13611_ ), .ZN(_13612_ ) );
NAND3_X1 _20625_ ( .A1(_12989_ ), .A2(fanout_net_31 ), .A3(\wbu.rf_18 [13] ), .ZN(_13613_ ) );
NAND2_X1 _20626_ ( .A1(_13096_ ), .A2(_13613_ ), .ZN(_13614_ ) );
OAI221_X1 _20627_ ( .A(_13101_ ), .B1(\wbu.rf_19 [13] ), .B2(_13096_ ), .C1(_13612_ ), .C2(_13614_ ), .ZN(_13615_ ) );
NAND4_X1 _20628_ ( .A1(_13007_ ), .A2(fanout_net_32 ), .A3(\wbu.rf_20 [13] ), .A4(_13228_ ), .ZN(_13616_ ) );
NAND2_X1 _20629_ ( .A1(_13615_ ), .A2(_13616_ ), .ZN(_13617_ ) );
MUX2_X1 _20630_ ( .A(\wbu.rf_21 [13] ), .B(_13617_ ), .S(_13109_ ), .Z(_13618_ ) );
MUX2_X1 _20631_ ( .A(\wbu.rf_22 [13] ), .B(_13618_ ), .S(_13115_ ), .Z(_13619_ ) );
MUX2_X1 _20632_ ( .A(\wbu.rf_23 [13] ), .B(_13619_ ), .S(_13125_ ), .Z(_13620_ ) );
MUX2_X1 _20633_ ( .A(\wbu.rf_24 [13] ), .B(_13620_ ), .S(_13130_ ), .Z(_13621_ ) );
MUX2_X1 _20634_ ( .A(\wbu.rf_25 [13] ), .B(_13621_ ), .S(_13139_ ), .Z(_13622_ ) );
MUX2_X1 _20635_ ( .A(\wbu.rf_26 [13] ), .B(_13622_ ), .S(_13143_ ), .Z(_13623_ ) );
MUX2_X1 _20636_ ( .A(\wbu.rf_27 [13] ), .B(_13623_ ), .S(_13152_ ), .Z(_13624_ ) );
MUX2_X1 _20637_ ( .A(\wbu.rf_28 [13] ), .B(_13624_ ), .S(_13156_ ), .Z(_13625_ ) );
MUX2_X1 _20638_ ( .A(\wbu.rf_29 [13] ), .B(_13625_ ), .S(_13164_ ), .Z(_13626_ ) );
MUX2_X1 _20639_ ( .A(\wbu.rf_30 [13] ), .B(_13626_ ), .S(_13268_ ), .Z(_13627_ ) );
AOI211_X1 _20640_ ( .A(_13473_ ), .B(_13593_ ), .C1(_13627_ ), .C2(_13271_ ), .ZN(_13628_ ) );
INV_X1 _20641_ ( .A(\wbu.io_in_bits_rd_wdata [13] ), .ZN(_13629_ ) );
AOI211_X1 _20642_ ( .A(fanout_net_24 ), .B(_13628_ ), .C1(_13629_ ), .C2(_13373_ ), .ZN(_00356_ ) );
AND3_X1 _20643_ ( .A1(_13474_ ), .A2(fanout_net_32 ), .A3(\wbu.rf_31 [12] ), .ZN(_13630_ ) );
OAI21_X1 _20644_ ( .A(_13363_ ), .B1(_13145_ ), .B2(\wbu.rf_26 [12] ), .ZN(_13631_ ) );
NAND4_X1 _20645_ ( .A1(_13007_ ), .A2(fanout_net_38 ), .A3(_12966_ ), .A4(\wbu.rf_7 [12] ), .ZN(_13632_ ) );
NAND3_X1 _20646_ ( .A1(_13008_ ), .A2(fanout_net_38 ), .A3(\wbu.rf_5 [12] ), .ZN(_13633_ ) );
NAND2_X1 _20647_ ( .A1(_13018_ ), .A2(_13633_ ), .ZN(_13634_ ) );
MUX2_X1 _20648_ ( .A(\wbu._GEN_71 [12] ), .B(\wbu.rf_2 [12] ), .S(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .Z(_13635_ ) );
MUX2_X1 _20649_ ( .A(\wbu.rf_3 [12] ), .B(_13635_ ), .S(_12998_ ), .Z(_13636_ ) );
MUX2_X1 _20650_ ( .A(\wbu.rf_4 [12] ), .B(_13636_ ), .S(_13004_ ), .Z(_13637_ ) );
AOI21_X1 _20651_ ( .A(_13634_ ), .B1(_13637_ ), .B2(_13012_ ), .ZN(_13638_ ) );
OAI21_X1 _20652_ ( .A(_13024_ ), .B1(_13018_ ), .B2(\wbu.rf_6 [12] ), .ZN(_13639_ ) );
OAI211_X1 _20653_ ( .A(_13030_ ), .B(_13632_ ), .C1(_13638_ ), .C2(_13639_ ), .ZN(_13640_ ) );
OAI211_X1 _20654_ ( .A(_13640_ ), .B(_13383_ ), .C1(\wbu.rf_8 [12] ), .C2(_13030_ ), .ZN(_13641_ ) );
NAND4_X1 _20655_ ( .A1(_13061_ ), .A2(_13046_ ), .A3(fanout_net_38 ), .A4(\wbu.rf_9 [12] ), .ZN(_13642_ ) );
NAND3_X1 _20656_ ( .A1(_13641_ ), .A2(_13039_ ), .A3(_13642_ ), .ZN(_13643_ ) );
OAI211_X1 _20657_ ( .A(_13643_ ), .B(_13038_ ), .C1(\wbu.rf_10 [12] ), .C2(_13039_ ), .ZN(_13644_ ) );
NAND4_X1 _20658_ ( .A1(_13148_ ), .A2(fanout_net_38 ), .A3(_13047_ ), .A4(\wbu.rf_11 [12] ), .ZN(_13645_ ) );
NAND3_X1 _20659_ ( .A1(_13644_ ), .A2(_13055_ ), .A3(_13645_ ), .ZN(_13646_ ) );
OAI211_X1 _20660_ ( .A(_13646_ ), .B(_13054_ ), .C1(\wbu.rf_12 [12] ), .C2(_13055_ ), .ZN(_13647_ ) );
NAND4_X1 _20661_ ( .A1(_13062_ ), .A2(fanout_net_38 ), .A3(_13078_ ), .A4(\wbu.rf_13 [12] ), .ZN(_13648_ ) );
NAND3_X1 _20662_ ( .A1(_13647_ ), .A2(_13071_ ), .A3(_13648_ ), .ZN(_13649_ ) );
OAI211_X1 _20663_ ( .A(_13649_ ), .B(_13070_ ), .C1(\wbu.rf_14 [12] ), .C2(_13071_ ), .ZN(_13650_ ) );
NAND4_X1 _20664_ ( .A1(_13105_ ), .A2(_13079_ ), .A3(fanout_net_38 ), .A4(\wbu.rf_15 [12] ), .ZN(_13651_ ) );
NAND3_X1 _20665_ ( .A1(_13650_ ), .A2(_13087_ ), .A3(_13651_ ), .ZN(_13652_ ) );
OAI211_X1 _20666_ ( .A(_13652_ ), .B(_13086_ ), .C1(\wbu.rf_16 [12] ), .C2(_13087_ ), .ZN(_13653_ ) );
NAND4_X1 _20667_ ( .A1(_13119_ ), .A2(fanout_net_32 ), .A3(\wbu.rf_17 [12] ), .A4(_13497_ ), .ZN(_13654_ ) );
NAND3_X1 _20668_ ( .A1(_13653_ ), .A2(_13099_ ), .A3(_13654_ ), .ZN(_13655_ ) );
OAI211_X1 _20669_ ( .A(_13655_ ), .B(_13098_ ), .C1(\wbu.rf_18 [12] ), .C2(_13099_ ), .ZN(_13656_ ) );
NAND4_X1 _20670_ ( .A1(_13134_ ), .A2(_08575_ ), .A3(fanout_net_32 ), .A4(\wbu.rf_19 [12] ), .ZN(_13657_ ) );
NAND3_X1 _20671_ ( .A1(_13656_ ), .A2(_13113_ ), .A3(_13657_ ), .ZN(_13658_ ) );
OAI211_X1 _20672_ ( .A(_13658_ ), .B(_13112_ ), .C1(\wbu.rf_20 [12] ), .C2(_13113_ ), .ZN(_13659_ ) );
NAND4_X1 _20673_ ( .A1(_13146_ ), .A2(_13186_ ), .A3(fanout_net_32 ), .A4(\wbu.rf_21 [12] ), .ZN(_13660_ ) );
NAND3_X1 _20674_ ( .A1(_13659_ ), .A2(_13128_ ), .A3(_13660_ ), .ZN(_13661_ ) );
OAI211_X1 _20675_ ( .A(_13661_ ), .B(_13231_ ), .C1(\wbu.rf_22 [12] ), .C2(_13128_ ), .ZN(_13662_ ) );
NAND4_X1 _20676_ ( .A1(_13133_ ), .A2(fanout_net_32 ), .A3(_13160_ ), .A4(\wbu.rf_23 [12] ), .ZN(_13663_ ) );
AOI21_X1 _20677_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_1_Y ), .B1(_13662_ ), .B2(_13663_ ), .ZN(_13664_ ) );
AND4_X1 _20678_ ( .A1(fanout_net_32 ), .A2(_13378_ ), .A3(\wbu.rf_24 [12] ), .A4(_13229_ ), .ZN(_13665_ ) );
OAI21_X1 _20679_ ( .A(_13140_ ), .B1(_13664_ ), .B2(_13665_ ), .ZN(_13666_ ) );
AOI22_X1 _20680_ ( .A1(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .A2(\wbu.rf_25 [12] ), .B1(fanout_net_32 ), .B2(_12980_ ), .ZN(_13667_ ) );
AOI21_X1 _20681_ ( .A(_13631_ ), .B1(_13666_ ), .B2(_13667_ ), .ZN(_13668_ ) );
NAND3_X1 _20682_ ( .A1(_13034_ ), .A2(fanout_net_32 ), .A3(\wbu.rf_27 [12] ), .ZN(_13669_ ) );
NAND2_X1 _20683_ ( .A1(_13156_ ), .A2(_13669_ ), .ZN(_13670_ ) );
OAI221_X1 _20684_ ( .A(_13164_ ), .B1(\wbu.rf_28 [12] ), .B2(_13166_ ), .C1(_13668_ ), .C2(_13670_ ), .ZN(_13671_ ) );
NAND4_X1 _20685_ ( .A1(_13326_ ), .A2(fanout_net_32 ), .A3(_13327_ ), .A4(\wbu.rf_29 [12] ), .ZN(_13672_ ) );
NAND2_X1 _20686_ ( .A1(_13671_ ), .A2(_13672_ ), .ZN(_13673_ ) );
MUX2_X1 _20687_ ( .A(\wbu.rf_30 [12] ), .B(_13673_ ), .S(_13268_ ), .Z(_13674_ ) );
AOI211_X1 _20688_ ( .A(_13473_ ), .B(_13630_ ), .C1(_13674_ ), .C2(_13271_ ), .ZN(_13675_ ) );
INV_X1 _20689_ ( .A(\wbu.io_in_bits_rd_wdata [12] ), .ZN(_13676_ ) );
AOI211_X1 _20690_ ( .A(fanout_net_24 ), .B(_13675_ ), .C1(_13676_ ), .C2(_13373_ ), .ZN(_00357_ ) );
AND3_X1 _20691_ ( .A1(_13474_ ), .A2(fanout_net_32 ), .A3(\wbu.rf_31 [29] ), .ZN(_13677_ ) );
NAND4_X1 _20692_ ( .A1(_13061_ ), .A2(fanout_net_38 ), .A3(_13064_ ), .A4(\wbu.rf_13 [29] ), .ZN(_13678_ ) );
AND4_X1 _20693_ ( .A1(fanout_net_38 ), .A2(_13063_ ), .A3(\wbu.rf_12 [29] ), .A4(_12960_ ), .ZN(_13679_ ) );
MUX2_X1 _20694_ ( .A(\wbu._GEN_71 [29] ), .B(\wbu.rf_2 [29] ), .S(_12992_ ), .Z(_13680_ ) );
MUX2_X1 _20695_ ( .A(\wbu.rf_3 [29] ), .B(_13680_ ), .S(_12997_ ), .Z(_13681_ ) );
MUX2_X1 _20696_ ( .A(\wbu.rf_4 [29] ), .B(_13681_ ), .S(_13003_ ), .Z(_13682_ ) );
MUX2_X1 _20697_ ( .A(\wbu.rf_5 [29] ), .B(_13682_ ), .S(_13011_ ), .Z(_13683_ ) );
MUX2_X1 _20698_ ( .A(\wbu.rf_6 [29] ), .B(_13683_ ), .S(_13017_ ), .Z(_13684_ ) );
MUX2_X1 _20699_ ( .A(\wbu.rf_7 [29] ), .B(_13684_ ), .S(_13023_ ), .Z(_13685_ ) );
MUX2_X1 _20700_ ( .A(\wbu.rf_8 [29] ), .B(_13685_ ), .S(_13029_ ), .Z(_13686_ ) );
MUX2_X1 _20701_ ( .A(\wbu.rf_9 [29] ), .B(_13686_ ), .S(_13383_ ), .Z(_13687_ ) );
MUX2_X1 _20702_ ( .A(\wbu.rf_10 [29] ), .B(_13687_ ), .S(_12984_ ), .Z(_13688_ ) );
MUX2_X1 _20703_ ( .A(\wbu.rf_11 [29] ), .B(_13688_ ), .S(_13038_ ), .Z(_13689_ ) );
AOI21_X1 _20704_ ( .A(_13679_ ), .B1(_13689_ ), .B2(_13045_ ), .ZN(_13690_ ) );
OAI211_X1 _20705_ ( .A(_13059_ ), .B(_13678_ ), .C1(_13690_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_13691_ ) );
OAI211_X1 _20706_ ( .A(_13691_ ), .B(_13069_ ), .C1(\wbu.rf_14 [29] ), .C2(_13060_ ), .ZN(_13692_ ) );
NAND4_X1 _20707_ ( .A1(_13047_ ), .A2(_13078_ ), .A3(fanout_net_38 ), .A4(\wbu.rf_15 [29] ), .ZN(_13693_ ) );
NAND3_X1 _20708_ ( .A1(_13692_ ), .A2(_13075_ ), .A3(_13693_ ), .ZN(_13694_ ) );
OAI211_X1 _20709_ ( .A(_13694_ ), .B(_13085_ ), .C1(\wbu.rf_16 [29] ), .C2(_13076_ ), .ZN(_13695_ ) );
NAND4_X1 _20710_ ( .A1(_13092_ ), .A2(fanout_net_32 ), .A3(\wbu.rf_17 [29] ), .A4(_13350_ ), .ZN(_13696_ ) );
NAND3_X1 _20711_ ( .A1(_13695_ ), .A2(_13091_ ), .A3(_13696_ ), .ZN(_13697_ ) );
OAI211_X1 _20712_ ( .A(_13697_ ), .B(_13097_ ), .C1(\wbu.rf_18 [29] ), .C2(_13450_ ), .ZN(_13698_ ) );
NAND4_X1 _20713_ ( .A1(_13105_ ), .A2(_13497_ ), .A3(fanout_net_32 ), .A4(\wbu.rf_19 [29] ), .ZN(_13699_ ) );
NAND3_X1 _20714_ ( .A1(_13698_ ), .A2(_13103_ ), .A3(_13699_ ), .ZN(_13700_ ) );
OAI211_X1 _20715_ ( .A(_13700_ ), .B(_13111_ ), .C1(\wbu.rf_20 [29] ), .C2(_13104_ ), .ZN(_13701_ ) );
NAND4_X1 _20716_ ( .A1(_13119_ ), .A2(_13121_ ), .A3(fanout_net_32 ), .A4(\wbu.rf_21 [29] ), .ZN(_13702_ ) );
NAND3_X1 _20717_ ( .A1(_13701_ ), .A2(_13117_ ), .A3(_13702_ ), .ZN(_13703_ ) );
OAI211_X1 _20718_ ( .A(_13703_ ), .B(_13126_ ), .C1(\wbu.rf_22 [29] ), .C2(_13118_ ), .ZN(_13704_ ) );
NAND4_X1 _20719_ ( .A1(_13186_ ), .A2(fanout_net_32 ), .A3(_13134_ ), .A4(\wbu.rf_23 [29] ), .ZN(_13705_ ) );
NAND3_X1 _20720_ ( .A1(_13704_ ), .A2(_13131_ ), .A3(_13705_ ), .ZN(_13706_ ) );
OAI211_X1 _20721_ ( .A(_13706_ ), .B(_13460_ ), .C1(\wbu.rf_24 [29] ), .C2(_13414_ ), .ZN(_13707_ ) );
NAND4_X1 _20722_ ( .A1(_13146_ ), .A2(_13378_ ), .A3(fanout_net_32 ), .A4(\wbu.rf_25 [29] ), .ZN(_13708_ ) );
NAND3_X1 _20723_ ( .A1(_13707_ ), .A2(_13144_ ), .A3(_13708_ ), .ZN(_13709_ ) );
OAI211_X1 _20724_ ( .A(_13709_ ), .B(_13363_ ), .C1(\wbu.rf_26 [29] ), .C2(_13260_ ), .ZN(_13710_ ) );
NAND4_X1 _20725_ ( .A1(_13158_ ), .A2(fanout_net_32 ), .A3(_13160_ ), .A4(\wbu.rf_27 [29] ), .ZN(_13711_ ) );
NAND3_X1 _20726_ ( .A1(_13710_ ), .A2(_13166_ ), .A3(_13711_ ), .ZN(_13712_ ) );
OAI211_X1 _20727_ ( .A(_13712_ ), .B(_13512_ ), .C1(\wbu.rf_28 [29] ), .C2(_13365_ ), .ZN(_13713_ ) );
NAND4_X1 _20728_ ( .A1(_13326_ ), .A2(fanout_net_32 ), .A3(_13327_ ), .A4(\wbu.rf_29 [29] ), .ZN(_13714_ ) );
NAND2_X1 _20729_ ( .A1(_13713_ ), .A2(_13714_ ), .ZN(_13715_ ) );
MUX2_X1 _20730_ ( .A(\wbu.rf_30 [29] ), .B(_13715_ ), .S(_13267_ ), .Z(_13716_ ) );
AOI211_X1 _20731_ ( .A(_13473_ ), .B(_13677_ ), .C1(_13716_ ), .C2(_13271_ ), .ZN(_13717_ ) );
INV_X1 _20732_ ( .A(\wbu.io_in_bits_rd_wdata [29] ), .ZN(_13718_ ) );
AOI211_X1 _20733_ ( .A(fanout_net_24 ), .B(_13717_ ), .C1(_13718_ ), .C2(_13373_ ), .ZN(_00358_ ) );
INV_X1 _20734_ ( .A(\wbu.io_in_bits_rd_wdata [11] ), .ZN(_13719_ ) );
NAND4_X1 _20735_ ( .A1(_13186_ ), .A2(fanout_net_32 ), .A3(_13134_ ), .A4(\wbu.rf_23 [11] ), .ZN(_13720_ ) );
AND4_X1 _20736_ ( .A1(fanout_net_32 ), .A2(_13174_ ), .A3(_13188_ ), .A4(\wbu.rf_22 [11] ), .ZN(_13721_ ) );
MUX2_X1 _20737_ ( .A(\wbu._GEN_71 [11] ), .B(\wbu.rf_2 [11] ), .S(_12991_ ), .Z(_13722_ ) );
MUX2_X1 _20738_ ( .A(\wbu.rf_3 [11] ), .B(_13722_ ), .S(_12996_ ), .Z(_13723_ ) );
MUX2_X1 _20739_ ( .A(\wbu.rf_4 [11] ), .B(_13723_ ), .S(_13002_ ), .Z(_13724_ ) );
MUX2_X1 _20740_ ( .A(\wbu.rf_5 [11] ), .B(_13724_ ), .S(_13010_ ), .Z(_13725_ ) );
MUX2_X1 _20741_ ( .A(\wbu.rf_6 [11] ), .B(_13725_ ), .S(_13016_ ), .Z(_13726_ ) );
MUX2_X1 _20742_ ( .A(\wbu.rf_7 [11] ), .B(_13726_ ), .S(_13022_ ), .Z(_13727_ ) );
MUX2_X1 _20743_ ( .A(\wbu.rf_8 [11] ), .B(_13727_ ), .S(_13028_ ), .Z(_13728_ ) );
MUX2_X1 _20744_ ( .A(\wbu.rf_9 [11] ), .B(_13728_ ), .S(_13197_ ), .Z(_13729_ ) );
MUX2_X1 _20745_ ( .A(\wbu.rf_10 [11] ), .B(_13729_ ), .S(_12982_ ), .Z(_13730_ ) );
MUX2_X1 _20746_ ( .A(\wbu.rf_11 [11] ), .B(_13730_ ), .S(_13036_ ), .Z(_13731_ ) );
MUX2_X1 _20747_ ( .A(\wbu.rf_12 [11] ), .B(_13731_ ), .S(_13043_ ), .Z(_13732_ ) );
MUX2_X1 _20748_ ( .A(\wbu.rf_13 [11] ), .B(_13732_ ), .S(_13052_ ), .Z(_13733_ ) );
MUX2_X1 _20749_ ( .A(\wbu.rf_14 [11] ), .B(_13733_ ), .S(_13058_ ), .Z(_13734_ ) );
MUX2_X1 _20750_ ( .A(\wbu.rf_15 [11] ), .B(_13734_ ), .S(_13068_ ), .Z(_13735_ ) );
MUX2_X1 _20751_ ( .A(\wbu.rf_16 [11] ), .B(_13735_ ), .S(_13074_ ), .Z(_13736_ ) );
MUX2_X1 _20752_ ( .A(\wbu.rf_17 [11] ), .B(_13736_ ), .S(_13084_ ), .Z(_13737_ ) );
MUX2_X1 _20753_ ( .A(\wbu.rf_18 [11] ), .B(_13737_ ), .S(_13090_ ), .Z(_13738_ ) );
MUX2_X1 _20754_ ( .A(\wbu.rf_19 [11] ), .B(_13738_ ), .S(_13097_ ), .Z(_13739_ ) );
MUX2_X1 _20755_ ( .A(\wbu.rf_20 [11] ), .B(_13739_ ), .S(_13103_ ), .Z(_13740_ ) );
MUX2_X1 _20756_ ( .A(\wbu.rf_21 [11] ), .B(_13740_ ), .S(_13111_ ), .Z(_13741_ ) );
AOI21_X1 _20757_ ( .A(_13721_ ), .B1(_13741_ ), .B2(_13212_ ), .ZN(_13742_ ) );
OAI211_X1 _20758_ ( .A(_13132_ ), .B(_13720_ ), .C1(_13742_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .ZN(_13743_ ) );
OAI211_X1 _20759_ ( .A(_13743_ ), .B(_13460_ ), .C1(\wbu.rf_24 [11] ), .C2(_13141_ ), .ZN(_13744_ ) );
NAND4_X1 _20760_ ( .A1(_13312_ ), .A2(_13149_ ), .A3(fanout_net_32 ), .A4(\wbu.rf_25 [11] ), .ZN(_13745_ ) );
NAND3_X1 _20761_ ( .A1(_13744_ ), .A2(_13145_ ), .A3(_13745_ ), .ZN(_13746_ ) );
OAI211_X1 _20762_ ( .A(_13746_ ), .B(_13218_ ), .C1(\wbu.rf_26 [11] ), .C2(_13154_ ), .ZN(_13747_ ) );
NAND4_X1 _20763_ ( .A1(_13159_ ), .A2(fanout_net_32 ), .A3(_13161_ ), .A4(\wbu.rf_27 [11] ), .ZN(_13748_ ) );
NAND3_X1 _20764_ ( .A1(_13747_ ), .A2(_13157_ ), .A3(_13748_ ), .ZN(_13749_ ) );
OAI211_X1 _20765_ ( .A(_13749_ ), .B(_13512_ ), .C1(\wbu.rf_28 [11] ), .C2(_13167_ ), .ZN(_13750_ ) );
NAND4_X1 _20766_ ( .A1(_13169_ ), .A2(fanout_net_32 ), .A3(_13176_ ), .A4(\wbu.rf_29 [11] ), .ZN(_13751_ ) );
AOI21_X1 _20767_ ( .A(_12975_ ), .B1(_13750_ ), .B2(_13751_ ), .ZN(_13752_ ) );
AND4_X1 _20768_ ( .A1(fanout_net_32 ), .A2(_13175_ ), .A3(\wbu.rf_30 [11] ), .A4(_13376_ ), .ZN(_13753_ ) );
OAI21_X1 _20769_ ( .A(_13369_ ), .B1(_13752_ ), .B2(_13753_ ), .ZN(_13754_ ) );
AOI22_X1 _20770_ ( .A1(_13179_ ), .A2(\wbu.rf_31 [11] ), .B1(_13180_ ), .B2(_13182_ ), .ZN(_13755_ ) );
AOI221_X4 _20771_ ( .A(fanout_net_24 ), .B1(_13719_ ), .B2(_12965_ ), .C1(_13754_ ), .C2(_13755_ ), .ZN(_00359_ ) );
INV_X1 _20772_ ( .A(\wbu.io_in_bits_rd_wdata [10] ), .ZN(_13756_ ) );
OR2_X1 _20773_ ( .A1(_13054_ ), .A2(\wbu.rf_13 [10] ), .ZN(_13757_ ) );
MUX2_X1 _20774_ ( .A(\wbu._GEN_71 [10] ), .B(\wbu.rf_2 [10] ), .S(_12992_ ), .Z(_13758_ ) );
MUX2_X1 _20775_ ( .A(\wbu.rf_3 [10] ), .B(_13758_ ), .S(_12997_ ), .Z(_13759_ ) );
MUX2_X1 _20776_ ( .A(\wbu.rf_4 [10] ), .B(_13759_ ), .S(_13003_ ), .Z(_13760_ ) );
MUX2_X1 _20777_ ( .A(\wbu.rf_5 [10] ), .B(_13760_ ), .S(_13011_ ), .Z(_13761_ ) );
MUX2_X1 _20778_ ( .A(\wbu.rf_6 [10] ), .B(_13761_ ), .S(_13017_ ), .Z(_13762_ ) );
MUX2_X1 _20779_ ( .A(\wbu.rf_7 [10] ), .B(_13762_ ), .S(_13023_ ), .Z(_13763_ ) );
MUX2_X1 _20780_ ( .A(\wbu.rf_8 [10] ), .B(_13763_ ), .S(_13029_ ), .Z(_13764_ ) );
MUX2_X1 _20781_ ( .A(\wbu.rf_9 [10] ), .B(_13764_ ), .S(_13383_ ), .Z(_13765_ ) );
MUX2_X1 _20782_ ( .A(\wbu.rf_10 [10] ), .B(_13765_ ), .S(_12984_ ), .Z(_13766_ ) );
MUX2_X1 _20783_ ( .A(\wbu.rf_11 [10] ), .B(_13766_ ), .S(_13038_ ), .Z(_13767_ ) );
MUX2_X1 _20784_ ( .A(\wbu.rf_12 [10] ), .B(_13767_ ), .S(_13055_ ), .Z(_13768_ ) );
OAI211_X1 _20785_ ( .A(_13060_ ), .B(_13757_ ), .C1(_13768_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_13769_ ) );
NAND4_X1 _20786_ ( .A1(_13173_ ), .A2(fanout_net_38 ), .A3(_13078_ ), .A4(\wbu.rf_14 [10] ), .ZN(_13770_ ) );
AOI21_X1 _20787_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .B1(_13769_ ), .B2(_13770_ ), .ZN(_13771_ ) );
NAND3_X1 _20788_ ( .A1(_12968_ ), .A2(fanout_net_38 ), .A3(\wbu.rf_15 [10] ), .ZN(_13772_ ) );
INV_X1 _20789_ ( .A(_12961_ ), .ZN(_13773_ ) );
OAI21_X1 _20790_ ( .A(_13772_ ), .B1(_08571_ ), .B2(_13773_ ), .ZN(_13774_ ) );
OAI221_X1 _20791_ ( .A(_13085_ ), .B1(\wbu.rf_16 [10] ), .B2(_13076_ ), .C1(_13771_ ), .C2(_13774_ ), .ZN(_13775_ ) );
NAND4_X1 _20792_ ( .A1(_13092_ ), .A2(fanout_net_32 ), .A3(\wbu.rf_17 [10] ), .A4(_08574_ ), .ZN(_13776_ ) );
NAND3_X1 _20793_ ( .A1(_13775_ ), .A2(_13091_ ), .A3(_13776_ ), .ZN(_13777_ ) );
OAI211_X1 _20794_ ( .A(_13777_ ), .B(_13097_ ), .C1(\wbu.rf_18 [10] ), .C2(_13450_ ), .ZN(_13778_ ) );
NAND4_X1 _20795_ ( .A1(_13106_ ), .A2(_13497_ ), .A3(fanout_net_32 ), .A4(\wbu.rf_19 [10] ), .ZN(_13779_ ) );
NAND3_X1 _20796_ ( .A1(_13778_ ), .A2(_13104_ ), .A3(_13779_ ), .ZN(_13780_ ) );
OAI211_X1 _20797_ ( .A(_13780_ ), .B(_13111_ ), .C1(\wbu.rf_20 [10] ), .C2(_13381_ ), .ZN(_13781_ ) );
NAND4_X1 _20798_ ( .A1(_13120_ ), .A2(_13188_ ), .A3(fanout_net_32 ), .A4(\wbu.rf_21 [10] ), .ZN(_13782_ ) );
NAND3_X1 _20799_ ( .A1(_13781_ ), .A2(_13118_ ), .A3(_13782_ ), .ZN(_13783_ ) );
OAI211_X1 _20800_ ( .A(_13783_ ), .B(_13127_ ), .C1(\wbu.rf_22 [10] ), .C2(_13212_ ), .ZN(_13784_ ) );
NAND4_X1 _20801_ ( .A1(_13133_ ), .A2(fanout_net_32 ), .A3(_13135_ ), .A4(\wbu.rf_23 [10] ), .ZN(_13785_ ) );
NAND3_X1 _20802_ ( .A1(_13784_ ), .A2(_13132_ ), .A3(_13785_ ), .ZN(_13786_ ) );
OAI211_X1 _20803_ ( .A(_13786_ ), .B(_13460_ ), .C1(\wbu.rf_24 [10] ), .C2(_13141_ ), .ZN(_13787_ ) );
NAND4_X1 _20804_ ( .A1(_13312_ ), .A2(_13149_ ), .A3(fanout_net_32 ), .A4(\wbu.rf_25 [10] ), .ZN(_13788_ ) );
NAND3_X1 _20805_ ( .A1(_13787_ ), .A2(_13145_ ), .A3(_13788_ ), .ZN(_13789_ ) );
OAI211_X1 _20806_ ( .A(_13789_ ), .B(_13218_ ), .C1(\wbu.rf_26 [10] ), .C2(_13260_ ), .ZN(_13790_ ) );
NAND4_X1 _20807_ ( .A1(_13159_ ), .A2(fanout_net_32 ), .A3(_13161_ ), .A4(\wbu.rf_27 [10] ), .ZN(_13791_ ) );
NAND3_X1 _20808_ ( .A1(_13790_ ), .A2(_13157_ ), .A3(_13791_ ), .ZN(_13792_ ) );
OAI211_X1 _20809_ ( .A(_13792_ ), .B(_13512_ ), .C1(\wbu.rf_28 [10] ), .C2(_13167_ ), .ZN(_13793_ ) );
NAND4_X1 _20810_ ( .A1(_13169_ ), .A2(fanout_net_33 ), .A3(_13176_ ), .A4(\wbu.rf_29 [10] ), .ZN(_13794_ ) );
AOI21_X1 _20811_ ( .A(_12975_ ), .B1(_13793_ ), .B2(_13794_ ), .ZN(_13795_ ) );
AND4_X1 _20812_ ( .A1(fanout_net_33 ), .A2(_13175_ ), .A3(\wbu.rf_30 [10] ), .A4(_13376_ ), .ZN(_13796_ ) );
OAI21_X1 _20813_ ( .A(_13369_ ), .B1(_13795_ ), .B2(_13796_ ), .ZN(_13797_ ) );
AOI22_X1 _20814_ ( .A1(_13179_ ), .A2(\wbu.rf_31 [10] ), .B1(_13180_ ), .B2(_13182_ ), .ZN(_13798_ ) );
AOI221_X4 _20815_ ( .A(fanout_net_24 ), .B1(_13756_ ), .B2(_12965_ ), .C1(_13797_ ), .C2(_13798_ ), .ZN(_00360_ ) );
INV_X1 _20816_ ( .A(\wbu.io_in_bits_rd_wdata [9] ), .ZN(_13799_ ) );
NAND4_X1 _20817_ ( .A1(_13077_ ), .A2(_13078_ ), .A3(fanout_net_38 ), .A4(\wbu.rf_15 [9] ), .ZN(_13800_ ) );
AND4_X1 _20818_ ( .A1(fanout_net_38 ), .A2(_13173_ ), .A3(\wbu.rf_14 [9] ), .A4(_13064_ ), .ZN(_13801_ ) );
NAND3_X1 _20819_ ( .A1(_13026_ ), .A2(fanout_net_38 ), .A3(\wbu.rf_8 [9] ), .ZN(_13802_ ) );
AND4_X1 _20820_ ( .A1(fanout_net_38 ), .A2(_12977_ ), .A3(_13007_ ), .A4(\wbu.rf_6 [9] ), .ZN(_13803_ ) );
MUX2_X1 _20821_ ( .A(\wbu._GEN_71 [9] ), .B(\wbu.rf_2 [9] ), .S(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .Z(_13804_ ) );
MUX2_X1 _20822_ ( .A(\wbu.rf_3 [9] ), .B(_13804_ ), .S(_12998_ ), .Z(_13805_ ) );
MUX2_X1 _20823_ ( .A(\wbu.rf_4 [9] ), .B(_13805_ ), .S(_13004_ ), .Z(_13806_ ) );
MUX2_X1 _20824_ ( .A(\wbu.rf_5 [9] ), .B(_13806_ ), .S(_13012_ ), .Z(_13807_ ) );
AOI211_X1 _20825_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_Y ), .B(_13803_ ), .C1(_13807_ ), .C2(_13018_ ), .ZN(_13808_ ) );
OAI21_X1 _20826_ ( .A(_13029_ ), .B1(_13024_ ), .B2(\wbu.rf_7 [9] ), .ZN(_13809_ ) );
OAI21_X1 _20827_ ( .A(_13802_ ), .B1(_13808_ ), .B2(_13809_ ), .ZN(_13810_ ) );
MUX2_X1 _20828_ ( .A(\wbu.rf_9 [9] ), .B(_13810_ ), .S(_13383_ ), .Z(_13811_ ) );
MUX2_X1 _20829_ ( .A(\wbu.rf_10 [9] ), .B(_13811_ ), .S(_12984_ ), .Z(_13812_ ) );
MUX2_X1 _20830_ ( .A(\wbu.rf_11 [9] ), .B(_13812_ ), .S(_13037_ ), .Z(_13813_ ) );
MUX2_X1 _20831_ ( .A(\wbu.rf_12 [9] ), .B(_13813_ ), .S(_13044_ ), .Z(_13814_ ) );
MUX2_X1 _20832_ ( .A(\wbu.rf_13 [9] ), .B(_13814_ ), .S(_13053_ ), .Z(_13815_ ) );
AOI21_X1 _20833_ ( .A(_13801_ ), .B1(_13815_ ), .B2(_13060_ ), .ZN(_13816_ ) );
OAI211_X1 _20834_ ( .A(_13075_ ), .B(_13800_ ), .C1(_13816_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .ZN(_13817_ ) );
OAI211_X1 _20835_ ( .A(_13817_ ), .B(_13086_ ), .C1(\wbu.rf_16 [9] ), .C2(_13087_ ), .ZN(_13818_ ) );
NAND4_X1 _20836_ ( .A1(_13092_ ), .A2(fanout_net_33 ), .A3(\wbu.rf_17 [9] ), .A4(_08574_ ), .ZN(_13819_ ) );
NAND3_X1 _20837_ ( .A1(_13818_ ), .A2(_13091_ ), .A3(_13819_ ), .ZN(_13820_ ) );
OAI211_X1 _20838_ ( .A(_13820_ ), .B(_13097_ ), .C1(\wbu.rf_18 [9] ), .C2(_13450_ ), .ZN(_13821_ ) );
NAND4_X1 _20839_ ( .A1(_13106_ ), .A2(_13497_ ), .A3(fanout_net_33 ), .A4(\wbu.rf_19 [9] ), .ZN(_13822_ ) );
NAND3_X1 _20840_ ( .A1(_13821_ ), .A2(_13104_ ), .A3(_13822_ ), .ZN(_13823_ ) );
OAI211_X1 _20841_ ( .A(_13823_ ), .B(_13111_ ), .C1(\wbu.rf_20 [9] ), .C2(_13381_ ), .ZN(_13824_ ) );
NAND4_X1 _20842_ ( .A1(_13120_ ), .A2(_13188_ ), .A3(fanout_net_33 ), .A4(\wbu.rf_21 [9] ), .ZN(_13825_ ) );
NAND3_X1 _20843_ ( .A1(_13824_ ), .A2(_13118_ ), .A3(_13825_ ), .ZN(_13826_ ) );
OAI211_X1 _20844_ ( .A(_13826_ ), .B(_13127_ ), .C1(\wbu.rf_22 [9] ), .C2(_13212_ ), .ZN(_13827_ ) );
NAND4_X1 _20845_ ( .A1(_13133_ ), .A2(fanout_net_33 ), .A3(_13135_ ), .A4(\wbu.rf_23 [9] ), .ZN(_13828_ ) );
NAND3_X1 _20846_ ( .A1(_13827_ ), .A2(_13132_ ), .A3(_13828_ ), .ZN(_13829_ ) );
OAI211_X1 _20847_ ( .A(_13829_ ), .B(_13460_ ), .C1(\wbu.rf_24 [9] ), .C2(_13141_ ), .ZN(_13830_ ) );
NAND4_X1 _20848_ ( .A1(_13312_ ), .A2(_13149_ ), .A3(fanout_net_33 ), .A4(\wbu.rf_25 [9] ), .ZN(_13831_ ) );
NAND3_X1 _20849_ ( .A1(_13830_ ), .A2(_13144_ ), .A3(_13831_ ), .ZN(_13832_ ) );
OAI211_X1 _20850_ ( .A(_13832_ ), .B(_13218_ ), .C1(\wbu.rf_26 [9] ), .C2(_13260_ ), .ZN(_13833_ ) );
NAND4_X1 _20851_ ( .A1(_13159_ ), .A2(fanout_net_33 ), .A3(_13160_ ), .A4(\wbu.rf_27 [9] ), .ZN(_13834_ ) );
NAND3_X1 _20852_ ( .A1(_13833_ ), .A2(_13166_ ), .A3(_13834_ ), .ZN(_13835_ ) );
OAI211_X1 _20853_ ( .A(_13835_ ), .B(_13512_ ), .C1(\wbu.rf_28 [9] ), .C2(_13167_ ), .ZN(_13836_ ) );
NAND4_X1 _20854_ ( .A1(_13169_ ), .A2(fanout_net_33 ), .A3(_13176_ ), .A4(\wbu.rf_29 [9] ), .ZN(_13837_ ) );
AOI21_X1 _20855_ ( .A(_12975_ ), .B1(_13836_ ), .B2(_13837_ ), .ZN(_13838_ ) );
AND4_X1 _20856_ ( .A1(fanout_net_33 ), .A2(_13175_ ), .A3(\wbu.rf_30 [9] ), .A4(_13376_ ), .ZN(_13839_ ) );
OAI21_X1 _20857_ ( .A(_13369_ ), .B1(_13838_ ), .B2(_13839_ ), .ZN(_13840_ ) );
AOI22_X1 _20858_ ( .A1(_12969_ ), .A2(\wbu.rf_31 [9] ), .B1(_13180_ ), .B2(_13182_ ), .ZN(_13841_ ) );
AOI221_X4 _20859_ ( .A(fanout_net_24 ), .B1(_13799_ ), .B2(_12965_ ), .C1(_13840_ ), .C2(_13841_ ), .ZN(_00361_ ) );
OR2_X1 _20860_ ( .A1(_13374_ ), .A2(\wbu.rf_31 [8] ), .ZN(_13842_ ) );
NAND4_X1 _20861_ ( .A1(_13046_ ), .A2(fanout_net_38 ), .A3(_13047_ ), .A4(\wbu.rf_11 [8] ), .ZN(_13843_ ) );
AND4_X1 _20862_ ( .A1(fanout_net_38 ), .A2(_12977_ ), .A3(_13046_ ), .A4(\wbu.rf_10 [8] ), .ZN(_13844_ ) );
MUX2_X1 _20863_ ( .A(\wbu._GEN_71 [8] ), .B(\wbu.rf_2 [8] ), .S(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .Z(_13845_ ) );
MUX2_X1 _20864_ ( .A(\wbu.rf_3 [8] ), .B(_13845_ ), .S(_12998_ ), .Z(_13846_ ) );
MUX2_X1 _20865_ ( .A(\wbu.rf_4 [8] ), .B(_13846_ ), .S(_13004_ ), .Z(_13847_ ) );
MUX2_X1 _20866_ ( .A(\wbu.rf_5 [8] ), .B(_13847_ ), .S(_13012_ ), .Z(_13848_ ) );
MUX2_X1 _20867_ ( .A(\wbu.rf_6 [8] ), .B(_13848_ ), .S(_13018_ ), .Z(_13849_ ) );
MUX2_X1 _20868_ ( .A(\wbu.rf_7 [8] ), .B(_13849_ ), .S(_13024_ ), .Z(_13850_ ) );
MUX2_X1 _20869_ ( .A(\wbu.rf_8 [8] ), .B(_13850_ ), .S(_13030_ ), .Z(_13851_ ) );
MUX2_X1 _20870_ ( .A(\wbu.rf_9 [8] ), .B(_13851_ ), .S(_13383_ ), .Z(_13852_ ) );
AOI21_X1 _20871_ ( .A(_13844_ ), .B1(_13852_ ), .B2(_13039_ ), .ZN(_13853_ ) );
OAI211_X1 _20872_ ( .A(_13045_ ), .B(_13843_ ), .C1(_13853_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .ZN(_13854_ ) );
OAI211_X1 _20873_ ( .A(_13854_ ), .B(_13054_ ), .C1(\wbu.rf_12 [8] ), .C2(_13055_ ), .ZN(_13855_ ) );
NAND4_X1 _20874_ ( .A1(_13062_ ), .A2(fanout_net_38 ), .A3(_13064_ ), .A4(\wbu.rf_13 [8] ), .ZN(_13856_ ) );
NAND3_X1 _20875_ ( .A1(_13855_ ), .A2(_13060_ ), .A3(_13856_ ), .ZN(_13857_ ) );
OAI211_X1 _20876_ ( .A(_13857_ ), .B(_13070_ ), .C1(\wbu.rf_14 [8] ), .C2(_13071_ ), .ZN(_13858_ ) );
NAND4_X1 _20877_ ( .A1(_13077_ ), .A2(_13079_ ), .A3(fanout_net_38 ), .A4(\wbu.rf_15 [8] ), .ZN(_13859_ ) );
NAND3_X1 _20878_ ( .A1(_13858_ ), .A2(_13076_ ), .A3(_13859_ ), .ZN(_13860_ ) );
OAI211_X1 _20879_ ( .A(_13860_ ), .B(_13086_ ), .C1(\wbu.rf_16 [8] ), .C2(_13087_ ), .ZN(_13861_ ) );
NAND4_X1 _20880_ ( .A1(_13119_ ), .A2(fanout_net_33 ), .A3(\wbu.rf_17 [8] ), .A4(_08574_ ), .ZN(_13862_ ) );
NAND3_X1 _20881_ ( .A1(_13861_ ), .A2(_13450_ ), .A3(_13862_ ), .ZN(_13863_ ) );
OAI211_X1 _20882_ ( .A(_13863_ ), .B(_13098_ ), .C1(\wbu.rf_18 [8] ), .C2(_13099_ ), .ZN(_13864_ ) );
NAND4_X1 _20883_ ( .A1(_13106_ ), .A2(_08575_ ), .A3(fanout_net_33 ), .A4(\wbu.rf_19 [8] ), .ZN(_13865_ ) );
NAND3_X1 _20884_ ( .A1(_13864_ ), .A2(_13381_ ), .A3(_13865_ ), .ZN(_13866_ ) );
OAI211_X1 _20885_ ( .A(_13866_ ), .B(_13112_ ), .C1(\wbu.rf_20 [8] ), .C2(_13113_ ), .ZN(_13867_ ) );
NAND4_X1 _20886_ ( .A1(_13120_ ), .A2(_13122_ ), .A3(fanout_net_33 ), .A4(\wbu.rf_21 [8] ), .ZN(_13868_ ) );
NAND3_X1 _20887_ ( .A1(_13867_ ), .A2(_13118_ ), .A3(_13868_ ), .ZN(_13869_ ) );
OAI211_X1 _20888_ ( .A(_13869_ ), .B(_13231_ ), .C1(\wbu.rf_22 [8] ), .C2(_13128_ ), .ZN(_13870_ ) );
NAND4_X1 _20889_ ( .A1(_13133_ ), .A2(fanout_net_33 ), .A3(_13135_ ), .A4(\wbu.rf_23 [8] ), .ZN(_13871_ ) );
NAND3_X1 _20890_ ( .A1(_13870_ ), .A2(_13414_ ), .A3(_13871_ ), .ZN(_13872_ ) );
OAI211_X1 _20891_ ( .A(_13872_ ), .B(_13140_ ), .C1(\wbu.rf_24 [8] ), .C2(_13141_ ), .ZN(_13873_ ) );
NAND4_X1 _20892_ ( .A1(_13147_ ), .A2(_13158_ ), .A3(fanout_net_33 ), .A4(\wbu.rf_25 [8] ), .ZN(_13874_ ) );
NAND3_X1 _20893_ ( .A1(_13873_ ), .A2(_13260_ ), .A3(_13874_ ), .ZN(_13875_ ) );
OAI211_X1 _20894_ ( .A(_13875_ ), .B(_13153_ ), .C1(\wbu.rf_26 [8] ), .C2(_13154_ ), .ZN(_13876_ ) );
NAND4_X1 _20895_ ( .A1(_13159_ ), .A2(fanout_net_33 ), .A3(_13161_ ), .A4(\wbu.rf_27 [8] ), .ZN(_13877_ ) );
NAND3_X1 _20896_ ( .A1(_13876_ ), .A2(_13365_ ), .A3(_13877_ ), .ZN(_13878_ ) );
OAI211_X1 _20897_ ( .A(_13878_ ), .B(_13165_ ), .C1(\wbu.rf_28 [8] ), .C2(_13167_ ), .ZN(_13879_ ) );
NAND4_X1 _20898_ ( .A1(_13169_ ), .A2(fanout_net_33 ), .A3(_13170_ ), .A4(\wbu.rf_29 [8] ), .ZN(_13880_ ) );
NAND2_X1 _20899_ ( .A1(_13879_ ), .A2(_13880_ ), .ZN(_13881_ ) );
MUX2_X1 _20900_ ( .A(\wbu.rf_30 [8] ), .B(_13881_ ), .S(_13268_ ), .Z(_13882_ ) );
OAI211_X1 _20901_ ( .A(_13276_ ), .B(_13842_ ), .C1(_13882_ ), .C2(_13179_ ), .ZN(_13883_ ) );
NAND3_X1 _20902_ ( .A1(_13181_ ), .A2(\wbu.io_in_bits_rd_wdata [8] ), .A3(_13183_ ), .ZN(_13884_ ) );
AOI21_X1 _20903_ ( .A(fanout_net_24 ), .B1(_13883_ ), .B2(_13884_ ), .ZN(_00362_ ) );
NAND4_X1 _20904_ ( .A1(_13376_ ), .A2(_13229_ ), .A3(fanout_net_33 ), .A4(\wbu.rf_28 [7] ), .ZN(_13885_ ) );
AND4_X1 _20905_ ( .A1(fanout_net_33 ), .A2(_13158_ ), .A3(\wbu.rf_27 [7] ), .A4(_13160_ ), .ZN(_13886_ ) );
MUX2_X1 _20906_ ( .A(\wbu._GEN_71 [7] ), .B(\wbu.rf_2 [7] ), .S(_12990_ ), .Z(_13887_ ) );
MUX2_X1 _20907_ ( .A(\wbu.rf_3 [7] ), .B(_13887_ ), .S(_12995_ ), .Z(_13888_ ) );
MUX2_X1 _20908_ ( .A(\wbu.rf_4 [7] ), .B(_13888_ ), .S(_13001_ ), .Z(_13889_ ) );
MUX2_X1 _20909_ ( .A(\wbu.rf_5 [7] ), .B(_13889_ ), .S(_13009_ ), .Z(_13890_ ) );
MUX2_X1 _20910_ ( .A(\wbu.rf_6 [7] ), .B(_13890_ ), .S(_13015_ ), .Z(_13891_ ) );
MUX2_X1 _20911_ ( .A(\wbu.rf_7 [7] ), .B(_13891_ ), .S(_13021_ ), .Z(_13892_ ) );
MUX2_X1 _20912_ ( .A(\wbu.rf_8 [7] ), .B(_13892_ ), .S(_13027_ ), .Z(_13893_ ) );
MUX2_X1 _20913_ ( .A(\wbu.rf_9 [7] ), .B(_13893_ ), .S(_13197_ ), .Z(_13894_ ) );
MUX2_X1 _20914_ ( .A(\wbu.rf_10 [7] ), .B(_13894_ ), .S(_12982_ ), .Z(_13895_ ) );
MUX2_X1 _20915_ ( .A(\wbu.rf_11 [7] ), .B(_13895_ ), .S(_13035_ ), .Z(_13896_ ) );
MUX2_X1 _20916_ ( .A(\wbu.rf_12 [7] ), .B(_13896_ ), .S(_13042_ ), .Z(_13897_ ) );
MUX2_X1 _20917_ ( .A(\wbu.rf_13 [7] ), .B(_13897_ ), .S(_13051_ ), .Z(_13898_ ) );
MUX2_X1 _20918_ ( .A(\wbu.rf_14 [7] ), .B(_13898_ ), .S(_13057_ ), .Z(_13899_ ) );
MUX2_X1 _20919_ ( .A(\wbu.rf_15 [7] ), .B(_13899_ ), .S(_13068_ ), .Z(_13900_ ) );
MUX2_X1 _20920_ ( .A(\wbu.rf_16 [7] ), .B(_13900_ ), .S(_13073_ ), .Z(_13901_ ) );
MUX2_X1 _20921_ ( .A(\wbu.rf_17 [7] ), .B(_13901_ ), .S(_13083_ ), .Z(_13902_ ) );
MUX2_X1 _20922_ ( .A(\wbu.rf_18 [7] ), .B(_13902_ ), .S(_13089_ ), .Z(_13903_ ) );
MUX2_X1 _20923_ ( .A(\wbu.rf_19 [7] ), .B(_13903_ ), .S(_13096_ ), .Z(_13904_ ) );
MUX2_X1 _20924_ ( .A(\wbu.rf_20 [7] ), .B(_13904_ ), .S(_13102_ ), .Z(_13905_ ) );
MUX2_X1 _20925_ ( .A(\wbu.rf_21 [7] ), .B(_13905_ ), .S(_13110_ ), .Z(_13906_ ) );
MUX2_X1 _20926_ ( .A(\wbu.rf_22 [7] ), .B(_13906_ ), .S(_13116_ ), .Z(_13907_ ) );
MUX2_X1 _20927_ ( .A(\wbu.rf_23 [7] ), .B(_13907_ ), .S(_13126_ ), .Z(_13908_ ) );
MUX2_X1 _20928_ ( .A(\wbu.rf_24 [7] ), .B(_13908_ ), .S(_13131_ ), .Z(_13909_ ) );
MUX2_X1 _20929_ ( .A(\wbu.rf_25 [7] ), .B(_13909_ ), .S(_13139_ ), .Z(_13910_ ) );
MUX2_X1 _20930_ ( .A(\wbu.rf_26 [7] ), .B(_13910_ ), .S(_13145_ ), .Z(_13911_ ) );
AOI21_X1 _20931_ ( .A(_13886_ ), .B1(_13911_ ), .B2(_13153_ ), .ZN(_13912_ ) );
OAI211_X1 _20932_ ( .A(_13165_ ), .B(_13885_ ), .C1(_13912_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_13913_ ) );
OAI211_X1 _20933_ ( .A(_13913_ ), .B(_13268_ ), .C1(\wbu.rf_29 [7] ), .C2(_13269_ ), .ZN(_13914_ ) );
NAND4_X1 _20934_ ( .A1(_13272_ ), .A2(fanout_net_33 ), .A3(_13273_ ), .A4(\wbu.rf_30 [7] ), .ZN(_13915_ ) );
NAND3_X1 _20935_ ( .A1(_13914_ ), .A2(_13374_ ), .A3(_13915_ ), .ZN(_13916_ ) );
OR2_X1 _20936_ ( .A1(_13369_ ), .A2(\wbu.rf_31 [7] ), .ZN(_13917_ ) );
AOI21_X1 _20937_ ( .A(_13324_ ), .B1(_13916_ ), .B2(_13917_ ), .ZN(_13918_ ) );
INV_X1 _20938_ ( .A(\wbu.io_in_bits_rd_wdata [7] ), .ZN(_13919_ ) );
AOI211_X1 _20939_ ( .A(fanout_net_24 ), .B(_13918_ ), .C1(_13919_ ), .C2(_13373_ ), .ZN(_00363_ ) );
OR2_X1 _20940_ ( .A1(_13374_ ), .A2(\wbu.rf_31 [6] ), .ZN(_13920_ ) );
NAND4_X1 _20941_ ( .A1(_13092_ ), .A2(fanout_net_33 ), .A3(\wbu.rf_17 [6] ), .A4(_08574_ ), .ZN(_13921_ ) );
AND4_X1 _20942_ ( .A1(fanout_net_33 ), .A2(_08573_ ), .A3(_13228_ ), .A4(\wbu.rf_16 [6] ), .ZN(_13922_ ) );
MUX2_X1 _20943_ ( .A(\wbu._GEN_71 [6] ), .B(\wbu.rf_2 [6] ), .S(_12992_ ), .Z(_13923_ ) );
MUX2_X1 _20944_ ( .A(\wbu.rf_3 [6] ), .B(_13923_ ), .S(_12997_ ), .Z(_13924_ ) );
MUX2_X1 _20945_ ( .A(\wbu.rf_4 [6] ), .B(_13924_ ), .S(_13003_ ), .Z(_13925_ ) );
MUX2_X1 _20946_ ( .A(\wbu.rf_5 [6] ), .B(_13925_ ), .S(_13011_ ), .Z(_13926_ ) );
MUX2_X1 _20947_ ( .A(\wbu.rf_6 [6] ), .B(_13926_ ), .S(_13017_ ), .Z(_13927_ ) );
MUX2_X1 _20948_ ( .A(\wbu.rf_7 [6] ), .B(_13927_ ), .S(_13023_ ), .Z(_13928_ ) );
MUX2_X1 _20949_ ( .A(\wbu.rf_8 [6] ), .B(_13928_ ), .S(_13029_ ), .Z(_13929_ ) );
MUX2_X1 _20950_ ( .A(\wbu.rf_9 [6] ), .B(_13929_ ), .S(_13198_ ), .Z(_13930_ ) );
MUX2_X1 _20951_ ( .A(\wbu.rf_10 [6] ), .B(_13930_ ), .S(_12983_ ), .Z(_00411_ ) );
MUX2_X1 _20952_ ( .A(\wbu.rf_11 [6] ), .B(_00411_ ), .S(_13037_ ), .Z(_00412_ ) );
MUX2_X1 _20953_ ( .A(\wbu.rf_12 [6] ), .B(_00412_ ), .S(_13044_ ), .Z(_00413_ ) );
MUX2_X1 _20954_ ( .A(\wbu.rf_13 [6] ), .B(_00413_ ), .S(_13053_ ), .Z(_00414_ ) );
MUX2_X1 _20955_ ( .A(\wbu.rf_14 [6] ), .B(_00414_ ), .S(_13059_ ), .Z(_00415_ ) );
MUX2_X1 _20956_ ( .A(\wbu.rf_15 [6] ), .B(_00415_ ), .S(_13070_ ), .Z(_00416_ ) );
AOI21_X1 _20957_ ( .A(_13922_ ), .B1(_00416_ ), .B2(_13087_ ), .ZN(_00417_ ) );
OAI211_X1 _20958_ ( .A(_13450_ ), .B(_13921_ ), .C1(_00417_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_00418_ ) );
OAI211_X1 _20959_ ( .A(_00418_ ), .B(_13098_ ), .C1(\wbu.rf_18 [6] ), .C2(_13099_ ), .ZN(_00419_ ) );
NAND4_X1 _20960_ ( .A1(_13106_ ), .A2(_08575_ ), .A3(fanout_net_33 ), .A4(\wbu.rf_19 [6] ), .ZN(_00420_ ) );
NAND3_X1 _20961_ ( .A1(_00419_ ), .A2(_13381_ ), .A3(_00420_ ), .ZN(_00421_ ) );
OAI211_X1 _20962_ ( .A(_00421_ ), .B(_13112_ ), .C1(\wbu.rf_20 [6] ), .C2(_13113_ ), .ZN(_00422_ ) );
NAND4_X1 _20963_ ( .A1(_13120_ ), .A2(_13122_ ), .A3(fanout_net_33 ), .A4(\wbu.rf_21 [6] ), .ZN(_00423_ ) );
NAND3_X1 _20964_ ( .A1(_00422_ ), .A2(_13118_ ), .A3(_00423_ ), .ZN(_00424_ ) );
OAI211_X1 _20965_ ( .A(_00424_ ), .B(_13231_ ), .C1(\wbu.rf_22 [6] ), .C2(_13128_ ), .ZN(_00425_ ) );
NAND4_X1 _20966_ ( .A1(_13133_ ), .A2(fanout_net_33 ), .A3(_13135_ ), .A4(\wbu.rf_23 [6] ), .ZN(_00426_ ) );
NAND3_X1 _20967_ ( .A1(_00425_ ), .A2(_13414_ ), .A3(_00426_ ), .ZN(_00427_ ) );
OAI211_X1 _20968_ ( .A(_00427_ ), .B(_13140_ ), .C1(\wbu.rf_24 [6] ), .C2(_13141_ ), .ZN(_00428_ ) );
NAND4_X1 _20969_ ( .A1(_13147_ ), .A2(_13158_ ), .A3(fanout_net_33 ), .A4(\wbu.rf_25 [6] ), .ZN(_00429_ ) );
NAND3_X1 _20970_ ( .A1(_00428_ ), .A2(_13260_ ), .A3(_00429_ ), .ZN(_00430_ ) );
OAI211_X1 _20971_ ( .A(_00430_ ), .B(_13153_ ), .C1(\wbu.rf_26 [6] ), .C2(_13154_ ), .ZN(_00431_ ) );
NAND4_X1 _20972_ ( .A1(_13159_ ), .A2(fanout_net_33 ), .A3(_13161_ ), .A4(\wbu.rf_27 [6] ), .ZN(_00432_ ) );
NAND3_X1 _20973_ ( .A1(_00431_ ), .A2(_13365_ ), .A3(_00432_ ), .ZN(_00433_ ) );
OAI211_X1 _20974_ ( .A(_00433_ ), .B(_13165_ ), .C1(\wbu.rf_28 [6] ), .C2(_13167_ ), .ZN(_00434_ ) );
NAND4_X1 _20975_ ( .A1(_13169_ ), .A2(fanout_net_33 ), .A3(_13170_ ), .A4(\wbu.rf_29 [6] ), .ZN(_00435_ ) );
NAND2_X1 _20976_ ( .A1(_00434_ ), .A2(_00435_ ), .ZN(_00436_ ) );
MUX2_X1 _20977_ ( .A(\wbu.rf_30 [6] ), .B(_00436_ ), .S(_13268_ ), .Z(_00437_ ) );
OAI211_X1 _20978_ ( .A(_13276_ ), .B(_13920_ ), .C1(_00437_ ), .C2(_13179_ ), .ZN(_00438_ ) );
NAND3_X1 _20979_ ( .A1(_13181_ ), .A2(\wbu.io_in_bits_rd_wdata [6] ), .A3(_13183_ ), .ZN(_00439_ ) );
AOI21_X1 _20980_ ( .A(fanout_net_24 ), .B1(_00438_ ), .B2(_00439_ ), .ZN(_00364_ ) );
OR2_X1 _20981_ ( .A1(_13153_ ), .A2(\wbu.rf_27 [5] ), .ZN(_00440_ ) );
OR2_X1 _20982_ ( .A1(_13030_ ), .A2(\wbu.rf_8 [5] ), .ZN(_00441_ ) );
MUX2_X1 _20983_ ( .A(\wbu._GEN_71 [5] ), .B(\wbu.rf_2 [5] ), .S(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .Z(_00442_ ) );
MUX2_X1 _20984_ ( .A(\wbu.rf_3 [5] ), .B(_00442_ ), .S(_12998_ ), .Z(_00443_ ) );
MUX2_X1 _20985_ ( .A(\wbu.rf_4 [5] ), .B(_00443_ ), .S(_13004_ ), .Z(_00444_ ) );
MUX2_X1 _20986_ ( .A(\wbu.rf_5 [5] ), .B(_00444_ ), .S(_13012_ ), .Z(_00445_ ) );
MUX2_X1 _20987_ ( .A(\wbu.rf_6 [5] ), .B(_00445_ ), .S(_13018_ ), .Z(_00446_ ) );
MUX2_X1 _20988_ ( .A(\wbu.rf_7 [5] ), .B(_00446_ ), .S(_13024_ ), .Z(_00447_ ) );
OAI211_X1 _20989_ ( .A(_13383_ ), .B(_00441_ ), .C1(_00447_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_Y ), .ZN(_00448_ ) );
NAND4_X1 _20990_ ( .A1(_12985_ ), .A2(_12986_ ), .A3(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A4(\wbu.rf_9 [5] ), .ZN(_00449_ ) );
NAND3_X1 _20991_ ( .A1(_00448_ ), .A2(_12984_ ), .A3(_00449_ ), .ZN(_00450_ ) );
OAI211_X1 _20992_ ( .A(_00450_ ), .B(_13038_ ), .C1(\wbu.rf_10 [5] ), .C2(_13039_ ), .ZN(_00451_ ) );
NAND4_X1 _20993_ ( .A1(_13046_ ), .A2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A3(_13047_ ), .A4(\wbu.rf_11 [5] ), .ZN(_00452_ ) );
NAND3_X1 _20994_ ( .A1(_00451_ ), .A2(_13045_ ), .A3(_00452_ ), .ZN(_00453_ ) );
OAI211_X1 _20995_ ( .A(_00453_ ), .B(_13054_ ), .C1(\wbu.rf_12 [5] ), .C2(_13055_ ), .ZN(_00454_ ) );
NAND4_X1 _20996_ ( .A1(_13061_ ), .A2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A3(_13064_ ), .A4(\wbu.rf_13 [5] ), .ZN(_00455_ ) );
NAND3_X1 _20997_ ( .A1(_00454_ ), .A2(_13059_ ), .A3(_00455_ ), .ZN(_00456_ ) );
OAI211_X1 _20998_ ( .A(_00456_ ), .B(_13070_ ), .C1(\wbu.rf_14 [5] ), .C2(_13060_ ), .ZN(_00457_ ) );
NAND4_X1 _20999_ ( .A1(_13077_ ), .A2(_13078_ ), .A3(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A4(\wbu.rf_15 [5] ), .ZN(_00458_ ) );
NAND3_X1 _21000_ ( .A1(_00457_ ), .A2(_13075_ ), .A3(_00458_ ), .ZN(_00459_ ) );
OAI211_X1 _21001_ ( .A(_00459_ ), .B(_13085_ ), .C1(\wbu.rf_16 [5] ), .C2(_13076_ ), .ZN(_00460_ ) );
NAND4_X1 _21002_ ( .A1(_13092_ ), .A2(fanout_net_33 ), .A3(\wbu.rf_17 [5] ), .A4(_13350_ ), .ZN(_00461_ ) );
NAND3_X1 _21003_ ( .A1(_00460_ ), .A2(_13091_ ), .A3(_00461_ ), .ZN(_00462_ ) );
OAI211_X1 _21004_ ( .A(_00462_ ), .B(_13097_ ), .C1(\wbu.rf_18 [5] ), .C2(_13450_ ), .ZN(_00463_ ) );
NAND4_X1 _21005_ ( .A1(_13105_ ), .A2(_13497_ ), .A3(fanout_net_33 ), .A4(\wbu.rf_19 [5] ), .ZN(_00464_ ) );
NAND3_X1 _21006_ ( .A1(_00463_ ), .A2(_13103_ ), .A3(_00464_ ), .ZN(_00465_ ) );
OAI211_X1 _21007_ ( .A(_00465_ ), .B(_13111_ ), .C1(\wbu.rf_20 [5] ), .C2(_13381_ ), .ZN(_00466_ ) );
NAND4_X1 _21008_ ( .A1(_13119_ ), .A2(_13188_ ), .A3(fanout_net_34 ), .A4(\wbu.rf_21 [5] ), .ZN(_00467_ ) );
NAND3_X1 _21009_ ( .A1(_00466_ ), .A2(_13117_ ), .A3(_00467_ ), .ZN(_00468_ ) );
OAI211_X1 _21010_ ( .A(_00468_ ), .B(_13127_ ), .C1(\wbu.rf_22 [5] ), .C2(_13212_ ), .ZN(_00469_ ) );
NAND4_X1 _21011_ ( .A1(_13186_ ), .A2(fanout_net_34 ), .A3(_13134_ ), .A4(\wbu.rf_23 [5] ), .ZN(_00470_ ) );
NAND3_X1 _21012_ ( .A1(_00469_ ), .A2(_13132_ ), .A3(_00470_ ), .ZN(_00471_ ) );
OAI211_X1 _21013_ ( .A(_00471_ ), .B(_13460_ ), .C1(\wbu.rf_24 [5] ), .C2(_13414_ ), .ZN(_00472_ ) );
NAND4_X1 _21014_ ( .A1(_13312_ ), .A2(_13378_ ), .A3(fanout_net_34 ), .A4(\wbu.rf_25 [5] ), .ZN(_00473_ ) );
NAND2_X1 _21015_ ( .A1(_00472_ ), .A2(_00473_ ), .ZN(_00474_ ) );
MUX2_X1 _21016_ ( .A(\wbu.rf_26 [5] ), .B(_00474_ ), .S(_13260_ ), .Z(_00475_ ) );
OAI211_X1 _21017_ ( .A(_13365_ ), .B(_00440_ ), .C1(_00475_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .ZN(_00476_ ) );
NAND4_X1 _21018_ ( .A1(_13376_ ), .A2(_13229_ ), .A3(fanout_net_34 ), .A4(\wbu.rf_28 [5] ), .ZN(_00477_ ) );
AOI21_X1 _21019_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .B1(_00476_ ), .B2(_00477_ ), .ZN(_00478_ ) );
NAND3_X1 _21020_ ( .A1(_13050_ ), .A2(fanout_net_34 ), .A3(\wbu.rf_29 [5] ), .ZN(_00479_ ) );
NAND2_X1 _21021_ ( .A1(_13267_ ), .A2(_00479_ ), .ZN(_00480_ ) );
OAI221_X1 _21022_ ( .A(_12970_ ), .B1(\wbu.rf_30 [5] ), .B2(_13268_ ), .C1(_00478_ ), .C2(_00480_ ), .ZN(_00481_ ) );
NAND4_X1 _21023_ ( .A1(_13161_ ), .A2(_13273_ ), .A3(fanout_net_34 ), .A4(\wbu.rf_31 [5] ), .ZN(_00482_ ) );
AND3_X1 _21024_ ( .A1(_00481_ ), .A2(_13276_ ), .A3(_00482_ ), .ZN(_00483_ ) );
INV_X1 _21025_ ( .A(\wbu.io_in_bits_rd_wdata [5] ), .ZN(_00484_ ) );
AOI211_X1 _21026_ ( .A(fanout_net_24 ), .B(_00483_ ), .C1(_00484_ ), .C2(_13373_ ), .ZN(_00365_ ) );
INV_X1 _21027_ ( .A(\wbu.io_in_bits_rd_wdata [4] ), .ZN(_00485_ ) );
NAND4_X1 _21028_ ( .A1(_13046_ ), .A2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A3(_12966_ ), .A4(\wbu.rf_11 [4] ), .ZN(_00486_ ) );
AND4_X1 _21029_ ( .A1(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A2(_12977_ ), .A3(_12986_ ), .A4(\wbu.rf_10 [4] ), .ZN(_00487_ ) );
MUX2_X1 _21030_ ( .A(\wbu._GEN_71 [4] ), .B(\wbu.rf_2 [4] ), .S(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .Z(_00488_ ) );
MUX2_X1 _21031_ ( .A(\wbu.rf_3 [4] ), .B(_00488_ ), .S(_12998_ ), .Z(_00489_ ) );
MUX2_X1 _21032_ ( .A(\wbu.rf_4 [4] ), .B(_00489_ ), .S(_13004_ ), .Z(_00490_ ) );
MUX2_X1 _21033_ ( .A(\wbu.rf_5 [4] ), .B(_00490_ ), .S(_13012_ ), .Z(_00491_ ) );
MUX2_X1 _21034_ ( .A(\wbu.rf_6 [4] ), .B(_00491_ ), .S(_13018_ ), .Z(_00492_ ) );
MUX2_X1 _21035_ ( .A(\wbu.rf_7 [4] ), .B(_00492_ ), .S(_13024_ ), .Z(_00493_ ) );
MUX2_X1 _21036_ ( .A(\wbu.rf_8 [4] ), .B(_00493_ ), .S(_13030_ ), .Z(_00494_ ) );
MUX2_X1 _21037_ ( .A(\wbu.rf_9 [4] ), .B(_00494_ ), .S(_13383_ ), .Z(_00495_ ) );
AOI21_X1 _21038_ ( .A(_00487_ ), .B1(_00495_ ), .B2(_13039_ ), .ZN(_00496_ ) );
OAI211_X1 _21039_ ( .A(_13045_ ), .B(_00486_ ), .C1(_00496_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .ZN(_00497_ ) );
OAI211_X1 _21040_ ( .A(_00497_ ), .B(_13054_ ), .C1(\wbu.rf_12 [4] ), .C2(_13055_ ), .ZN(_00498_ ) );
NAND4_X1 _21041_ ( .A1(_13061_ ), .A2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A3(_13064_ ), .A4(\wbu.rf_13 [4] ), .ZN(_00499_ ) );
NAND3_X1 _21042_ ( .A1(_00498_ ), .A2(_13059_ ), .A3(_00499_ ), .ZN(_00500_ ) );
OAI211_X1 _21043_ ( .A(_00500_ ), .B(_13070_ ), .C1(\wbu.rf_14 [4] ), .C2(_13071_ ), .ZN(_00501_ ) );
NAND4_X1 _21044_ ( .A1(_13077_ ), .A2(_13078_ ), .A3(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A4(\wbu.rf_15 [4] ), .ZN(_00502_ ) );
NAND3_X1 _21045_ ( .A1(_00501_ ), .A2(_13076_ ), .A3(_00502_ ), .ZN(_00503_ ) );
OAI211_X1 _21046_ ( .A(_00503_ ), .B(_13085_ ), .C1(\wbu.rf_16 [4] ), .C2(_13087_ ), .ZN(_00504_ ) );
NAND4_X1 _21047_ ( .A1(_13092_ ), .A2(fanout_net_34 ), .A3(\wbu.rf_17 [4] ), .A4(_13350_ ), .ZN(_00505_ ) );
NAND3_X1 _21048_ ( .A1(_00504_ ), .A2(_13091_ ), .A3(_00505_ ), .ZN(_00506_ ) );
OAI211_X1 _21049_ ( .A(_00506_ ), .B(_13097_ ), .C1(\wbu.rf_18 [4] ), .C2(_13450_ ), .ZN(_00507_ ) );
NAND4_X1 _21050_ ( .A1(_13106_ ), .A2(_13497_ ), .A3(fanout_net_34 ), .A4(\wbu.rf_19 [4] ), .ZN(_00508_ ) );
NAND3_X1 _21051_ ( .A1(_00507_ ), .A2(_13104_ ), .A3(_00508_ ), .ZN(_00509_ ) );
OAI211_X1 _21052_ ( .A(_00509_ ), .B(_13111_ ), .C1(\wbu.rf_20 [4] ), .C2(_13381_ ), .ZN(_00510_ ) );
NAND4_X1 _21053_ ( .A1(_13120_ ), .A2(_13188_ ), .A3(fanout_net_34 ), .A4(\wbu.rf_21 [4] ), .ZN(_00511_ ) );
NAND3_X1 _21054_ ( .A1(_00510_ ), .A2(_13118_ ), .A3(_00511_ ), .ZN(_00512_ ) );
OAI211_X1 _21055_ ( .A(_00512_ ), .B(_13127_ ), .C1(\wbu.rf_22 [4] ), .C2(_13212_ ), .ZN(_00513_ ) );
NAND4_X1 _21056_ ( .A1(_13133_ ), .A2(fanout_net_34 ), .A3(_13135_ ), .A4(\wbu.rf_23 [4] ), .ZN(_00514_ ) );
NAND3_X1 _21057_ ( .A1(_00513_ ), .A2(_13132_ ), .A3(_00514_ ), .ZN(_00515_ ) );
OAI211_X1 _21058_ ( .A(_00515_ ), .B(_13460_ ), .C1(\wbu.rf_24 [4] ), .C2(_13414_ ), .ZN(_00516_ ) );
NAND4_X1 _21059_ ( .A1(_13312_ ), .A2(_13149_ ), .A3(fanout_net_34 ), .A4(\wbu.rf_25 [4] ), .ZN(_00517_ ) );
NAND3_X1 _21060_ ( .A1(_00516_ ), .A2(_13144_ ), .A3(_00517_ ), .ZN(_00518_ ) );
OAI211_X1 _21061_ ( .A(_00518_ ), .B(_13218_ ), .C1(\wbu.rf_26 [4] ), .C2(_13260_ ), .ZN(_00519_ ) );
NAND4_X1 _21062_ ( .A1(_13158_ ), .A2(fanout_net_34 ), .A3(_13160_ ), .A4(\wbu.rf_27 [4] ), .ZN(_00520_ ) );
NAND3_X1 _21063_ ( .A1(_00519_ ), .A2(_13166_ ), .A3(_00520_ ), .ZN(_00521_ ) );
OAI211_X1 _21064_ ( .A(_00521_ ), .B(_13512_ ), .C1(\wbu.rf_28 [4] ), .C2(_13365_ ), .ZN(_00522_ ) );
NAND4_X1 _21065_ ( .A1(_13326_ ), .A2(fanout_net_34 ), .A3(_13176_ ), .A4(\wbu.rf_29 [4] ), .ZN(_00523_ ) );
AOI21_X1 _21066_ ( .A(_12975_ ), .B1(_00522_ ), .B2(_00523_ ), .ZN(_00524_ ) );
AND4_X1 _21067_ ( .A1(fanout_net_34 ), .A2(_13175_ ), .A3(\wbu.rf_30 [4] ), .A4(_13376_ ), .ZN(_00525_ ) );
OAI21_X1 _21068_ ( .A(_13369_ ), .B1(_00524_ ), .B2(_00525_ ), .ZN(_00526_ ) );
AOI22_X1 _21069_ ( .A1(_12969_ ), .A2(\wbu.rf_31 [4] ), .B1(_13180_ ), .B2(_13182_ ), .ZN(_00527_ ) );
AOI221_X4 _21070_ ( .A(fanout_net_25 ), .B1(_00485_ ), .B2(_12965_ ), .C1(_00526_ ), .C2(_00527_ ), .ZN(_00366_ ) );
NAND4_X1 _21071_ ( .A1(_13272_ ), .A2(fanout_net_34 ), .A3(_13273_ ), .A4(\wbu.rf_30 [3] ), .ZN(_00528_ ) );
AND4_X1 _21072_ ( .A1(fanout_net_34 ), .A2(_13147_ ), .A3(\wbu.rf_29 [3] ), .A4(_13327_ ), .ZN(_00529_ ) );
NOR2_X1 _21073_ ( .A1(_13110_ ), .A2(\wbu.rf_21 [3] ), .ZN(_00530_ ) );
OAI21_X1 _21074_ ( .A(_13102_ ), .B1(_13096_ ), .B2(\wbu.rf_19 [3] ), .ZN(_00531_ ) );
INV_X1 _21075_ ( .A(_00531_ ), .ZN(_00532_ ) );
NAND3_X1 _21076_ ( .A1(_13026_ ), .A2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A3(\wbu.rf_8 [3] ), .ZN(_00533_ ) );
AND4_X1 _21077_ ( .A1(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A2(_12977_ ), .A3(_13007_ ), .A4(\wbu.rf_6 [3] ), .ZN(_00534_ ) );
MUX2_X1 _21078_ ( .A(\wbu._GEN_71 [3] ), .B(\wbu.rf_2 [3] ), .S(_12991_ ), .Z(_00535_ ) );
MUX2_X1 _21079_ ( .A(\wbu.rf_3 [3] ), .B(_00535_ ), .S(_12996_ ), .Z(_00536_ ) );
MUX2_X1 _21080_ ( .A(\wbu.rf_4 [3] ), .B(_00536_ ), .S(_13002_ ), .Z(_00537_ ) );
MUX2_X1 _21081_ ( .A(\wbu.rf_5 [3] ), .B(_00537_ ), .S(_13010_ ), .Z(_00538_ ) );
AOI211_X1 _21082_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_Y ), .B(_00534_ ), .C1(_00538_ ), .C2(_13016_ ), .ZN(_00539_ ) );
OAI21_X1 _21083_ ( .A(_13027_ ), .B1(_13022_ ), .B2(\wbu.rf_7 [3] ), .ZN(_00540_ ) );
OAI21_X1 _21084_ ( .A(_00533_ ), .B1(_00539_ ), .B2(_00540_ ), .ZN(_00541_ ) );
MUX2_X1 _21085_ ( .A(\wbu.rf_9 [3] ), .B(_00541_ ), .S(_13197_ ), .Z(_00542_ ) );
MUX2_X1 _21086_ ( .A(\wbu.rf_10 [3] ), .B(_00542_ ), .S(_12982_ ), .Z(_00543_ ) );
MUX2_X1 _21087_ ( .A(\wbu.rf_11 [3] ), .B(_00543_ ), .S(_13036_ ), .Z(_00544_ ) );
MUX2_X1 _21088_ ( .A(\wbu.rf_12 [3] ), .B(_00544_ ), .S(_13043_ ), .Z(_00545_ ) );
MUX2_X1 _21089_ ( .A(\wbu.rf_13 [3] ), .B(_00545_ ), .S(_13052_ ), .Z(_00546_ ) );
MUX2_X1 _21090_ ( .A(\wbu.rf_14 [3] ), .B(_00546_ ), .S(_13057_ ), .Z(_00547_ ) );
MUX2_X1 _21091_ ( .A(\wbu.rf_15 [3] ), .B(_00547_ ), .S(_13068_ ), .Z(_00548_ ) );
MUX2_X1 _21092_ ( .A(\wbu.rf_16 [3] ), .B(_00548_ ), .S(_13074_ ), .Z(_00549_ ) );
MUX2_X1 _21093_ ( .A(\wbu.rf_17 [3] ), .B(_00549_ ), .S(_13084_ ), .Z(_00550_ ) );
MUX2_X1 _21094_ ( .A(\wbu.rf_18 [3] ), .B(_00550_ ), .S(_13090_ ), .Z(_00551_ ) );
OAI21_X1 _21095_ ( .A(_00532_ ), .B1(_00551_ ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .ZN(_00552_ ) );
AOI22_X1 _21096_ ( .A1(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .A2(\wbu.rf_20 [3] ), .B1(fanout_net_34 ), .B2(_13008_ ), .ZN(_00553_ ) );
AOI21_X1 _21097_ ( .A(_00530_ ), .B1(_00552_ ), .B2(_00553_ ), .ZN(_00554_ ) );
MUX2_X1 _21098_ ( .A(\wbu.rf_22 [3] ), .B(_00554_ ), .S(_13116_ ), .Z(_00555_ ) );
MUX2_X1 _21099_ ( .A(\wbu.rf_23 [3] ), .B(_00555_ ), .S(_13126_ ), .Z(_00556_ ) );
MUX2_X1 _21100_ ( .A(\wbu.rf_24 [3] ), .B(_00556_ ), .S(_13130_ ), .Z(_00557_ ) );
MUX2_X1 _21101_ ( .A(\wbu.rf_25 [3] ), .B(_00557_ ), .S(_13139_ ), .Z(_00558_ ) );
MUX2_X1 _21102_ ( .A(\wbu.rf_26 [3] ), .B(_00558_ ), .S(_13143_ ), .Z(_00559_ ) );
MUX2_X1 _21103_ ( .A(\wbu.rf_27 [3] ), .B(_00559_ ), .S(_13363_ ), .Z(_00560_ ) );
MUX2_X1 _21104_ ( .A(\wbu.rf_28 [3] ), .B(_00560_ ), .S(_13157_ ), .Z(_00561_ ) );
AOI21_X1 _21105_ ( .A(_00529_ ), .B1(_00561_ ), .B2(_13269_ ), .ZN(_00562_ ) );
OAI211_X1 _21106_ ( .A(_12971_ ), .B(_00528_ ), .C1(_00562_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_00563_ ) );
OR2_X1 _21107_ ( .A1(_13369_ ), .A2(\wbu.rf_31 [3] ), .ZN(_00564_ ) );
AOI21_X1 _21108_ ( .A(_13324_ ), .B1(_00563_ ), .B2(_00564_ ), .ZN(_00565_ ) );
INV_X1 _21109_ ( .A(\wbu.io_in_bits_rd_wdata [3] ), .ZN(_00566_ ) );
AOI211_X1 _21110_ ( .A(fanout_net_25 ), .B(_00565_ ), .C1(_00566_ ), .C2(_13373_ ), .ZN(_00367_ ) );
OR2_X1 _21111_ ( .A1(_12971_ ), .A2(\wbu.rf_31 [2] ), .ZN(_00567_ ) );
NAND3_X1 _21112_ ( .A1(_12961_ ), .A2(fanout_net_34 ), .A3(\wbu.rf_16 [2] ), .ZN(_00568_ ) );
AND3_X1 _21113_ ( .A1(_12973_ ), .A2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A3(\wbu.rf_14 [2] ), .ZN(_00569_ ) );
NAND3_X1 _21114_ ( .A1(_13032_ ), .A2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A3(\wbu.rf_9 [2] ), .ZN(_00570_ ) );
AND4_X1 _21115_ ( .A1(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A2(_12979_ ), .A3(\wbu.rf_8 [2] ), .A4(_12959_ ), .ZN(_00571_ ) );
OR2_X1 _21116_ ( .A1(_13010_ ), .A2(\wbu.rf_5 [2] ), .ZN(_00572_ ) );
MUX2_X1 _21117_ ( .A(\wbu._GEN_71 [2] ), .B(\wbu.rf_2 [2] ), .S(_12991_ ), .Z(_00573_ ) );
MUX2_X1 _21118_ ( .A(\wbu.rf_3 [2] ), .B(_00573_ ), .S(_12996_ ), .Z(_00574_ ) );
MUX2_X1 _21119_ ( .A(\wbu.rf_4 [2] ), .B(_00574_ ), .S(_13002_ ), .Z(_00575_ ) );
OAI211_X1 _21120_ ( .A(_13016_ ), .B(_00572_ ), .C1(_00575_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_00576_ ) );
NAND4_X1 _21121_ ( .A1(_12977_ ), .A2(_13007_ ), .A3(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A4(\wbu.rf_6 [2] ), .ZN(_00577_ ) );
NAND3_X1 _21122_ ( .A1(_00576_ ), .A2(_13022_ ), .A3(_00577_ ), .ZN(_00578_ ) );
NOR2_X1 _21123_ ( .A1(_13021_ ), .A2(\wbu.rf_7 [2] ), .ZN(_00579_ ) );
NOR2_X1 _21124_ ( .A1(_00579_ ), .A2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_Y ), .ZN(_00580_ ) );
AOI21_X1 _21125_ ( .A(_00571_ ), .B1(_00578_ ), .B2(_00580_ ), .ZN(_00581_ ) );
OAI21_X1 _21126_ ( .A(_00570_ ), .B1(_00581_ ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_Y ), .ZN(_00582_ ) );
MUX2_X1 _21127_ ( .A(\wbu.rf_10 [2] ), .B(_00582_ ), .S(_12982_ ), .Z(_00583_ ) );
MUX2_X1 _21128_ ( .A(\wbu.rf_11 [2] ), .B(_00583_ ), .S(_13036_ ), .Z(_00584_ ) );
MUX2_X1 _21129_ ( .A(\wbu.rf_12 [2] ), .B(_00584_ ), .S(_13043_ ), .Z(_00585_ ) );
MUX2_X1 _21130_ ( .A(\wbu.rf_13 [2] ), .B(_00585_ ), .S(_13052_ ), .Z(_00586_ ) );
AOI211_X1 _21131_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .B(_00569_ ), .C1(_00586_ ), .C2(_13057_ ), .ZN(_00587_ ) );
OAI21_X1 _21132_ ( .A(_13073_ ), .B1(_13068_ ), .B2(\wbu.rf_15 [2] ), .ZN(_00588_ ) );
OAI21_X1 _21133_ ( .A(_00568_ ), .B1(_00587_ ), .B2(_00588_ ), .ZN(_00589_ ) );
MUX2_X1 _21134_ ( .A(\wbu.rf_17 [2] ), .B(_00589_ ), .S(_13083_ ), .Z(_00590_ ) );
MUX2_X1 _21135_ ( .A(\wbu.rf_18 [2] ), .B(_00590_ ), .S(_13089_ ), .Z(_00591_ ) );
MUX2_X1 _21136_ ( .A(\wbu.rf_19 [2] ), .B(_00591_ ), .S(_13096_ ), .Z(_00592_ ) );
MUX2_X1 _21137_ ( .A(\wbu.rf_20 [2] ), .B(_00592_ ), .S(_13101_ ), .Z(_00593_ ) );
MUX2_X1 _21138_ ( .A(\wbu.rf_21 [2] ), .B(_00593_ ), .S(_13110_ ), .Z(_00594_ ) );
MUX2_X1 _21139_ ( .A(\wbu.rf_22 [2] ), .B(_00594_ ), .S(_13115_ ), .Z(_00595_ ) );
MUX2_X1 _21140_ ( .A(\wbu.rf_23 [2] ), .B(_00595_ ), .S(_13126_ ), .Z(_00596_ ) );
MUX2_X1 _21141_ ( .A(\wbu.rf_24 [2] ), .B(_00596_ ), .S(_13130_ ), .Z(_00597_ ) );
MUX2_X1 _21142_ ( .A(\wbu.rf_25 [2] ), .B(_00597_ ), .S(_13139_ ), .Z(_00598_ ) );
MUX2_X1 _21143_ ( .A(\wbu.rf_26 [2] ), .B(_00598_ ), .S(_13143_ ), .Z(_00599_ ) );
MUX2_X1 _21144_ ( .A(\wbu.rf_27 [2] ), .B(_00599_ ), .S(_13152_ ), .Z(_00600_ ) );
MUX2_X1 _21145_ ( .A(\wbu.rf_28 [2] ), .B(_00600_ ), .S(_13156_ ), .Z(_00601_ ) );
MUX2_X1 _21146_ ( .A(\wbu.rf_29 [2] ), .B(_00601_ ), .S(_13512_ ), .Z(_00602_ ) );
MUX2_X1 _21147_ ( .A(\wbu.rf_30 [2] ), .B(_00602_ ), .S(_13268_ ), .Z(_00603_ ) );
OAI211_X1 _21148_ ( .A(_13276_ ), .B(_00567_ ), .C1(_00603_ ), .C2(_13179_ ), .ZN(_00604_ ) );
NAND3_X1 _21149_ ( .A1(_13181_ ), .A2(\wbu.io_in_bits_rd_wdata [2] ), .A3(_13183_ ), .ZN(_00605_ ) );
AOI21_X1 _21150_ ( .A(fanout_net_25 ), .B1(_00604_ ), .B2(_00605_ ), .ZN(_00368_ ) );
AND3_X1 _21151_ ( .A1(_13474_ ), .A2(fanout_net_34 ), .A3(\wbu.rf_31 [28] ), .ZN(_00606_ ) );
NAND4_X1 _21152_ ( .A1(_13272_ ), .A2(fanout_net_34 ), .A3(_13170_ ), .A4(\wbu.rf_30 [28] ), .ZN(_00607_ ) );
AND4_X1 _21153_ ( .A1(fanout_net_34 ), .A2(_13147_ ), .A3(\wbu.rf_29 [28] ), .A4(_13327_ ), .ZN(_00608_ ) );
MUX2_X1 _21154_ ( .A(\wbu._GEN_71 [28] ), .B(\wbu.rf_2 [28] ), .S(_12990_ ), .Z(_00609_ ) );
MUX2_X1 _21155_ ( .A(\wbu.rf_3 [28] ), .B(_00609_ ), .S(_12995_ ), .Z(_00610_ ) );
MUX2_X1 _21156_ ( .A(\wbu.rf_4 [28] ), .B(_00610_ ), .S(_13001_ ), .Z(_00611_ ) );
MUX2_X1 _21157_ ( .A(\wbu.rf_5 [28] ), .B(_00611_ ), .S(_13009_ ), .Z(_00612_ ) );
MUX2_X1 _21158_ ( .A(\wbu.rf_6 [28] ), .B(_00612_ ), .S(_13015_ ), .Z(_00613_ ) );
MUX2_X1 _21159_ ( .A(\wbu.rf_7 [28] ), .B(_00613_ ), .S(_13021_ ), .Z(_00614_ ) );
MUX2_X1 _21160_ ( .A(\wbu.rf_8 [28] ), .B(_00614_ ), .S(_13027_ ), .Z(_00615_ ) );
MUX2_X1 _21161_ ( .A(\wbu.rf_9 [28] ), .B(_00615_ ), .S(_13197_ ), .Z(_00616_ ) );
MUX2_X1 _21162_ ( .A(\wbu.rf_10 [28] ), .B(_00616_ ), .S(_12981_ ), .Z(_00617_ ) );
MUX2_X1 _21163_ ( .A(\wbu.rf_11 [28] ), .B(_00617_ ), .S(_13035_ ), .Z(_00618_ ) );
MUX2_X1 _21164_ ( .A(\wbu.rf_12 [28] ), .B(_00618_ ), .S(_13042_ ), .Z(_00619_ ) );
MUX2_X1 _21165_ ( .A(\wbu.rf_13 [28] ), .B(_00619_ ), .S(_13051_ ), .Z(_00620_ ) );
MUX2_X1 _21166_ ( .A(\wbu.rf_14 [28] ), .B(_00620_ ), .S(_13057_ ), .Z(_00621_ ) );
MUX2_X1 _21167_ ( .A(\wbu.rf_15 [28] ), .B(_00621_ ), .S(_13067_ ), .Z(_00622_ ) );
MUX2_X1 _21168_ ( .A(\wbu.rf_16 [28] ), .B(_00622_ ), .S(_13073_ ), .Z(_00623_ ) );
MUX2_X1 _21169_ ( .A(\wbu.rf_17 [28] ), .B(_00623_ ), .S(_13083_ ), .Z(_00624_ ) );
MUX2_X1 _21170_ ( .A(\wbu.rf_18 [28] ), .B(_00624_ ), .S(_13089_ ), .Z(_00625_ ) );
MUX2_X1 _21171_ ( .A(\wbu.rf_19 [28] ), .B(_00625_ ), .S(_13096_ ), .Z(_00626_ ) );
MUX2_X1 _21172_ ( .A(\wbu.rf_20 [28] ), .B(_00626_ ), .S(_13102_ ), .Z(_00627_ ) );
MUX2_X1 _21173_ ( .A(\wbu.rf_21 [28] ), .B(_00627_ ), .S(_13110_ ), .Z(_00628_ ) );
MUX2_X1 _21174_ ( .A(\wbu.rf_22 [28] ), .B(_00628_ ), .S(_13116_ ), .Z(_00629_ ) );
MUX2_X1 _21175_ ( .A(\wbu.rf_23 [28] ), .B(_00629_ ), .S(_13126_ ), .Z(_00630_ ) );
MUX2_X1 _21176_ ( .A(\wbu.rf_24 [28] ), .B(_00630_ ), .S(_13130_ ), .Z(_00631_ ) );
MUX2_X1 _21177_ ( .A(\wbu.rf_25 [28] ), .B(_00631_ ), .S(_13139_ ), .Z(_00632_ ) );
MUX2_X1 _21178_ ( .A(\wbu.rf_26 [28] ), .B(_00632_ ), .S(_13143_ ), .Z(_00633_ ) );
MUX2_X1 _21179_ ( .A(\wbu.rf_27 [28] ), .B(_00633_ ), .S(_13363_ ), .Z(_00634_ ) );
MUX2_X1 _21180_ ( .A(\wbu.rf_28 [28] ), .B(_00634_ ), .S(_13166_ ), .Z(_00635_ ) );
AOI21_X1 _21181_ ( .A(_00608_ ), .B1(_00635_ ), .B2(_13269_ ), .ZN(_00636_ ) );
OAI21_X1 _21182_ ( .A(_00607_ ), .B1(_00636_ ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_00637_ ) );
AOI211_X1 _21183_ ( .A(_13473_ ), .B(_00606_ ), .C1(_00637_ ), .C2(_13374_ ), .ZN(_00638_ ) );
INV_X1 _21184_ ( .A(\wbu.io_in_bits_rd_wdata [28] ), .ZN(_00639_ ) );
AOI211_X1 _21185_ ( .A(fanout_net_25 ), .B(_00638_ ), .C1(_00639_ ), .C2(_13373_ ), .ZN(_00369_ ) );
INV_X1 _21186_ ( .A(\wbu.io_in_bits_rd_wdata [1] ), .ZN(_00640_ ) );
OR2_X1 _21187_ ( .A1(_13090_ ), .A2(\wbu.rf_18 [1] ), .ZN(_00641_ ) );
MUX2_X1 _21188_ ( .A(\wbu._GEN_71 [1] ), .B(\wbu.rf_2 [1] ), .S(_12991_ ), .Z(_00642_ ) );
MUX2_X1 _21189_ ( .A(\wbu.rf_3 [1] ), .B(_00642_ ), .S(_12996_ ), .Z(_00643_ ) );
MUX2_X1 _21190_ ( .A(\wbu.rf_4 [1] ), .B(_00643_ ), .S(_13002_ ), .Z(_00644_ ) );
MUX2_X1 _21191_ ( .A(\wbu.rf_5 [1] ), .B(_00644_ ), .S(_13010_ ), .Z(_00645_ ) );
MUX2_X1 _21192_ ( .A(\wbu.rf_6 [1] ), .B(_00645_ ), .S(_13016_ ), .Z(_00646_ ) );
MUX2_X1 _21193_ ( .A(\wbu.rf_7 [1] ), .B(_00646_ ), .S(_13023_ ), .Z(_00647_ ) );
MUX2_X1 _21194_ ( .A(\wbu.rf_8 [1] ), .B(_00647_ ), .S(_13028_ ), .Z(_00648_ ) );
MUX2_X1 _21195_ ( .A(\wbu.rf_9 [1] ), .B(_00648_ ), .S(_13198_ ), .Z(_00649_ ) );
MUX2_X1 _21196_ ( .A(\wbu.rf_10 [1] ), .B(_00649_ ), .S(_12983_ ), .Z(_00650_ ) );
MUX2_X1 _21197_ ( .A(\wbu.rf_11 [1] ), .B(_00650_ ), .S(_13037_ ), .Z(_00651_ ) );
MUX2_X1 _21198_ ( .A(\wbu.rf_12 [1] ), .B(_00651_ ), .S(_13044_ ), .Z(_00652_ ) );
MUX2_X1 _21199_ ( .A(\wbu.rf_13 [1] ), .B(_00652_ ), .S(_13053_ ), .Z(_00653_ ) );
MUX2_X1 _21200_ ( .A(\wbu.rf_14 [1] ), .B(_00653_ ), .S(_13058_ ), .Z(_00654_ ) );
MUX2_X1 _21201_ ( .A(\wbu.rf_15 [1] ), .B(_00654_ ), .S(_13069_ ), .Z(_00655_ ) );
MUX2_X1 _21202_ ( .A(\wbu.rf_16 [1] ), .B(_00655_ ), .S(_13075_ ), .Z(_00656_ ) );
MUX2_X1 _21203_ ( .A(\wbu.rf_17 [1] ), .B(_00656_ ), .S(_13085_ ), .Z(_00657_ ) );
OAI211_X1 _21204_ ( .A(_13098_ ), .B(_00641_ ), .C1(_00657_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .ZN(_00658_ ) );
NAND4_X1 _21205_ ( .A1(_13105_ ), .A2(_13497_ ), .A3(fanout_net_34 ), .A4(\wbu.rf_19 [1] ), .ZN(_00659_ ) );
NAND3_X1 _21206_ ( .A1(_00658_ ), .A2(_13104_ ), .A3(_00659_ ), .ZN(_00660_ ) );
OAI211_X1 _21207_ ( .A(_00660_ ), .B(_13111_ ), .C1(\wbu.rf_20 [1] ), .C2(_13381_ ), .ZN(_00661_ ) );
NAND4_X1 _21208_ ( .A1(_13119_ ), .A2(_13188_ ), .A3(fanout_net_34 ), .A4(\wbu.rf_21 [1] ), .ZN(_00662_ ) );
NAND3_X1 _21209_ ( .A1(_00661_ ), .A2(_13117_ ), .A3(_00662_ ), .ZN(_00663_ ) );
OAI211_X1 _21210_ ( .A(_00663_ ), .B(_13127_ ), .C1(\wbu.rf_22 [1] ), .C2(_13212_ ), .ZN(_00664_ ) );
NAND4_X1 _21211_ ( .A1(_13186_ ), .A2(fanout_net_34 ), .A3(_13135_ ), .A4(\wbu.rf_23 [1] ), .ZN(_00665_ ) );
NAND3_X1 _21212_ ( .A1(_00664_ ), .A2(_13132_ ), .A3(_00665_ ), .ZN(_00666_ ) );
OAI211_X1 _21213_ ( .A(_00666_ ), .B(_13460_ ), .C1(\wbu.rf_24 [1] ), .C2(_13414_ ), .ZN(_00667_ ) );
NAND4_X1 _21214_ ( .A1(_13312_ ), .A2(_13378_ ), .A3(fanout_net_34 ), .A4(\wbu.rf_25 [1] ), .ZN(_00668_ ) );
NAND3_X1 _21215_ ( .A1(_00667_ ), .A2(_13144_ ), .A3(_00668_ ), .ZN(_00669_ ) );
OAI211_X1 _21216_ ( .A(_00669_ ), .B(_13218_ ), .C1(\wbu.rf_26 [1] ), .C2(_13260_ ), .ZN(_00670_ ) );
NAND4_X1 _21217_ ( .A1(_13158_ ), .A2(fanout_net_34 ), .A3(_13160_ ), .A4(\wbu.rf_27 [1] ), .ZN(_00671_ ) );
NAND3_X1 _21218_ ( .A1(_00670_ ), .A2(_13166_ ), .A3(_00671_ ), .ZN(_00672_ ) );
OAI211_X1 _21219_ ( .A(_00672_ ), .B(_13512_ ), .C1(\wbu.rf_28 [1] ), .C2(_13365_ ), .ZN(_00673_ ) );
NAND4_X1 _21220_ ( .A1(_13326_ ), .A2(fanout_net_34 ), .A3(_13176_ ), .A4(\wbu.rf_29 [1] ), .ZN(_00674_ ) );
AOI21_X1 _21221_ ( .A(_12975_ ), .B1(_00673_ ), .B2(_00674_ ), .ZN(_00675_ ) );
AND4_X1 _21222_ ( .A1(fanout_net_34 ), .A2(_13174_ ), .A3(\wbu.rf_30 [1] ), .A4(_13376_ ), .ZN(_00676_ ) );
OAI21_X1 _21223_ ( .A(_13369_ ), .B1(_00675_ ), .B2(_00676_ ), .ZN(_00677_ ) );
AOI22_X1 _21224_ ( .A1(_12969_ ), .A2(\wbu.rf_31 [1] ), .B1(_13180_ ), .B2(_13182_ ), .ZN(_00678_ ) );
AOI221_X4 _21225_ ( .A(fanout_net_25 ), .B1(_00640_ ), .B2(_12965_ ), .C1(_00677_ ), .C2(_00678_ ), .ZN(_00370_ ) );
NAND4_X1 _21226_ ( .A1(_13272_ ), .A2(\wbu.rf_30 [0] ), .A3(_13273_ ), .A4(fanout_net_34 ), .ZN(_00679_ ) );
AND4_X1 _21227_ ( .A1(\wbu.rf_29 [0] ), .A2(_13326_ ), .A3(fanout_net_34 ), .A4(_13376_ ), .ZN(_00680_ ) );
NAND4_X1 _21228_ ( .A1(_13170_ ), .A2(_13229_ ), .A3(\wbu.rf_28 [0] ), .A4(fanout_net_35 ), .ZN(_00681_ ) );
NAND4_X1 _21229_ ( .A1(_13174_ ), .A2(_13158_ ), .A3(\wbu.rf_26 [0] ), .A4(fanout_net_35 ), .ZN(_00682_ ) );
AND4_X1 _21230_ ( .A1(\wbu.rf_25 [0] ), .A2(_13312_ ), .A3(_13378_ ), .A4(fanout_net_35 ), .ZN(_00683_ ) );
NAND4_X1 _21231_ ( .A1(_13149_ ), .A2(\wbu.rf_24 [0] ), .A3(fanout_net_35 ), .A4(_13229_ ), .ZN(_00684_ ) );
AND4_X1 _21232_ ( .A1(\wbu.rf_22 [0] ), .A2(_13174_ ), .A3(_13122_ ), .A4(fanout_net_35 ), .ZN(_00685_ ) );
NAND4_X1 _21233_ ( .A1(_13120_ ), .A2(_13122_ ), .A3(\wbu.rf_21 [0] ), .A4(fanout_net_35 ), .ZN(_00686_ ) );
AND4_X1 _21234_ ( .A1(\wbu.rf_20 [0] ), .A2(_13121_ ), .A3(fanout_net_35 ), .A4(_13228_ ), .ZN(_00687_ ) );
NAND4_X1 _21235_ ( .A1(_13106_ ), .A2(_08575_ ), .A3(\wbu.rf_19 [0] ), .A4(fanout_net_35 ), .ZN(_00688_ ) );
AND4_X1 _21236_ ( .A1(\wbu.rf_18 [0] ), .A2(_13173_ ), .A3(fanout_net_35 ), .A4(_08574_ ), .ZN(_00689_ ) );
INV_X1 _21237_ ( .A(\wbu.rf_17 [0] ), .ZN(_00690_ ) );
AND4_X1 _21238_ ( .A1(_00690_ ), .A2(_13062_ ), .A3(fanout_net_35 ), .A4(_13350_ ), .ZN(_00691_ ) );
AND4_X1 _21239_ ( .A1(\wbu.rf_16 [0] ), .A2(_13350_ ), .A3(_13228_ ), .A4(fanout_net_35 ), .ZN(_00692_ ) );
NAND4_X1 _21240_ ( .A1(_13077_ ), .A2(_13079_ ), .A3(\wbu.rf_15 [0] ), .A4(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .ZN(_00693_ ) );
AND4_X1 _21241_ ( .A1(\wbu.rf_13 [0] ), .A2(_13061_ ), .A3(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A4(_13063_ ), .ZN(_00694_ ) );
NAND4_X1 _21242_ ( .A1(_13064_ ), .A2(_13228_ ), .A3(\wbu.rf_12 [0] ), .A4(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .ZN(_00695_ ) );
INV_X1 _21243_ ( .A(\wbu.rf_11 [0] ), .ZN(_00696_ ) );
AND4_X1 _21244_ ( .A1(\wbu.rf_10 [0] ), .A2(_12977_ ), .A3(_12986_ ), .A4(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .ZN(_00697_ ) );
MUX2_X1 _21245_ ( .A(\wbu._GEN_71 [0] ), .B(\wbu.rf_2 [0] ), .S(_12992_ ), .Z(_00698_ ) );
MUX2_X1 _21246_ ( .A(\wbu.rf_3 [0] ), .B(_00698_ ), .S(_12998_ ), .Z(_00699_ ) );
MUX2_X1 _21247_ ( .A(\wbu.rf_4 [0] ), .B(_00699_ ), .S(_13004_ ), .Z(_00700_ ) );
MUX2_X1 _21248_ ( .A(\wbu.rf_5 [0] ), .B(_00700_ ), .S(_13012_ ), .Z(_00701_ ) );
MUX2_X1 _21249_ ( .A(\wbu.rf_6 [0] ), .B(_00701_ ), .S(_13017_ ), .Z(_00702_ ) );
MUX2_X1 _21250_ ( .A(\wbu.rf_7 [0] ), .B(_00702_ ), .S(_13024_ ), .Z(_00703_ ) );
MUX2_X1 _21251_ ( .A(\wbu.rf_8 [0] ), .B(_00703_ ), .S(_13030_ ), .Z(_00704_ ) );
MUX2_X1 _21252_ ( .A(\wbu.rf_9 [0] ), .B(_00704_ ), .S(_13383_ ), .Z(_00705_ ) );
AOI21_X1 _21253_ ( .A(_00697_ ), .B1(_00705_ ), .B2(_12984_ ), .ZN(_00706_ ) );
MUX2_X1 _21254_ ( .A(_00696_ ), .B(_00706_ ), .S(_13038_ ), .Z(_00707_ ) );
OAI21_X1 _21255_ ( .A(_00695_ ), .B1(_00707_ ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_00708_ ) );
AOI21_X1 _21256_ ( .A(_00694_ ), .B1(_00708_ ), .B2(_13054_ ), .ZN(_00709_ ) );
NAND2_X1 _21257_ ( .A1(_00709_ ), .A2(_13071_ ), .ZN(_00710_ ) );
OAI21_X1 _21258_ ( .A(_00710_ ), .B1(\wbu.rf_14 [0] ), .B2(_13071_ ), .ZN(_00711_ ) );
OAI21_X1 _21259_ ( .A(_00693_ ), .B1(_00711_ ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .ZN(_00712_ ) );
AOI21_X1 _21260_ ( .A(_00692_ ), .B1(_00712_ ), .B2(_13087_ ), .ZN(_00713_ ) );
AOI21_X1 _21261_ ( .A(_00691_ ), .B1(_00713_ ), .B2(_13086_ ), .ZN(_00714_ ) );
AOI21_X1 _21262_ ( .A(_00689_ ), .B1(_00714_ ), .B2(_13099_ ), .ZN(_00715_ ) );
OAI21_X1 _21263_ ( .A(_00688_ ), .B1(_00715_ ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .ZN(_00716_ ) );
AOI21_X1 _21264_ ( .A(_00687_ ), .B1(_00716_ ), .B2(_13113_ ), .ZN(_00717_ ) );
OAI21_X1 _21265_ ( .A(_00686_ ), .B1(_00717_ ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_00718_ ) );
AOI21_X1 _21266_ ( .A(_00685_ ), .B1(_00718_ ), .B2(_13128_ ), .ZN(_00719_ ) );
NAND2_X1 _21267_ ( .A1(_00719_ ), .A2(_13231_ ), .ZN(_00720_ ) );
OAI21_X1 _21268_ ( .A(_00720_ ), .B1(\wbu.rf_23 [0] ), .B2(_13231_ ), .ZN(_00721_ ) );
OAI21_X1 _21269_ ( .A(_00684_ ), .B1(_00721_ ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_1_Y ), .ZN(_00722_ ) );
AOI21_X1 _21270_ ( .A(_00683_ ), .B1(_00722_ ), .B2(_13140_ ), .ZN(_00723_ ) );
OAI211_X1 _21271_ ( .A(_13153_ ), .B(_00682_ ), .C1(_00723_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_00724_ ) );
OAI21_X1 _21272_ ( .A(_00724_ ), .B1(\wbu.rf_27 [0] ), .B2(_13153_ ), .ZN(_00725_ ) );
OAI21_X1 _21273_ ( .A(_00681_ ), .B1(_00725_ ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_00726_ ) );
AOI21_X1 _21274_ ( .A(_00680_ ), .B1(_00726_ ), .B2(_13269_ ), .ZN(_00727_ ) );
OAI211_X1 _21275_ ( .A(_13374_ ), .B(_00679_ ), .C1(_00727_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_00728_ ) );
OAI211_X1 _21276_ ( .A(_00728_ ), .B(_13276_ ), .C1(\wbu.rf_31 [0] ), .C2(_13271_ ), .ZN(_00729_ ) );
NAND3_X1 _21277_ ( .A1(_13181_ ), .A2(\wbu.io_in_bits_rd_wdata [0] ), .A3(_13183_ ), .ZN(_00730_ ) );
AOI21_X1 _21278_ ( .A(fanout_net_25 ), .B1(_00729_ ), .B2(_00730_ ), .ZN(_00371_ ) );
AND3_X1 _21279_ ( .A1(_13474_ ), .A2(fanout_net_35 ), .A3(\wbu.rf_31 [27] ), .ZN(_00731_ ) );
AND3_X1 _21280_ ( .A1(_12994_ ), .A2(fanout_net_35 ), .A3(\wbu.rf_19 [27] ), .ZN(_00732_ ) );
NAND4_X1 _21281_ ( .A1(_13174_ ), .A2(fanout_net_35 ), .A3(\wbu.rf_18 [27] ), .A4(_13497_ ), .ZN(_00733_ ) );
AND4_X1 _21282_ ( .A1(fanout_net_35 ), .A2(_13062_ ), .A3(\wbu.rf_17 [27] ), .A4(_13350_ ), .ZN(_00734_ ) );
MUX2_X1 _21283_ ( .A(\wbu._GEN_71 [27] ), .B(\wbu.rf_2 [27] ), .S(_12992_ ), .Z(_00735_ ) );
MUX2_X1 _21284_ ( .A(\wbu.rf_3 [27] ), .B(_00735_ ), .S(_12997_ ), .Z(_00736_ ) );
MUX2_X1 _21285_ ( .A(\wbu.rf_4 [27] ), .B(_00736_ ), .S(_13003_ ), .Z(_00737_ ) );
MUX2_X1 _21286_ ( .A(\wbu.rf_5 [27] ), .B(_00737_ ), .S(_13011_ ), .Z(_00738_ ) );
MUX2_X1 _21287_ ( .A(\wbu.rf_6 [27] ), .B(_00738_ ), .S(_13017_ ), .Z(_00739_ ) );
MUX2_X1 _21288_ ( .A(\wbu.rf_7 [27] ), .B(_00739_ ), .S(_13023_ ), .Z(_00740_ ) );
MUX2_X1 _21289_ ( .A(\wbu.rf_8 [27] ), .B(_00740_ ), .S(_13029_ ), .Z(_00741_ ) );
MUX2_X1 _21290_ ( .A(\wbu.rf_9 [27] ), .B(_00741_ ), .S(_13198_ ), .Z(_00742_ ) );
MUX2_X1 _21291_ ( .A(\wbu.rf_10 [27] ), .B(_00742_ ), .S(_12983_ ), .Z(_00743_ ) );
MUX2_X1 _21292_ ( .A(\wbu.rf_11 [27] ), .B(_00743_ ), .S(_13037_ ), .Z(_00744_ ) );
MUX2_X1 _21293_ ( .A(\wbu.rf_12 [27] ), .B(_00744_ ), .S(_13044_ ), .Z(_00745_ ) );
MUX2_X1 _21294_ ( .A(\wbu.rf_13 [27] ), .B(_00745_ ), .S(_13053_ ), .Z(_00746_ ) );
MUX2_X1 _21295_ ( .A(\wbu.rf_14 [27] ), .B(_00746_ ), .S(_13059_ ), .Z(_00747_ ) );
MUX2_X1 _21296_ ( .A(\wbu.rf_15 [27] ), .B(_00747_ ), .S(_13069_ ), .Z(_00748_ ) );
MUX2_X1 _21297_ ( .A(\wbu.rf_16 [27] ), .B(_00748_ ), .S(_13075_ ), .Z(_00749_ ) );
AOI21_X1 _21298_ ( .A(_00734_ ), .B1(_00749_ ), .B2(_13086_ ), .ZN(_00750_ ) );
OAI21_X1 _21299_ ( .A(_00733_ ), .B1(_00750_ ), .B2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .ZN(_00751_ ) );
AOI211_X1 _21300_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .B(_00732_ ), .C1(_00751_ ), .C2(_13098_ ), .ZN(_00752_ ) );
NOR2_X1 _21301_ ( .A1(_13104_ ), .A2(\wbu.rf_20 [27] ), .ZN(_00753_ ) );
NOR3_X1 _21302_ ( .A1(_00752_ ), .A2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_1_Y ), .A3(_00753_ ), .ZN(_00754_ ) );
NAND3_X1 _21303_ ( .A1(_13008_ ), .A2(fanout_net_35 ), .A3(\wbu.rf_21 [27] ), .ZN(_00755_ ) );
NAND2_X1 _21304_ ( .A1(_13117_ ), .A2(_00755_ ), .ZN(_00756_ ) );
OAI221_X1 _21305_ ( .A(_13126_ ), .B1(\wbu.rf_22 [27] ), .B2(_13117_ ), .C1(_00754_ ), .C2(_00756_ ), .ZN(_00757_ ) );
NAND4_X1 _21306_ ( .A1(_13186_ ), .A2(fanout_net_35 ), .A3(_13134_ ), .A4(\wbu.rf_23 [27] ), .ZN(_00758_ ) );
NAND3_X1 _21307_ ( .A1(_00757_ ), .A2(_13131_ ), .A3(_00758_ ), .ZN(_00759_ ) );
OAI211_X1 _21308_ ( .A(_00759_ ), .B(_13460_ ), .C1(\wbu.rf_24 [27] ), .C2(_13414_ ), .ZN(_00760_ ) );
NAND4_X1 _21309_ ( .A1(_13146_ ), .A2(_13378_ ), .A3(fanout_net_35 ), .A4(\wbu.rf_25 [27] ), .ZN(_00761_ ) );
NAND3_X1 _21310_ ( .A1(_00760_ ), .A2(_13144_ ), .A3(_00761_ ), .ZN(_00762_ ) );
OAI211_X1 _21311_ ( .A(_00762_ ), .B(_13363_ ), .C1(\wbu.rf_26 [27] ), .C2(_13145_ ), .ZN(_00763_ ) );
NAND4_X1 _21312_ ( .A1(_13158_ ), .A2(fanout_net_35 ), .A3(_13160_ ), .A4(\wbu.rf_27 [27] ), .ZN(_00764_ ) );
NAND3_X1 _21313_ ( .A1(_00763_ ), .A2(_13166_ ), .A3(_00764_ ), .ZN(_00765_ ) );
OAI211_X1 _21314_ ( .A(_00765_ ), .B(_13512_ ), .C1(\wbu.rf_28 [27] ), .C2(_13365_ ), .ZN(_00766_ ) );
NAND4_X1 _21315_ ( .A1(_13326_ ), .A2(fanout_net_35 ), .A3(_13327_ ), .A4(\wbu.rf_29 [27] ), .ZN(_00767_ ) );
NAND2_X1 _21316_ ( .A1(_00766_ ), .A2(_00767_ ), .ZN(_00768_ ) );
MUX2_X1 _21317_ ( .A(\wbu.rf_30 [27] ), .B(_00768_ ), .S(_13267_ ), .Z(_00769_ ) );
AOI211_X1 _21318_ ( .A(_13473_ ), .B(_00731_ ), .C1(_00769_ ), .C2(_13374_ ), .ZN(_00770_ ) );
INV_X1 _21319_ ( .A(\wbu.io_in_bits_rd_wdata [27] ), .ZN(_00771_ ) );
AOI211_X1 _21320_ ( .A(fanout_net_25 ), .B(_00770_ ), .C1(_00771_ ), .C2(_13324_ ), .ZN(_00372_ ) );
AND3_X1 _21321_ ( .A1(_13474_ ), .A2(fanout_net_35 ), .A3(\wbu.rf_31 [26] ), .ZN(_00772_ ) );
NAND4_X1 _21322_ ( .A1(_13173_ ), .A2(fanout_net_35 ), .A3(\wbu.rf_18 [26] ), .A4(_08573_ ), .ZN(_00773_ ) );
AND4_X1 _21323_ ( .A1(fanout_net_35 ), .A2(_13061_ ), .A3(\wbu.rf_17 [26] ), .A4(_08573_ ), .ZN(_00774_ ) );
MUX2_X1 _21324_ ( .A(\wbu._GEN_71 [26] ), .B(\wbu.rf_2 [26] ), .S(_12990_ ), .Z(_00775_ ) );
MUX2_X1 _21325_ ( .A(\wbu.rf_3 [26] ), .B(_00775_ ), .S(_12995_ ), .Z(_00776_ ) );
MUX2_X1 _21326_ ( .A(\wbu.rf_4 [26] ), .B(_00776_ ), .S(_13001_ ), .Z(_00777_ ) );
MUX2_X1 _21327_ ( .A(\wbu.rf_5 [26] ), .B(_00777_ ), .S(_13009_ ), .Z(_00778_ ) );
MUX2_X1 _21328_ ( .A(\wbu.rf_6 [26] ), .B(_00778_ ), .S(_13015_ ), .Z(_00779_ ) );
MUX2_X1 _21329_ ( .A(\wbu.rf_7 [26] ), .B(_00779_ ), .S(_13021_ ), .Z(_00780_ ) );
MUX2_X1 _21330_ ( .A(\wbu.rf_8 [26] ), .B(_00780_ ), .S(_13028_ ), .Z(_00781_ ) );
MUX2_X1 _21331_ ( .A(\wbu.rf_9 [26] ), .B(_00781_ ), .S(_13197_ ), .Z(_00782_ ) );
MUX2_X1 _21332_ ( .A(\wbu.rf_10 [26] ), .B(_00782_ ), .S(_12982_ ), .Z(_00783_ ) );
MUX2_X1 _21333_ ( .A(\wbu.rf_11 [26] ), .B(_00783_ ), .S(_13036_ ), .Z(_00784_ ) );
MUX2_X1 _21334_ ( .A(\wbu.rf_12 [26] ), .B(_00784_ ), .S(_13043_ ), .Z(_00785_ ) );
MUX2_X1 _21335_ ( .A(\wbu.rf_13 [26] ), .B(_00785_ ), .S(_13052_ ), .Z(_00786_ ) );
MUX2_X1 _21336_ ( .A(\wbu.rf_14 [26] ), .B(_00786_ ), .S(_13058_ ), .Z(_00787_ ) );
MUX2_X1 _21337_ ( .A(\wbu.rf_15 [26] ), .B(_00787_ ), .S(_13068_ ), .Z(_00788_ ) );
MUX2_X1 _21338_ ( .A(\wbu.rf_16 [26] ), .B(_00788_ ), .S(_13074_ ), .Z(_00789_ ) );
AOI21_X1 _21339_ ( .A(_00774_ ), .B1(_00789_ ), .B2(_13084_ ), .ZN(_00790_ ) );
OAI211_X1 _21340_ ( .A(_13096_ ), .B(_00773_ ), .C1(_00790_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .ZN(_00791_ ) );
OAI211_X1 _21341_ ( .A(_00791_ ), .B(_13102_ ), .C1(\wbu.rf_19 [26] ), .C2(_13096_ ), .ZN(_00792_ ) );
NAND4_X1 _21342_ ( .A1(_13121_ ), .A2(fanout_net_35 ), .A3(\wbu.rf_20 [26] ), .A4(_13228_ ), .ZN(_00793_ ) );
AOI21_X1 _21343_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_1_Y ), .B1(_00792_ ), .B2(_00793_ ), .ZN(_00794_ ) );
NAND3_X1 _21344_ ( .A1(_13008_ ), .A2(fanout_net_35 ), .A3(\wbu.rf_21 [26] ), .ZN(_00795_ ) );
NAND2_X1 _21345_ ( .A1(_13116_ ), .A2(_00795_ ), .ZN(_00796_ ) );
OAI221_X1 _21346_ ( .A(_13125_ ), .B1(\wbu.rf_22 [26] ), .B2(_13116_ ), .C1(_00794_ ), .C2(_00796_ ), .ZN(_00797_ ) );
NAND4_X1 _21347_ ( .A1(_13121_ ), .A2(fanout_net_35 ), .A3(_13105_ ), .A4(\wbu.rf_23 [26] ), .ZN(_00798_ ) );
NAND2_X1 _21348_ ( .A1(_00797_ ), .A2(_00798_ ), .ZN(_00799_ ) );
MUX2_X1 _21349_ ( .A(\wbu.rf_24 [26] ), .B(_00799_ ), .S(_13130_ ), .Z(_00800_ ) );
MUX2_X1 _21350_ ( .A(\wbu.rf_25 [26] ), .B(_00800_ ), .S(_13139_ ), .Z(_00801_ ) );
MUX2_X1 _21351_ ( .A(\wbu.rf_26 [26] ), .B(_00801_ ), .S(_13143_ ), .Z(_00802_ ) );
MUX2_X1 _21352_ ( .A(\wbu.rf_27 [26] ), .B(_00802_ ), .S(_13152_ ), .Z(_00803_ ) );
MUX2_X1 _21353_ ( .A(\wbu.rf_28 [26] ), .B(_00803_ ), .S(_13156_ ), .Z(_00804_ ) );
MUX2_X1 _21354_ ( .A(\wbu.rf_29 [26] ), .B(_00804_ ), .S(_13164_ ), .Z(_00805_ ) );
MUX2_X1 _21355_ ( .A(\wbu.rf_30 [26] ), .B(_00805_ ), .S(_13267_ ), .Z(_00806_ ) );
AOI211_X1 _21356_ ( .A(_13473_ ), .B(_00772_ ), .C1(_00806_ ), .C2(_13374_ ), .ZN(_00807_ ) );
INV_X1 _21357_ ( .A(\wbu.io_in_bits_rd_wdata [26] ), .ZN(_00808_ ) );
AOI211_X1 _21358_ ( .A(fanout_net_25 ), .B(_00807_ ), .C1(_00808_ ), .C2(_13324_ ), .ZN(_00373_ ) );
AND3_X1 _21359_ ( .A1(_13474_ ), .A2(fanout_net_35 ), .A3(\wbu.rf_31 [25] ), .ZN(_00809_ ) );
NAND4_X1 _21360_ ( .A1(_08572_ ), .A2(_12960_ ), .A3(fanout_net_35 ), .A4(\wbu.rf_16 [25] ), .ZN(_00810_ ) );
AND4_X1 _21361_ ( .A1(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A2(_12966_ ), .A3(_13063_ ), .A4(\wbu.rf_15 [25] ), .ZN(_00811_ ) );
MUX2_X1 _21362_ ( .A(\wbu._GEN_71 [25] ), .B(\wbu.rf_2 [25] ), .S(_12990_ ), .Z(_00812_ ) );
MUX2_X1 _21363_ ( .A(\wbu.rf_3 [25] ), .B(_00812_ ), .S(_12996_ ), .Z(_00813_ ) );
MUX2_X1 _21364_ ( .A(\wbu.rf_4 [25] ), .B(_00813_ ), .S(_13002_ ), .Z(_00814_ ) );
MUX2_X1 _21365_ ( .A(\wbu.rf_5 [25] ), .B(_00814_ ), .S(_13010_ ), .Z(_00815_ ) );
MUX2_X1 _21366_ ( .A(\wbu.rf_6 [25] ), .B(_00815_ ), .S(_13015_ ), .Z(_00816_ ) );
MUX2_X1 _21367_ ( .A(\wbu.rf_7 [25] ), .B(_00816_ ), .S(_13022_ ), .Z(_00817_ ) );
MUX2_X1 _21368_ ( .A(\wbu.rf_8 [25] ), .B(_00817_ ), .S(_13028_ ), .Z(_00818_ ) );
MUX2_X1 _21369_ ( .A(\wbu.rf_9 [25] ), .B(_00818_ ), .S(_13197_ ), .Z(_00819_ ) );
MUX2_X1 _21370_ ( .A(\wbu.rf_10 [25] ), .B(_00819_ ), .S(_12982_ ), .Z(_00820_ ) );
MUX2_X1 _21371_ ( .A(\wbu.rf_11 [25] ), .B(_00820_ ), .S(_13036_ ), .Z(_00821_ ) );
MUX2_X1 _21372_ ( .A(\wbu.rf_12 [25] ), .B(_00821_ ), .S(_13043_ ), .Z(_00822_ ) );
MUX2_X1 _21373_ ( .A(\wbu.rf_13 [25] ), .B(_00822_ ), .S(_13052_ ), .Z(_00823_ ) );
MUX2_X1 _21374_ ( .A(\wbu.rf_14 [25] ), .B(_00823_ ), .S(_13058_ ), .Z(_00824_ ) );
AOI21_X1 _21375_ ( .A(_00811_ ), .B1(_00824_ ), .B2(_13068_ ), .ZN(_00825_ ) );
OAI211_X1 _21376_ ( .A(_13084_ ), .B(_00810_ ), .C1(_00825_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__B_Y ), .ZN(_00826_ ) );
OAI211_X1 _21377_ ( .A(_00826_ ), .B(_13089_ ), .C1(\wbu.rf_17 [25] ), .C2(_13084_ ), .ZN(_00827_ ) );
NAND4_X1 _21378_ ( .A1(_13173_ ), .A2(fanout_net_35 ), .A3(\wbu.rf_18 [25] ), .A4(_08573_ ), .ZN(_00828_ ) );
AOI21_X1 _21379_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .B1(_00827_ ), .B2(_00828_ ), .ZN(_00829_ ) );
NAND3_X1 _21380_ ( .A1(_12994_ ), .A2(fanout_net_35 ), .A3(\wbu.rf_19 [25] ), .ZN(_00830_ ) );
NAND2_X1 _21381_ ( .A1(_13101_ ), .A2(_00830_ ), .ZN(_00831_ ) );
OAI221_X1 _21382_ ( .A(_13110_ ), .B1(\wbu.rf_20 [25] ), .B2(_13102_ ), .C1(_00829_ ), .C2(_00831_ ), .ZN(_00832_ ) );
NAND4_X1 _21383_ ( .A1(_13061_ ), .A2(_13007_ ), .A3(fanout_net_36 ), .A4(\wbu.rf_21 [25] ), .ZN(_00833_ ) );
NAND2_X1 _21384_ ( .A1(_00832_ ), .A2(_00833_ ), .ZN(_00834_ ) );
MUX2_X1 _21385_ ( .A(\wbu.rf_22 [25] ), .B(_00834_ ), .S(_13115_ ), .Z(_00835_ ) );
MUX2_X1 _21386_ ( .A(\wbu.rf_23 [25] ), .B(_00835_ ), .S(_13125_ ), .Z(_00836_ ) );
MUX2_X1 _21387_ ( .A(\wbu.rf_24 [25] ), .B(_00836_ ), .S(_13130_ ), .Z(_00837_ ) );
MUX2_X1 _21388_ ( .A(\wbu.rf_25 [25] ), .B(_00837_ ), .S(_13138_ ), .Z(_00838_ ) );
MUX2_X1 _21389_ ( .A(\wbu.rf_26 [25] ), .B(_00838_ ), .S(_13143_ ), .Z(_00839_ ) );
MUX2_X1 _21390_ ( .A(\wbu.rf_27 [25] ), .B(_00839_ ), .S(_13152_ ), .Z(_00840_ ) );
MUX2_X1 _21391_ ( .A(\wbu.rf_28 [25] ), .B(_00840_ ), .S(_13156_ ), .Z(_00841_ ) );
MUX2_X1 _21392_ ( .A(\wbu.rf_29 [25] ), .B(_00841_ ), .S(_13164_ ), .Z(_00842_ ) );
MUX2_X1 _21393_ ( .A(\wbu.rf_30 [25] ), .B(_00842_ ), .S(_13267_ ), .Z(_00843_ ) );
AOI211_X1 _21394_ ( .A(_13473_ ), .B(_00809_ ), .C1(_00843_ ), .C2(_13374_ ), .ZN(_00844_ ) );
INV_X1 _21395_ ( .A(\wbu.io_in_bits_rd_wdata [25] ), .ZN(_00845_ ) );
AOI211_X1 _21396_ ( .A(fanout_net_25 ), .B(_00844_ ), .C1(_00845_ ), .C2(_13324_ ), .ZN(_00374_ ) );
AND3_X1 _21397_ ( .A1(_13474_ ), .A2(fanout_net_36 ), .A3(\wbu.rf_31 [24] ), .ZN(_00846_ ) );
OAI21_X1 _21398_ ( .A(_13363_ ), .B1(_13145_ ), .B2(\wbu.rf_26 [24] ), .ZN(_00847_ ) );
NAND4_X1 _21399_ ( .A1(_13134_ ), .A2(_08575_ ), .A3(fanout_net_36 ), .A4(\wbu.rf_19 [24] ), .ZN(_00848_ ) );
AND4_X1 _21400_ ( .A1(fanout_net_36 ), .A2(_13173_ ), .A3(\wbu.rf_18 [24] ), .A4(_08574_ ), .ZN(_00849_ ) );
MUX2_X1 _21401_ ( .A(\wbu._GEN_71 [24] ), .B(\wbu.rf_2 [24] ), .S(_12992_ ), .Z(_00850_ ) );
MUX2_X1 _21402_ ( .A(\wbu.rf_3 [24] ), .B(_00850_ ), .S(_12997_ ), .Z(_00851_ ) );
MUX2_X1 _21403_ ( .A(\wbu.rf_4 [24] ), .B(_00851_ ), .S(_13003_ ), .Z(_00852_ ) );
MUX2_X1 _21404_ ( .A(\wbu.rf_5 [24] ), .B(_00852_ ), .S(_13011_ ), .Z(_00853_ ) );
MUX2_X1 _21405_ ( .A(\wbu.rf_6 [24] ), .B(_00853_ ), .S(_13017_ ), .Z(_00854_ ) );
MUX2_X1 _21406_ ( .A(\wbu.rf_7 [24] ), .B(_00854_ ), .S(_13023_ ), .Z(_00855_ ) );
MUX2_X1 _21407_ ( .A(\wbu.rf_8 [24] ), .B(_00855_ ), .S(_13029_ ), .Z(_00856_ ) );
MUX2_X1 _21408_ ( .A(\wbu.rf_9 [24] ), .B(_00856_ ), .S(_13198_ ), .Z(_00857_ ) );
MUX2_X1 _21409_ ( .A(\wbu.rf_10 [24] ), .B(_00857_ ), .S(_12983_ ), .Z(_00858_ ) );
MUX2_X1 _21410_ ( .A(\wbu.rf_11 [24] ), .B(_00858_ ), .S(_13037_ ), .Z(_00859_ ) );
MUX2_X1 _21411_ ( .A(\wbu.rf_12 [24] ), .B(_00859_ ), .S(_13044_ ), .Z(_00860_ ) );
MUX2_X1 _21412_ ( .A(\wbu.rf_13 [24] ), .B(_00860_ ), .S(_13053_ ), .Z(_00861_ ) );
MUX2_X1 _21413_ ( .A(\wbu.rf_14 [24] ), .B(_00861_ ), .S(_13059_ ), .Z(_00862_ ) );
MUX2_X1 _21414_ ( .A(\wbu.rf_15 [24] ), .B(_00862_ ), .S(_13069_ ), .Z(_00863_ ) );
MUX2_X1 _21415_ ( .A(\wbu.rf_16 [24] ), .B(_00863_ ), .S(_13075_ ), .Z(_00864_ ) );
MUX2_X1 _21416_ ( .A(\wbu.rf_17 [24] ), .B(_00864_ ), .S(_13086_ ), .Z(_00865_ ) );
AOI21_X1 _21417_ ( .A(_00849_ ), .B1(_00865_ ), .B2(_13099_ ), .ZN(_00866_ ) );
OAI211_X1 _21418_ ( .A(_13113_ ), .B(_00848_ ), .C1(_00866_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .ZN(_00867_ ) );
OAI211_X1 _21419_ ( .A(_00867_ ), .B(_13112_ ), .C1(\wbu.rf_20 [24] ), .C2(_13113_ ), .ZN(_00868_ ) );
NAND4_X1 _21420_ ( .A1(_13146_ ), .A2(_13186_ ), .A3(fanout_net_36 ), .A4(\wbu.rf_21 [24] ), .ZN(_00869_ ) );
NAND3_X1 _21421_ ( .A1(_00868_ ), .A2(_13128_ ), .A3(_00869_ ), .ZN(_00870_ ) );
OAI211_X1 _21422_ ( .A(_00870_ ), .B(_13231_ ), .C1(\wbu.rf_22 [24] ), .C2(_13128_ ), .ZN(_00871_ ) );
NAND4_X1 _21423_ ( .A1(_13133_ ), .A2(fanout_net_36 ), .A3(_13160_ ), .A4(\wbu.rf_23 [24] ), .ZN(_00872_ ) );
AOI21_X1 _21424_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_1_Y ), .B1(_00871_ ), .B2(_00872_ ), .ZN(_00873_ ) );
AND4_X1 _21425_ ( .A1(fanout_net_36 ), .A2(_13378_ ), .A3(\wbu.rf_24 [24] ), .A4(_13229_ ), .ZN(_00874_ ) );
OAI21_X1 _21426_ ( .A(_13140_ ), .B1(_00873_ ), .B2(_00874_ ), .ZN(_00875_ ) );
AOI22_X1 _21427_ ( .A1(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .A2(\wbu.rf_25 [24] ), .B1(fanout_net_36 ), .B2(_12980_ ), .ZN(_00876_ ) );
AOI21_X1 _21428_ ( .A(_00847_ ), .B1(_00875_ ), .B2(_00876_ ), .ZN(_00877_ ) );
NAND3_X1 _21429_ ( .A1(_13034_ ), .A2(fanout_net_36 ), .A3(\wbu.rf_27 [24] ), .ZN(_00878_ ) );
NAND2_X1 _21430_ ( .A1(_13156_ ), .A2(_00878_ ), .ZN(_00879_ ) );
OAI221_X1 _21431_ ( .A(_13164_ ), .B1(\wbu.rf_28 [24] ), .B2(_13166_ ), .C1(_00877_ ), .C2(_00879_ ), .ZN(_00880_ ) );
NAND4_X1 _21432_ ( .A1(_13326_ ), .A2(fanout_net_36 ), .A3(_13327_ ), .A4(\wbu.rf_29 [24] ), .ZN(_00881_ ) );
NAND2_X1 _21433_ ( .A1(_00880_ ), .A2(_00881_ ), .ZN(_00882_ ) );
MUX2_X1 _21434_ ( .A(\wbu.rf_30 [24] ), .B(_00882_ ), .S(_13267_ ), .Z(_00883_ ) );
AOI211_X1 _21435_ ( .A(_13473_ ), .B(_00846_ ), .C1(_00883_ ), .C2(_13374_ ), .ZN(_00884_ ) );
INV_X1 _21436_ ( .A(\wbu.io_in_bits_rd_wdata [24] ), .ZN(_00885_ ) );
AOI211_X1 _21437_ ( .A(fanout_net_25 ), .B(_00884_ ), .C1(_00885_ ), .C2(_13324_ ), .ZN(_00375_ ) );
AND3_X1 _21438_ ( .A1(_12980_ ), .A2(fanout_net_36 ), .A3(\wbu.rf_26 [23] ), .ZN(_00886_ ) );
NAND4_X1 _21439_ ( .A1(_13188_ ), .A2(fanout_net_36 ), .A3(\wbu.rf_20 [23] ), .A4(_13228_ ), .ZN(_00887_ ) );
AND4_X1 _21440_ ( .A1(fanout_net_36 ), .A2(_13105_ ), .A3(\wbu.rf_19 [23] ), .A4(_13497_ ), .ZN(_00888_ ) );
MUX2_X1 _21441_ ( .A(\wbu._GEN_71 [23] ), .B(\wbu.rf_2 [23] ), .S(_12991_ ), .Z(_00889_ ) );
MUX2_X1 _21442_ ( .A(\wbu.rf_3 [23] ), .B(_00889_ ), .S(_12996_ ), .Z(_00890_ ) );
MUX2_X1 _21443_ ( .A(\wbu.rf_4 [23] ), .B(_00890_ ), .S(_13002_ ), .Z(_00891_ ) );
MUX2_X1 _21444_ ( .A(\wbu.rf_5 [23] ), .B(_00891_ ), .S(_13010_ ), .Z(_00892_ ) );
MUX2_X1 _21445_ ( .A(\wbu.rf_6 [23] ), .B(_00892_ ), .S(_13016_ ), .Z(_00893_ ) );
MUX2_X1 _21446_ ( .A(\wbu.rf_7 [23] ), .B(_00893_ ), .S(_13022_ ), .Z(_00894_ ) );
MUX2_X1 _21447_ ( .A(\wbu.rf_8 [23] ), .B(_00894_ ), .S(_13028_ ), .Z(_00895_ ) );
MUX2_X1 _21448_ ( .A(\wbu.rf_9 [23] ), .B(_00895_ ), .S(_13198_ ), .Z(_00896_ ) );
MUX2_X1 _21449_ ( .A(\wbu.rf_10 [23] ), .B(_00896_ ), .S(_12983_ ), .Z(_00897_ ) );
MUX2_X1 _21450_ ( .A(\wbu.rf_11 [23] ), .B(_00897_ ), .S(_13037_ ), .Z(_00898_ ) );
MUX2_X1 _21451_ ( .A(\wbu.rf_12 [23] ), .B(_00898_ ), .S(_13044_ ), .Z(_00899_ ) );
MUX2_X1 _21452_ ( .A(\wbu.rf_13 [23] ), .B(_00899_ ), .S(_13053_ ), .Z(_00900_ ) );
MUX2_X1 _21453_ ( .A(\wbu.rf_14 [23] ), .B(_00900_ ), .S(_13058_ ), .Z(_00901_ ) );
MUX2_X1 _21454_ ( .A(\wbu.rf_15 [23] ), .B(_00901_ ), .S(_13069_ ), .Z(_00902_ ) );
MUX2_X1 _21455_ ( .A(\wbu.rf_16 [23] ), .B(_00902_ ), .S(_13074_ ), .Z(_00903_ ) );
MUX2_X1 _21456_ ( .A(\wbu.rf_17 [23] ), .B(_00903_ ), .S(_13085_ ), .Z(_00904_ ) );
MUX2_X1 _21457_ ( .A(\wbu.rf_18 [23] ), .B(_00904_ ), .S(_13450_ ), .Z(_00905_ ) );
AOI21_X1 _21458_ ( .A(_00888_ ), .B1(_00905_ ), .B2(_13098_ ), .ZN(_00906_ ) );
OAI211_X1 _21459_ ( .A(_13112_ ), .B(_00887_ ), .C1(_00906_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .ZN(_00907_ ) );
OAI211_X1 _21460_ ( .A(_00907_ ), .B(_13128_ ), .C1(\wbu.rf_21 [23] ), .C2(_13112_ ), .ZN(_00908_ ) );
NAND4_X1 _21461_ ( .A1(_13174_ ), .A2(_13186_ ), .A3(fanout_net_36 ), .A4(\wbu.rf_22 [23] ), .ZN(_00909_ ) );
NAND3_X1 _21462_ ( .A1(_00908_ ), .A2(_13231_ ), .A3(_00909_ ), .ZN(_00910_ ) );
OAI211_X1 _21463_ ( .A(_00910_ ), .B(_13141_ ), .C1(\wbu.rf_23 [23] ), .C2(_13231_ ), .ZN(_00911_ ) );
NAND4_X1 _21464_ ( .A1(_13149_ ), .A2(fanout_net_36 ), .A3(\wbu.rf_24 [23] ), .A4(_13229_ ), .ZN(_00912_ ) );
NAND2_X1 _21465_ ( .A1(_00911_ ), .A2(_00912_ ), .ZN(_00913_ ) );
MUX2_X1 _21466_ ( .A(\wbu.rf_25 [23] ), .B(_00913_ ), .S(_13140_ ), .Z(_00914_ ) );
AOI211_X1 _21467_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .B(_00886_ ), .C1(_00914_ ), .C2(_13154_ ), .ZN(_00915_ ) );
NOR2_X1 _21468_ ( .A1(_13153_ ), .A2(\wbu.rf_27 [23] ), .ZN(_00916_ ) );
NOR3_X1 _21469_ ( .A1(_00915_ ), .A2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .A3(_00916_ ), .ZN(_00917_ ) );
NAND3_X1 _21470_ ( .A1(_13041_ ), .A2(fanout_net_36 ), .A3(\wbu.rf_28 [23] ), .ZN(_00918_ ) );
NAND2_X1 _21471_ ( .A1(_13165_ ), .A2(_00918_ ), .ZN(_00919_ ) );
OAI221_X1 _21472_ ( .A(_13268_ ), .B1(\wbu.rf_29 [23] ), .B2(_13269_ ), .C1(_00917_ ), .C2(_00919_ ), .ZN(_00920_ ) );
NAND4_X1 _21473_ ( .A1(_13272_ ), .A2(fanout_net_36 ), .A3(_13273_ ), .A4(\wbu.rf_30 [23] ), .ZN(_00921_ ) );
NAND3_X1 _21474_ ( .A1(_00920_ ), .A2(_13271_ ), .A3(_00921_ ), .ZN(_00922_ ) );
OAI211_X1 _21475_ ( .A(_00922_ ), .B(_13276_ ), .C1(\wbu.rf_31 [23] ), .C2(_13271_ ), .ZN(_00923_ ) );
NAND3_X1 _21476_ ( .A1(_13181_ ), .A2(\wbu.io_in_bits_rd_wdata [23] ), .A3(_13183_ ), .ZN(_00924_ ) );
AOI21_X1 _21477_ ( .A(fanout_net_25 ), .B1(_00923_ ), .B2(_00924_ ), .ZN(_00376_ ) );
NAND4_X1 _21478_ ( .A1(_13272_ ), .A2(fanout_net_36 ), .A3(_13273_ ), .A4(\wbu.rf_30 [22] ), .ZN(_00925_ ) );
AND4_X1 _21479_ ( .A1(fanout_net_36 ), .A2(_13147_ ), .A3(\wbu.rf_29 [22] ), .A4(_13327_ ), .ZN(_00926_ ) );
NAND4_X1 _21480_ ( .A1(_13105_ ), .A2(_13350_ ), .A3(fanout_net_36 ), .A4(\wbu.rf_19 [22] ), .ZN(_00927_ ) );
AND4_X1 _21481_ ( .A1(fanout_net_36 ), .A2(_13173_ ), .A3(\wbu.rf_18 [22] ), .A4(_08573_ ), .ZN(_00928_ ) );
NAND3_X1 _21482_ ( .A1(_13026_ ), .A2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A3(\wbu.rf_8 [22] ), .ZN(_00929_ ) );
AND4_X1 _21483_ ( .A1(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .A2(_12977_ ), .A3(_13007_ ), .A4(\wbu.rf_6 [22] ), .ZN(_00930_ ) );
MUX2_X1 _21484_ ( .A(\wbu._GEN_71 [22] ), .B(\wbu.rf_2 [22] ), .S(_12992_ ), .Z(_00931_ ) );
MUX2_X1 _21485_ ( .A(\wbu.rf_3 [22] ), .B(_00931_ ), .S(_12997_ ), .Z(_00932_ ) );
MUX2_X1 _21486_ ( .A(\wbu.rf_4 [22] ), .B(_00932_ ), .S(_13003_ ), .Z(_00933_ ) );
MUX2_X1 _21487_ ( .A(\wbu.rf_5 [22] ), .B(_00933_ ), .S(_13011_ ), .Z(_00934_ ) );
AOI211_X1 _21488_ ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_Y ), .B(_00930_ ), .C1(_00934_ ), .C2(_13017_ ), .ZN(_00935_ ) );
OAI21_X1 _21489_ ( .A(_13028_ ), .B1(_13022_ ), .B2(\wbu.rf_7 [22] ), .ZN(_00936_ ) );
OAI21_X1 _21490_ ( .A(_00929_ ), .B1(_00935_ ), .B2(_00936_ ), .ZN(_00937_ ) );
MUX2_X1 _21491_ ( .A(\wbu.rf_9 [22] ), .B(_00937_ ), .S(_13198_ ), .Z(_00938_ ) );
MUX2_X1 _21492_ ( .A(\wbu.rf_10 [22] ), .B(_00938_ ), .S(_12983_ ), .Z(_00939_ ) );
MUX2_X1 _21493_ ( .A(\wbu.rf_11 [22] ), .B(_00939_ ), .S(_13037_ ), .Z(_00940_ ) );
MUX2_X1 _21494_ ( .A(\wbu.rf_12 [22] ), .B(_00940_ ), .S(_13044_ ), .Z(_00941_ ) );
MUX2_X1 _21495_ ( .A(\wbu.rf_13 [22] ), .B(_00941_ ), .S(_13053_ ), .Z(_00942_ ) );
MUX2_X1 _21496_ ( .A(\wbu.rf_14 [22] ), .B(_00942_ ), .S(_13058_ ), .Z(_00943_ ) );
MUX2_X1 _21497_ ( .A(\wbu.rf_15 [22] ), .B(_00943_ ), .S(_13069_ ), .Z(_00944_ ) );
MUX2_X1 _21498_ ( .A(\wbu.rf_16 [22] ), .B(_00944_ ), .S(_13074_ ), .Z(_00945_ ) );
MUX2_X1 _21499_ ( .A(\wbu.rf_17 [22] ), .B(_00945_ ), .S(_13084_ ), .Z(_00946_ ) );
AOI21_X1 _21500_ ( .A(_00928_ ), .B1(_00946_ ), .B2(_13090_ ), .ZN(_00947_ ) );
OAI211_X1 _21501_ ( .A(_13103_ ), .B(_00927_ ), .C1(_00947_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .ZN(_00948_ ) );
OAI211_X1 _21502_ ( .A(_00948_ ), .B(_13110_ ), .C1(\wbu.rf_20 [22] ), .C2(_13103_ ), .ZN(_00949_ ) );
NAND4_X1 _21503_ ( .A1(_13119_ ), .A2(_13121_ ), .A3(fanout_net_36 ), .A4(\wbu.rf_21 [22] ), .ZN(_00950_ ) );
NAND3_X1 _21504_ ( .A1(_00949_ ), .A2(_13116_ ), .A3(_00950_ ), .ZN(_00951_ ) );
OAI211_X1 _21505_ ( .A(_00951_ ), .B(_13126_ ), .C1(\wbu.rf_22 [22] ), .C2(_13116_ ), .ZN(_00952_ ) );
NAND4_X1 _21506_ ( .A1(_13188_ ), .A2(fanout_net_36 ), .A3(_13134_ ), .A4(\wbu.rf_23 [22] ), .ZN(_00953_ ) );
NAND3_X1 _21507_ ( .A1(_00952_ ), .A2(_13130_ ), .A3(_00953_ ), .ZN(_00954_ ) );
OAI211_X1 _21508_ ( .A(_00954_ ), .B(_13139_ ), .C1(\wbu.rf_24 [22] ), .C2(_13131_ ), .ZN(_00955_ ) );
NAND4_X1 _21509_ ( .A1(_13146_ ), .A2(_13148_ ), .A3(fanout_net_36 ), .A4(\wbu.rf_25 [22] ), .ZN(_00956_ ) );
NAND2_X1 _21510_ ( .A1(_00955_ ), .A2(_00956_ ), .ZN(_00957_ ) );
MUX2_X1 _21511_ ( .A(\wbu.rf_26 [22] ), .B(_00957_ ), .S(_13143_ ), .Z(_00958_ ) );
MUX2_X1 _21512_ ( .A(\wbu.rf_27 [22] ), .B(_00958_ ), .S(_13363_ ), .Z(_00959_ ) );
MUX2_X1 _21513_ ( .A(\wbu.rf_28 [22] ), .B(_00959_ ), .S(_13157_ ), .Z(_00960_ ) );
AOI21_X1 _21514_ ( .A(_00926_ ), .B1(_00960_ ), .B2(_13269_ ), .ZN(_00961_ ) );
OAI211_X1 _21515_ ( .A(_12971_ ), .B(_00925_ ), .C1(_00961_ ), .C2(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .ZN(_00962_ ) );
OR2_X1 _21516_ ( .A1(_13369_ ), .A2(\wbu.rf_31 [22] ), .ZN(_00963_ ) );
AOI21_X1 _21517_ ( .A(_13473_ ), .B1(_00962_ ), .B2(_00963_ ), .ZN(_00964_ ) );
INV_X1 _21518_ ( .A(\wbu.io_in_bits_rd_wdata [22] ), .ZN(_00965_ ) );
AOI211_X1 _21519_ ( .A(fanout_net_25 ), .B(_00964_ ), .C1(_00965_ ), .C2(_13324_ ), .ZN(_00377_ ) );
NOR2_X1 _21520_ ( .A1(_12958_ ), .A2(fanout_net_25 ), .ZN(_00378_ ) );
NOR2_X1 _21521_ ( .A1(_13185_ ), .A2(fanout_net_25 ), .ZN(_00379_ ) );
AND2_X1 _21522_ ( .A1(\ifu.ren_REG_$_DFF_P__Q_D_$_NAND__Y_B ), .A2(\wbu.io_in_bits_rd_wdata [21] ), .ZN(_00380_ ) );
NOR2_X1 _21523_ ( .A1(_13279_ ), .A2(fanout_net_25 ), .ZN(_00381_ ) );
NOR2_X1 _21524_ ( .A1(_13372_ ), .A2(fanout_net_25 ), .ZN(_00382_ ) );
AND2_X1 _21525_ ( .A1(\ifu.ren_REG_$_DFF_P__Q_D_$_NAND__Y_B ), .A2(\wbu.io_in_bits_rd_wdata [18] ), .ZN(_00383_ ) );
NOR2_X1 _21526_ ( .A1(_13427_ ), .A2(fanout_net_25 ), .ZN(_00384_ ) );
NOR2_X1 _21527_ ( .A1(_13518_ ), .A2(fanout_net_25 ), .ZN(_00385_ ) );
NOR2_X1 _21528_ ( .A1(_13519_ ), .A2(fanout_net_25 ), .ZN(_00386_ ) );
NOR2_X1 _21529_ ( .A1(_13592_ ), .A2(fanout_net_25 ), .ZN(_00387_ ) );
NOR2_X1 _21530_ ( .A1(_13629_ ), .A2(fanout_net_25 ), .ZN(_00388_ ) );
NOR2_X1 _21531_ ( .A1(_13676_ ), .A2(fanout_net_25 ), .ZN(_00389_ ) );
NOR2_X1 _21532_ ( .A1(_13718_ ), .A2(fanout_net_25 ), .ZN(_00390_ ) );
NOR2_X1 _21533_ ( .A1(_13719_ ), .A2(fanout_net_25 ), .ZN(_00391_ ) );
NOR2_X1 _21534_ ( .A1(_13756_ ), .A2(fanout_net_25 ), .ZN(_00392_ ) );
NOR2_X1 _21535_ ( .A1(_13799_ ), .A2(fanout_net_25 ), .ZN(_00393_ ) );
AND2_X1 _21536_ ( .A1(\ifu.ren_REG_$_DFF_P__Q_D_$_NAND__Y_B ), .A2(\wbu.io_in_bits_rd_wdata [8] ), .ZN(_00394_ ) );
NOR2_X1 _21537_ ( .A1(_13919_ ), .A2(fanout_net_25 ), .ZN(_00395_ ) );
AND2_X1 _21538_ ( .A1(\ifu.ren_REG_$_DFF_P__Q_D_$_NAND__Y_B ), .A2(\wbu.io_in_bits_rd_wdata [6] ), .ZN(_00396_ ) );
NOR2_X1 _21539_ ( .A1(_00484_ ), .A2(fanout_net_25 ), .ZN(_00397_ ) );
NOR2_X1 _21540_ ( .A1(_00485_ ), .A2(fanout_net_25 ), .ZN(_00398_ ) );
NOR2_X1 _21541_ ( .A1(_00566_ ), .A2(fanout_net_25 ), .ZN(_00399_ ) );
INV_X1 _21542_ ( .A(\wbu.io_in_bits_rd_wdata [2] ), .ZN(_00966_ ) );
NOR2_X1 _21543_ ( .A1(_00966_ ), .A2(fanout_net_26 ), .ZN(_00400_ ) );
NOR2_X1 _21544_ ( .A1(_00639_ ), .A2(fanout_net_26 ), .ZN(_00401_ ) );
NOR2_X1 _21545_ ( .A1(_00640_ ), .A2(fanout_net_26 ), .ZN(_00402_ ) );
AND2_X1 _21546_ ( .A1(_10987_ ), .A2(\wbu.io_in_bits_rd_wdata [0] ), .ZN(_00403_ ) );
NOR2_X1 _21547_ ( .A1(_00771_ ), .A2(fanout_net_26 ), .ZN(_00404_ ) );
NOR2_X1 _21548_ ( .A1(_00808_ ), .A2(fanout_net_26 ), .ZN(_00405_ ) );
NOR2_X1 _21549_ ( .A1(_00845_ ), .A2(fanout_net_26 ), .ZN(_00406_ ) );
NOR2_X1 _21550_ ( .A1(_00885_ ), .A2(fanout_net_26 ), .ZN(_00407_ ) );
AND2_X1 _21551_ ( .A1(_10987_ ), .A2(\wbu.io_in_bits_rd_wdata [23] ), .ZN(_00408_ ) );
NOR2_X1 _21552_ ( .A1(_00965_ ), .A2(fanout_net_26 ), .ZN(_00409_ ) );
AOI21_X1 _21553_ ( .A(fanout_net_26 ), .B1(_08567_ ), .B2(_08569_ ), .ZN(_00410_ ) );
BUF_X2 _21554_ ( .A(_08547_ ), .Z(_00967_ ) );
BUF_X2 _21555_ ( .A(_00967_ ), .Z(_00968_ ) );
BUF_X2 _21556_ ( .A(_08560_ ), .Z(_00969_ ) );
BUF_X2 _21557_ ( .A(_00969_ ), .Z(_00970_ ) );
NOR2_X1 _21558_ ( .A1(_10823_ ), .A2(\lsu.state [1] ), .ZN(_00971_ ) );
NOR2_X1 _21559_ ( .A1(_00971_ ), .A2(io_master_wready_$_ANDNOT__B_Y_$_OR__A_B ), .ZN(_00972_ ) );
INV_X1 _21560_ ( .A(_00972_ ), .ZN(_00973_ ) );
NOR3_X1 _21561_ ( .A1(_00968_ ), .A2(_00970_ ), .A3(_00973_ ), .ZN(\arbiter.clink.io_axi_arvalid ) );
BUF_X4 _21562_ ( .A(_08562_ ), .Z(_00974_ ) );
BUF_X4 _21563_ ( .A(_00974_ ), .Z(_00975_ ) );
BUF_X4 _21564_ ( .A(_00972_ ), .Z(_00976_ ) );
BUF_X4 _21565_ ( .A(_00976_ ), .Z(_00977_ ) );
NAND4_X1 _21566_ ( .A1(_00975_ ), .A2(\arbiter.clink.mtime [63] ), .A3(\io_master_awaddr [2] ), .A4(_00977_ ), .ZN(_00978_ ) );
BUF_X4 _21567_ ( .A(_00974_ ), .Z(_00979_ ) );
INV_X1 _21568_ ( .A(\io_master_awaddr [2] ), .ZN(_00980_ ) );
BUF_X4 _21569_ ( .A(_00980_ ), .Z(_00981_ ) );
BUF_X4 _21570_ ( .A(_00976_ ), .Z(_00982_ ) );
NAND4_X1 _21571_ ( .A1(_00979_ ), .A2(\arbiter.clink.mtime [31] ), .A3(_00981_ ), .A4(_00982_ ), .ZN(_00983_ ) );
NAND2_X1 _21572_ ( .A1(_00978_ ), .A2(_00983_ ), .ZN(_00002_ ) );
NAND4_X1 _21573_ ( .A1(_00975_ ), .A2(\arbiter.clink.mtime [62] ), .A3(\io_master_awaddr [2] ), .A4(_00977_ ), .ZN(_00984_ ) );
NAND4_X1 _21574_ ( .A1(_00979_ ), .A2(\arbiter.clink.mtime [30] ), .A3(_00981_ ), .A4(_00982_ ), .ZN(_00985_ ) );
NAND2_X1 _21575_ ( .A1(_00984_ ), .A2(_00985_ ), .ZN(_00003_ ) );
NAND4_X1 _21576_ ( .A1(_00975_ ), .A2(\arbiter.clink.mtime [53] ), .A3(\io_master_awaddr [2] ), .A4(_00977_ ), .ZN(_00986_ ) );
NAND4_X1 _21577_ ( .A1(_00979_ ), .A2(\arbiter.clink.mtime [21] ), .A3(_00981_ ), .A4(_00982_ ), .ZN(_00987_ ) );
NAND2_X1 _21578_ ( .A1(_00986_ ), .A2(_00987_ ), .ZN(_00004_ ) );
NAND4_X1 _21579_ ( .A1(_00975_ ), .A2(\arbiter.clink.mtime [52] ), .A3(\io_master_awaddr [2] ), .A4(_00977_ ), .ZN(_00988_ ) );
NAND4_X1 _21580_ ( .A1(_00979_ ), .A2(\arbiter.clink.mtime [20] ), .A3(_00981_ ), .A4(_00982_ ), .ZN(_00989_ ) );
NAND2_X1 _21581_ ( .A1(_00988_ ), .A2(_00989_ ), .ZN(_00005_ ) );
NAND4_X1 _21582_ ( .A1(_00975_ ), .A2(\arbiter.clink.mtime [51] ), .A3(\io_master_awaddr [2] ), .A4(_00977_ ), .ZN(_00990_ ) );
NAND4_X1 _21583_ ( .A1(_00979_ ), .A2(\arbiter.clink.mtime [19] ), .A3(_00981_ ), .A4(_00982_ ), .ZN(_00991_ ) );
NAND2_X1 _21584_ ( .A1(_00990_ ), .A2(_00991_ ), .ZN(_00006_ ) );
NAND4_X1 _21585_ ( .A1(_00975_ ), .A2(\arbiter.clink.mtime [50] ), .A3(\io_master_awaddr [2] ), .A4(_00977_ ), .ZN(_00992_ ) );
NAND4_X1 _21586_ ( .A1(_00979_ ), .A2(\arbiter.clink.mtime [18] ), .A3(_00981_ ), .A4(_00982_ ), .ZN(_00993_ ) );
NAND2_X1 _21587_ ( .A1(_00992_ ), .A2(_00993_ ), .ZN(_00007_ ) );
NAND4_X1 _21588_ ( .A1(_00975_ ), .A2(\arbiter.clink.mtime [49] ), .A3(\io_master_awaddr [2] ), .A4(_00977_ ), .ZN(_00994_ ) );
NAND4_X1 _21589_ ( .A1(_00979_ ), .A2(\arbiter.clink.mtime [17] ), .A3(_00981_ ), .A4(_00982_ ), .ZN(_00995_ ) );
NAND2_X1 _21590_ ( .A1(_00994_ ), .A2(_00995_ ), .ZN(_00008_ ) );
NAND4_X1 _21591_ ( .A1(_00975_ ), .A2(\arbiter.clink.mtime [48] ), .A3(\io_master_awaddr [2] ), .A4(_00977_ ), .ZN(_00996_ ) );
NAND4_X1 _21592_ ( .A1(_00979_ ), .A2(\arbiter.clink.mtime [16] ), .A3(_00981_ ), .A4(_00982_ ), .ZN(_00997_ ) );
NAND2_X1 _21593_ ( .A1(_00996_ ), .A2(_00997_ ), .ZN(_00009_ ) );
NAND4_X1 _21594_ ( .A1(_00975_ ), .A2(\arbiter.clink.mtime [47] ), .A3(\io_master_awaddr [2] ), .A4(_00977_ ), .ZN(_00998_ ) );
BUF_X4 _21595_ ( .A(_00974_ ), .Z(_00999_ ) );
BUF_X4 _21596_ ( .A(_00976_ ), .Z(_01000_ ) );
NAND4_X1 _21597_ ( .A1(_00999_ ), .A2(\arbiter.clink.mtime [15] ), .A3(_00981_ ), .A4(_01000_ ), .ZN(_01001_ ) );
NAND2_X1 _21598_ ( .A1(_00998_ ), .A2(_01001_ ), .ZN(_00010_ ) );
NAND4_X1 _21599_ ( .A1(_00975_ ), .A2(\arbiter.clink.mtime [46] ), .A3(\io_master_awaddr [2] ), .A4(_00977_ ), .ZN(_01002_ ) );
BUF_X4 _21600_ ( .A(_00980_ ), .Z(_01003_ ) );
NAND4_X1 _21601_ ( .A1(_00999_ ), .A2(\arbiter.clink.mtime [14] ), .A3(_01003_ ), .A4(_01000_ ), .ZN(_01004_ ) );
NAND2_X1 _21602_ ( .A1(_01002_ ), .A2(_01004_ ), .ZN(_00011_ ) );
BUF_X4 _21603_ ( .A(_00974_ ), .Z(_01005_ ) );
BUF_X4 _21604_ ( .A(_00976_ ), .Z(_01006_ ) );
NAND4_X1 _21605_ ( .A1(_01005_ ), .A2(\arbiter.clink.mtime [45] ), .A3(\io_master_awaddr [2] ), .A4(_01006_ ), .ZN(_01007_ ) );
NAND4_X1 _21606_ ( .A1(_00999_ ), .A2(\arbiter.clink.mtime [13] ), .A3(_01003_ ), .A4(_01000_ ), .ZN(_01008_ ) );
NAND2_X1 _21607_ ( .A1(_01007_ ), .A2(_01008_ ), .ZN(_00012_ ) );
NAND4_X1 _21608_ ( .A1(_01005_ ), .A2(\arbiter.clink.mtime [44] ), .A3(\io_master_awaddr [2] ), .A4(_01006_ ), .ZN(_01009_ ) );
NAND4_X1 _21609_ ( .A1(_00999_ ), .A2(\arbiter.clink.mtime [12] ), .A3(_01003_ ), .A4(_01000_ ), .ZN(_01010_ ) );
NAND2_X1 _21610_ ( .A1(_01009_ ), .A2(_01010_ ), .ZN(_00013_ ) );
NAND4_X1 _21611_ ( .A1(_01005_ ), .A2(\arbiter.clink.mtime [61] ), .A3(\io_master_awaddr [2] ), .A4(_01006_ ), .ZN(_01011_ ) );
NAND4_X1 _21612_ ( .A1(_00999_ ), .A2(\arbiter.clink.mtime [29] ), .A3(_01003_ ), .A4(_01000_ ), .ZN(_01012_ ) );
NAND2_X1 _21613_ ( .A1(_01011_ ), .A2(_01012_ ), .ZN(_00014_ ) );
NAND4_X1 _21614_ ( .A1(_01005_ ), .A2(\arbiter.clink.mtime [43] ), .A3(\io_master_awaddr [2] ), .A4(_01006_ ), .ZN(_01013_ ) );
NAND4_X1 _21615_ ( .A1(_00999_ ), .A2(\arbiter.clink.mtime [11] ), .A3(_01003_ ), .A4(_01000_ ), .ZN(_01014_ ) );
NAND2_X1 _21616_ ( .A1(_01013_ ), .A2(_01014_ ), .ZN(_00015_ ) );
NAND4_X1 _21617_ ( .A1(_01005_ ), .A2(\arbiter.clink.mtime [42] ), .A3(\io_master_awaddr [2] ), .A4(_01006_ ), .ZN(_01015_ ) );
NAND4_X1 _21618_ ( .A1(_00999_ ), .A2(\arbiter.clink.mtime [10] ), .A3(_01003_ ), .A4(_01000_ ), .ZN(_01016_ ) );
NAND2_X1 _21619_ ( .A1(_01015_ ), .A2(_01016_ ), .ZN(_00016_ ) );
NAND4_X1 _21620_ ( .A1(_01005_ ), .A2(\arbiter.clink.mtime [41] ), .A3(\io_master_awaddr [2] ), .A4(_01006_ ), .ZN(_01017_ ) );
NAND4_X1 _21621_ ( .A1(_00999_ ), .A2(\arbiter.clink.mtime [9] ), .A3(_01003_ ), .A4(_01000_ ), .ZN(_01018_ ) );
NAND2_X1 _21622_ ( .A1(_01017_ ), .A2(_01018_ ), .ZN(_00017_ ) );
NAND4_X1 _21623_ ( .A1(_01005_ ), .A2(\arbiter.clink.mtime [40] ), .A3(\io_master_awaddr [2] ), .A4(_01006_ ), .ZN(_01019_ ) );
NAND4_X1 _21624_ ( .A1(_00999_ ), .A2(\arbiter.clink.mtime [8] ), .A3(_01003_ ), .A4(_01000_ ), .ZN(_01020_ ) );
NAND2_X1 _21625_ ( .A1(_01019_ ), .A2(_01020_ ), .ZN(_00018_ ) );
NAND4_X1 _21626_ ( .A1(_01005_ ), .A2(\arbiter.clink.mtime [39] ), .A3(\io_master_awaddr [2] ), .A4(_01006_ ), .ZN(_01021_ ) );
NAND4_X1 _21627_ ( .A1(_00999_ ), .A2(\arbiter.clink.mtime [7] ), .A3(_01003_ ), .A4(_01000_ ), .ZN(_01022_ ) );
NAND2_X1 _21628_ ( .A1(_01021_ ), .A2(_01022_ ), .ZN(_00019_ ) );
NAND4_X1 _21629_ ( .A1(_01005_ ), .A2(\arbiter.clink.mtime [38] ), .A3(\io_master_awaddr [2] ), .A4(_01006_ ), .ZN(_01023_ ) );
BUF_X4 _21630_ ( .A(_00974_ ), .Z(_01024_ ) );
BUF_X4 _21631_ ( .A(_00976_ ), .Z(_01025_ ) );
NAND4_X1 _21632_ ( .A1(_01024_ ), .A2(\arbiter.clink.mtime [6] ), .A3(_01003_ ), .A4(_01025_ ), .ZN(_01026_ ) );
NAND2_X1 _21633_ ( .A1(_01023_ ), .A2(_01026_ ), .ZN(_00020_ ) );
NAND4_X1 _21634_ ( .A1(_01005_ ), .A2(\arbiter.clink.mtime [37] ), .A3(\io_master_awaddr [2] ), .A4(_01006_ ), .ZN(_01027_ ) );
BUF_X4 _21635_ ( .A(_00980_ ), .Z(_01028_ ) );
NAND4_X1 _21636_ ( .A1(_01024_ ), .A2(\arbiter.clink.mtime [5] ), .A3(_01028_ ), .A4(_01025_ ), .ZN(_01029_ ) );
NAND2_X1 _21637_ ( .A1(_01027_ ), .A2(_01029_ ), .ZN(_00021_ ) );
BUF_X4 _21638_ ( .A(_00974_ ), .Z(_01030_ ) );
BUF_X4 _21639_ ( .A(_00976_ ), .Z(_01031_ ) );
NAND4_X1 _21640_ ( .A1(_01030_ ), .A2(\arbiter.clink.mtime [36] ), .A3(\io_master_awaddr [2] ), .A4(_01031_ ), .ZN(_01032_ ) );
NAND4_X1 _21641_ ( .A1(_01024_ ), .A2(\arbiter.clink.mtime [4] ), .A3(_01028_ ), .A4(_01025_ ), .ZN(_01033_ ) );
NAND2_X1 _21642_ ( .A1(_01032_ ), .A2(_01033_ ), .ZN(_00022_ ) );
NAND4_X1 _21643_ ( .A1(_01030_ ), .A2(\arbiter.clink.mtime [35] ), .A3(\io_master_awaddr [2] ), .A4(_01031_ ), .ZN(_01034_ ) );
NAND4_X1 _21644_ ( .A1(_01024_ ), .A2(\arbiter.clink.mtime [3] ), .A3(_01028_ ), .A4(_01025_ ), .ZN(_01035_ ) );
NAND2_X1 _21645_ ( .A1(_01034_ ), .A2(_01035_ ), .ZN(_00023_ ) );
NAND4_X1 _21646_ ( .A1(_01030_ ), .A2(\arbiter.clink.mtime [34] ), .A3(\io_master_awaddr [2] ), .A4(_01031_ ), .ZN(_01036_ ) );
NAND4_X1 _21647_ ( .A1(_01024_ ), .A2(\arbiter.clink.mtime [2] ), .A3(_01028_ ), .A4(_01025_ ), .ZN(_01037_ ) );
NAND2_X1 _21648_ ( .A1(_01036_ ), .A2(_01037_ ), .ZN(_00024_ ) );
NAND4_X1 _21649_ ( .A1(_01030_ ), .A2(\arbiter.clink.mtime [60] ), .A3(\io_master_awaddr [2] ), .A4(_01031_ ), .ZN(_01038_ ) );
NAND4_X1 _21650_ ( .A1(_01024_ ), .A2(\arbiter.clink.mtime [28] ), .A3(_01028_ ), .A4(_01025_ ), .ZN(_01039_ ) );
NAND2_X1 _21651_ ( .A1(_01038_ ), .A2(_01039_ ), .ZN(_00025_ ) );
NAND4_X1 _21652_ ( .A1(_01030_ ), .A2(\arbiter.clink.mtime [33] ), .A3(\io_master_awaddr [2] ), .A4(_01031_ ), .ZN(_01040_ ) );
NAND4_X1 _21653_ ( .A1(_01024_ ), .A2(\arbiter.clink.mtime [1] ), .A3(_01028_ ), .A4(_01025_ ), .ZN(_01041_ ) );
NAND2_X1 _21654_ ( .A1(_01040_ ), .A2(_01041_ ), .ZN(_00026_ ) );
NAND4_X1 _21655_ ( .A1(_01030_ ), .A2(\arbiter.clink.mtime [32] ), .A3(\io_master_awaddr [2] ), .A4(_01031_ ), .ZN(_01042_ ) );
NAND4_X1 _21656_ ( .A1(_01024_ ), .A2(\arbiter.clink.mtime [0] ), .A3(_01028_ ), .A4(_01025_ ), .ZN(_01043_ ) );
NAND2_X1 _21657_ ( .A1(_01042_ ), .A2(_01043_ ), .ZN(_00027_ ) );
NAND4_X1 _21658_ ( .A1(_01030_ ), .A2(\arbiter.clink.mtime [59] ), .A3(\io_master_awaddr [2] ), .A4(_01031_ ), .ZN(_01044_ ) );
NAND4_X1 _21659_ ( .A1(_01024_ ), .A2(\arbiter.clink.mtime [27] ), .A3(_01028_ ), .A4(_01025_ ), .ZN(_01045_ ) );
NAND2_X1 _21660_ ( .A1(_01044_ ), .A2(_01045_ ), .ZN(_00028_ ) );
NAND4_X1 _21661_ ( .A1(_01030_ ), .A2(\arbiter.clink.mtime [58] ), .A3(\io_master_awaddr [2] ), .A4(_01031_ ), .ZN(_01046_ ) );
NAND4_X1 _21662_ ( .A1(_01024_ ), .A2(\arbiter.clink.mtime [26] ), .A3(_01028_ ), .A4(_01025_ ), .ZN(_01047_ ) );
NAND2_X1 _21663_ ( .A1(_01046_ ), .A2(_01047_ ), .ZN(_00029_ ) );
NAND4_X1 _21664_ ( .A1(_01030_ ), .A2(\arbiter.clink.mtime [57] ), .A3(fanout_net_16 ), .A4(_01031_ ), .ZN(_01048_ ) );
NAND4_X1 _21665_ ( .A1(_00974_ ), .A2(\arbiter.clink.mtime [25] ), .A3(_01028_ ), .A4(_00976_ ), .ZN(_01049_ ) );
NAND2_X1 _21666_ ( .A1(_01048_ ), .A2(_01049_ ), .ZN(_00030_ ) );
NAND4_X1 _21667_ ( .A1(_01030_ ), .A2(\arbiter.clink.mtime [56] ), .A3(fanout_net_16 ), .A4(_01031_ ), .ZN(_01050_ ) );
NAND4_X1 _21668_ ( .A1(_00974_ ), .A2(\arbiter.clink.mtime [24] ), .A3(_00980_ ), .A4(_00976_ ), .ZN(_01051_ ) );
NAND2_X1 _21669_ ( .A1(_01050_ ), .A2(_01051_ ), .ZN(_00031_ ) );
NAND4_X1 _21670_ ( .A1(_00979_ ), .A2(\arbiter.clink.mtime [55] ), .A3(fanout_net_16 ), .A4(_00982_ ), .ZN(_01052_ ) );
NAND4_X1 _21671_ ( .A1(_00974_ ), .A2(\arbiter.clink.mtime [23] ), .A3(_00980_ ), .A4(_00976_ ), .ZN(_01053_ ) );
NAND2_X1 _21672_ ( .A1(_01052_ ), .A2(_01053_ ), .ZN(_00032_ ) );
NAND4_X1 _21673_ ( .A1(_00979_ ), .A2(\arbiter.clink.mtime [54] ), .A3(fanout_net_16 ), .A4(_00982_ ), .ZN(_01054_ ) );
NAND4_X1 _21674_ ( .A1(_00974_ ), .A2(\arbiter.clink.mtime [22] ), .A3(_00980_ ), .A4(_00976_ ), .ZN(_01055_ ) );
NAND2_X1 _21675_ ( .A1(_01054_ ), .A2(_01055_ ), .ZN(_00033_ ) );
NOR2_X1 _21676_ ( .A1(_10824_ ), .A2(\lsu._io_axi_awvalid_T_1 ), .ZN(_01056_ ) );
AND2_X1 _21677_ ( .A1(_00971_ ), .A2(_01056_ ), .ZN(_01057_ ) );
BUF_X2 _21678_ ( .A(_10844_ ), .Z(_01058_ ) );
AND3_X1 _21679_ ( .A1(_01057_ ), .A2(_01058_ ), .A3(\arbiter._clink_io_axi_araddr_T ), .ZN(_01059_ ) );
INV_X1 _21680_ ( .A(_11977_ ), .ZN(_01060_ ) );
AOI21_X1 _21681_ ( .A(_10703_ ), .B1(_01060_ ), .B2(_12018_ ), .ZN(_01061_ ) );
OAI221_X1 _21682_ ( .A(_01059_ ), .B1(_12204_ ), .B2(_12019_ ), .C1(_01061_ ), .C2(\icache._io_out_arvalid_T_2 ), .ZN(_01062_ ) );
INV_X1 _21683_ ( .A(\arbiter._io_axi_araddr_T_6 ), .ZN(_01063_ ) );
BUF_X4 _21684_ ( .A(_01063_ ), .Z(_01064_ ) );
BUF_X2 _21685_ ( .A(_01064_ ), .Z(_01065_ ) );
OR3_X1 _21686_ ( .A1(_01065_ ), .A2(fanout_net_26 ), .A3(\arbiter.ifu_end ), .ZN(_01066_ ) );
NAND2_X1 _21687_ ( .A1(_01062_ ), .A2(_01066_ ), .ZN(\arbiter.state_$_DFF_P__Q_1_D ) );
NOR2_X1 _21688_ ( .A1(_01061_ ), .A2(\icache._io_out_arvalid_T_2 ), .ZN(_01067_ ) );
OAI21_X1 _21689_ ( .A(_01059_ ), .B1(_01067_ ), .B2(_10708_ ), .ZN(_01068_ ) );
AOI221_X4 _21690_ ( .A(fanout_net_26 ), .B1(\arbiter.ifu_end ), .B2(\arbiter._io_axi_araddr_T_6 ), .C1(\arbiter.lsu_end ), .C2(fanout_net_1 ), .ZN(_01069_ ) );
NAND2_X1 _21691_ ( .A1(_01068_ ), .A2(_01069_ ), .ZN(\arbiter.state_$_DFF_P__Q_2_D ) );
INV_X1 _21692_ ( .A(\arbiter.lsu_end ), .ZN(_01070_ ) );
NAND3_X1 _21693_ ( .A1(_10979_ ), .A2(_01070_ ), .A3(fanout_net_1 ), .ZN(_01071_ ) );
NAND2_X1 _21694_ ( .A1(_10917_ ), .A2(\arbiter._clink_io_axi_araddr_T ), .ZN(_01072_ ) );
OAI21_X1 _21695_ ( .A(_01071_ ), .B1(_01057_ ), .B2(_01072_ ), .ZN(\arbiter.state_$_DFF_P__Q_D ) );
INV_X1 _21696_ ( .A(_10093_ ), .ZN(\exu.addi._io_rd_T_4 [17] ) );
INV_X1 _21697_ ( .A(_11473_ ), .ZN(\exu.addi._io_rd_T_4 [3] ) );
BUF_X4 _21698_ ( .A(_11397_ ), .Z(\exu._io_out_bits_wdata_T_1 [3] ) );
NOR2_X1 _21699_ ( .A1(_09553_ ), .A2(_09514_ ), .ZN(\exu.addi._io_rd_T_4 [22] ) );
MUX2_X1 _21700_ ( .A(\exu._GEN_0 [31] ), .B(\exu._GEN_0 [23] ), .S(\exu._io_out_bits_wdata_T_1 [3] ), .Z(_01073_ ) );
MUX2_X1 _21701_ ( .A(_01073_ ), .B(_12824_ ), .S(\exu._io_out_bits_wdata_T_1 [4] ), .Z(\exu._io_out_bits_wdata_T_2 [31] ) );
MUX2_X1 _21702_ ( .A(\exu._GEN_0 [30] ), .B(\exu._GEN_0 [22] ), .S(\exu._io_out_bits_wdata_T_1 [3] ), .Z(_01074_ ) );
MUX2_X1 _21703_ ( .A(_01074_ ), .B(_12826_ ), .S(\exu._io_out_bits_wdata_T_1 [4] ), .Z(\exu._io_out_bits_wdata_T_2 [30] ) );
NAND3_X1 _21704_ ( .A1(\exu._io_out_bits_wdata_T_1 [4] ), .A2(\exu._GEN_0 [5] ), .A3(_12828_ ), .ZN(_01075_ ) );
MUX2_X1 _21705_ ( .A(_08895_ ), .B(_08857_ ), .S(\exu._io_out_bits_wdata_T_1 [3] ), .Z(_01076_ ) );
OAI21_X1 _21706_ ( .A(_01075_ ), .B1(_01076_ ), .B2(\exu._io_out_bits_wdata_T_1 [4] ), .ZN(\exu._io_out_bits_wdata_T_2 [21] ) );
MUX2_X1 _21707_ ( .A(\exu._GEN_0 [20] ), .B(\exu._GEN_0 [12] ), .S(\exu._io_out_bits_wdata_T_1 [3] ), .Z(_01077_ ) );
BUF_X4 _21708_ ( .A(_11358_ ), .Z(_01078_ ) );
MUX2_X1 _21709_ ( .A(_01077_ ), .B(_12830_ ), .S(_01078_ ), .Z(\exu._io_out_bits_wdata_T_2 [20] ) );
OR2_X1 _21710_ ( .A1(\exu._io_out_bits_wdata_T_1 [3] ), .A2(\exu._GEN_0 [19] ), .ZN(_01079_ ) );
OAI211_X1 _21711_ ( .A(_12825_ ), .B(_01079_ ), .C1(\exu._GEN_0 [11] ), .C2(_12828_ ), .ZN(_01080_ ) );
NAND3_X1 _21712_ ( .A1(\exu._io_out_bits_wdata_T_1 [4] ), .A2(_12831_ ), .A3(_12828_ ), .ZN(_01081_ ) );
NAND2_X1 _21713_ ( .A1(_01080_ ), .A2(_01081_ ), .ZN(\exu._io_out_bits_wdata_T_2 [19] ) );
NAND3_X1 _21714_ ( .A1(\exu._io_out_bits_wdata_T_1 [4] ), .A2(_12832_ ), .A3(_12828_ ), .ZN(_01082_ ) );
INV_X1 _21715_ ( .A(\exu._GEN_0 [18] ), .ZN(_01083_ ) );
INV_X1 _21716_ ( .A(\exu._GEN_0 [10] ), .ZN(_01084_ ) );
MUX2_X1 _21717_ ( .A(_01083_ ), .B(_01084_ ), .S(\exu._io_out_bits_wdata_T_1 [3] ), .Z(_01085_ ) );
OAI21_X1 _21718_ ( .A(_01082_ ), .B1(_01085_ ), .B2(\exu._io_out_bits_wdata_T_1 [4] ), .ZN(\exu._io_out_bits_wdata_T_2 [18] ) );
NAND3_X1 _21719_ ( .A1(\exu._io_out_bits_wdata_T_1 [4] ), .A2(_12833_ ), .A3(_12828_ ), .ZN(_01086_ ) );
MUX2_X1 _21720_ ( .A(_08879_ ), .B(_08845_ ), .S(\exu._io_out_bits_wdata_T_1 [3] ), .Z(_01087_ ) );
OAI21_X1 _21721_ ( .A(_01086_ ), .B1(_01087_ ), .B2(\exu._io_out_bits_wdata_T_1 [4] ), .ZN(\exu._io_out_bits_wdata_T_2 [17] ) );
MUX2_X1 _21722_ ( .A(\exu._GEN_0 [16] ), .B(\exu._GEN_0 [8] ), .S(\exu._io_out_bits_wdata_T_1 [3] ), .Z(_01088_ ) );
INV_X1 _21723_ ( .A(\exu._GEN_0 [0] ), .ZN(_01089_ ) );
AOI21_X1 _21724_ ( .A(_01089_ ), .B1(_09054_ ), .B2(_12829_ ), .ZN(_01090_ ) );
MUX2_X1 _21725_ ( .A(_01088_ ), .B(_01090_ ), .S(_01078_ ), .Z(\exu._io_out_bits_wdata_T_2 [16] ) );
MUX2_X1 _21726_ ( .A(\exu._GEN_0 [29] ), .B(\exu._GEN_0 [21] ), .S(\exu._io_out_bits_wdata_T_1 [3] ), .Z(_01091_ ) );
MUX2_X1 _21727_ ( .A(_01091_ ), .B(_12834_ ), .S(_01078_ ), .Z(\exu._io_out_bits_wdata_T_2 [29] ) );
MUX2_X1 _21728_ ( .A(\exu._GEN_0 [28] ), .B(\exu._GEN_0 [20] ), .S(_12823_ ), .Z(_01092_ ) );
MUX2_X1 _21729_ ( .A(_01092_ ), .B(_12835_ ), .S(_01078_ ), .Z(\exu._io_out_bits_wdata_T_2 [28] ) );
MUX2_X1 _21730_ ( .A(\exu._GEN_0 [27] ), .B(\exu._GEN_0 [19] ), .S(_12823_ ), .Z(_01093_ ) );
MUX2_X1 _21731_ ( .A(_01093_ ), .B(_12836_ ), .S(_01078_ ), .Z(\exu._io_out_bits_wdata_T_2 [27] ) );
MUX2_X1 _21732_ ( .A(\exu._GEN_0 [26] ), .B(\exu._GEN_0 [18] ), .S(_12823_ ), .Z(_01094_ ) );
MUX2_X1 _21733_ ( .A(_01094_ ), .B(_12837_ ), .S(_01078_ ), .Z(\exu._io_out_bits_wdata_T_2 [26] ) );
MUX2_X1 _21734_ ( .A(\exu._GEN_0 [25] ), .B(\exu._GEN_0 [17] ), .S(_12823_ ), .Z(_01095_ ) );
MUX2_X1 _21735_ ( .A(_01095_ ), .B(_12838_ ), .S(_01078_ ), .Z(\exu._io_out_bits_wdata_T_2 [25] ) );
MUX2_X1 _21736_ ( .A(\exu._GEN_0 [24] ), .B(\exu._GEN_0 [16] ), .S(_12823_ ), .Z(_01096_ ) );
MUX2_X1 _21737_ ( .A(_01096_ ), .B(_12839_ ), .S(_01078_ ), .Z(\exu._io_out_bits_wdata_T_2 [24] ) );
MUX2_X1 _21738_ ( .A(\exu._GEN_0 [23] ), .B(\exu._GEN_0 [15] ), .S(_12823_ ), .Z(_01097_ ) );
MUX2_X1 _21739_ ( .A(_01097_ ), .B(_12840_ ), .S(_01078_ ), .Z(\exu._io_out_bits_wdata_T_2 [23] ) );
MUX2_X1 _21740_ ( .A(\exu._GEN_0 [22] ), .B(\exu._GEN_0 [14] ), .S(_12823_ ), .Z(_01098_ ) );
MUX2_X1 _21741_ ( .A(_01098_ ), .B(_12842_ ), .S(_01078_ ), .Z(\exu._io_out_bits_wdata_T_2 [22] ) );
BUF_X2 _21742_ ( .A(_11125_ ), .Z(_01099_ ) );
BUF_X2 _21743_ ( .A(_01099_ ), .Z(_01100_ ) );
BUF_X2 _21744_ ( .A(_01100_ ), .Z(_01101_ ) );
BUF_X4 _21745_ ( .A(_01101_ ), .Z(_01102_ ) );
BUF_X2 _21746_ ( .A(_01102_ ), .Z(\idu.immI [4] ) );
NAND3_X1 _21747_ ( .A1(_10979_ ), .A2(fanout_net_8 ), .A3(\exu.auipc.io_rs1_data [31] ), .ZN(_01103_ ) );
NAND2_X1 _21748_ ( .A1(_10844_ ), .A2(\exu.csrrs.io_is ), .ZN(_01104_ ) );
NOR2_X1 _21749_ ( .A1(_01104_ ), .A2(\exu.csrrw.io_is ), .ZN(_01105_ ) );
BUF_X4 _21750_ ( .A(_01105_ ), .Z(_01106_ ) );
AOI21_X1 _21751_ ( .A(\exu.add.io_rs1_data [31] ), .B1(_01106_ ), .B2(\exu.csrrs.io_csr_rdata [31] ), .ZN(_01107_ ) );
NOR2_X2 _21752_ ( .A1(\exu.csrrs.io_is ), .A2(\exu.csrrw.io_is ), .ZN(_01108_ ) );
BUF_X4 _21753_ ( .A(_01108_ ), .Z(_01109_ ) );
NOR2_X1 _21754_ ( .A1(_01109_ ), .A2(fanout_net_26 ), .ZN(_01110_ ) );
NAND2_X1 _21755_ ( .A1(_01110_ ), .A2(_08989_ ), .ZN(_01111_ ) );
BUF_X4 _21756_ ( .A(_01111_ ), .Z(_01112_ ) );
OAI21_X1 _21757_ ( .A(_01103_ ), .B1(_01107_ ), .B2(_01112_ ), .ZN(\exu.io_out_bits_csr_wdata [31] ) );
NAND3_X1 _21758_ ( .A1(_10979_ ), .A2(fanout_net_8 ), .A3(\exu.auipc.io_rs1_data [30] ), .ZN(_01113_ ) );
AOI21_X1 _21759_ ( .A(\exu.add.io_rs1_data [30] ), .B1(_01106_ ), .B2(\exu.csrrs.io_csr_rdata [30] ), .ZN(_01114_ ) );
OAI21_X1 _21760_ ( .A(_01113_ ), .B1(_01114_ ), .B2(_01112_ ), .ZN(\exu.io_out_bits_csr_wdata [30] ) );
NAND3_X1 _21761_ ( .A1(_10979_ ), .A2(fanout_net_8 ), .A3(\exu.auipc.io_rs1_data [21] ), .ZN(_01115_ ) );
AOI21_X1 _21762_ ( .A(\exu.add.io_rs1_data [21] ), .B1(_01106_ ), .B2(\exu.csrrs.io_csr_rdata [21] ), .ZN(_01116_ ) );
OAI21_X1 _21763_ ( .A(_01115_ ), .B1(_01116_ ), .B2(_01112_ ), .ZN(\exu.io_out_bits_csr_wdata [21] ) );
BUF_X4 _21764_ ( .A(_10922_ ), .Z(_01117_ ) );
NAND3_X1 _21765_ ( .A1(_01117_ ), .A2(fanout_net_8 ), .A3(\exu.auipc.io_rs1_data [20] ), .ZN(_01118_ ) );
AOI21_X1 _21766_ ( .A(\exu.add.io_rs1_data [20] ), .B1(_01106_ ), .B2(\exu.csrrs.io_csr_rdata [20] ), .ZN(_01119_ ) );
OAI21_X1 _21767_ ( .A(_01118_ ), .B1(_01119_ ), .B2(_01112_ ), .ZN(\exu.io_out_bits_csr_wdata [20] ) );
NAND3_X1 _21768_ ( .A1(_01117_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [19] ), .ZN(_01120_ ) );
AOI21_X1 _21769_ ( .A(\exu.add.io_rs1_data [19] ), .B1(_01106_ ), .B2(\exu.csrrs.io_csr_rdata [19] ), .ZN(_01121_ ) );
OAI21_X1 _21770_ ( .A(_01120_ ), .B1(_01121_ ), .B2(_01112_ ), .ZN(\exu.io_out_bits_csr_wdata [19] ) );
BUF_X4 _21771_ ( .A(_01105_ ), .Z(_01122_ ) );
AOI21_X1 _21772_ ( .A(\exu.add.io_rs1_data [18] ), .B1(_01122_ ), .B2(\exu.csrrs.io_csr_rdata [18] ), .ZN(_01123_ ) );
BUF_X4 _21773_ ( .A(_01111_ ), .Z(_01124_ ) );
BUF_X4 _21774_ ( .A(_09456_ ), .Z(_01125_ ) );
OAI22_X1 _21775_ ( .A1(_01123_ ), .A2(_01124_ ), .B1(_09974_ ), .B2(_01125_ ), .ZN(\exu.io_out_bits_csr_wdata [18] ) );
NAND3_X1 _21776_ ( .A1(_01117_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [17] ), .ZN(_01126_ ) );
AOI21_X1 _21777_ ( .A(\exu.add.io_rs1_data [17] ), .B1(_01106_ ), .B2(\exu.csrrs.io_csr_rdata [17] ), .ZN(_01127_ ) );
OAI21_X1 _21778_ ( .A(_01126_ ), .B1(_01127_ ), .B2(_01112_ ), .ZN(\exu.io_out_bits_csr_wdata [17] ) );
NAND3_X1 _21779_ ( .A1(_01117_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [16] ), .ZN(_01128_ ) );
AOI21_X1 _21780_ ( .A(\exu.add.io_rs1_data [16] ), .B1(_01106_ ), .B2(\exu.csrrs.io_csr_rdata [16] ), .ZN(_01129_ ) );
OAI21_X1 _21781_ ( .A(_01128_ ), .B1(_01129_ ), .B2(_01112_ ), .ZN(\exu.io_out_bits_csr_wdata [16] ) );
NAND3_X1 _21782_ ( .A1(_01117_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [15] ), .ZN(_01130_ ) );
AOI21_X1 _21783_ ( .A(\exu.add.io_rs1_data [15] ), .B1(_01106_ ), .B2(\exu.csrrs.io_csr_rdata [15] ), .ZN(_01131_ ) );
OAI21_X1 _21784_ ( .A(_01130_ ), .B1(_01131_ ), .B2(_01112_ ), .ZN(\exu.io_out_bits_csr_wdata [15] ) );
AOI21_X1 _21785_ ( .A(\exu.add.io_rs1_data [14] ), .B1(_01122_ ), .B2(\exu.csrrs.io_csr_rdata [14] ), .ZN(_01132_ ) );
OAI22_X1 _21786_ ( .A1(_01132_ ), .A2(_01124_ ), .B1(_10120_ ), .B2(_01125_ ), .ZN(\exu.io_out_bits_csr_wdata [14] ) );
AOI21_X1 _21787_ ( .A(\exu.add.io_rs1_data [13] ), .B1(_01122_ ), .B2(\exu.csrrs.io_csr_rdata [13] ), .ZN(_01133_ ) );
OAI22_X1 _21788_ ( .A1(_01133_ ), .A2(_01124_ ), .B1(_08648_ ), .B2(_01125_ ), .ZN(\exu.io_out_bits_csr_wdata [13] ) );
AOI21_X1 _21789_ ( .A(\exu.add.io_rs1_data [12] ), .B1(_01122_ ), .B2(\exu.csrrs.io_csr_rdata [12] ), .ZN(_01134_ ) );
OAI22_X1 _21790_ ( .A1(_01134_ ), .A2(_01124_ ), .B1(_08800_ ), .B2(_01125_ ), .ZN(\exu.io_out_bits_csr_wdata [12] ) );
NAND3_X1 _21791_ ( .A1(_01117_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [29] ), .ZN(_01135_ ) );
AOI21_X1 _21792_ ( .A(\exu.add.io_rs1_data [29] ), .B1(_01106_ ), .B2(\exu.csrrs.io_csr_rdata [29] ), .ZN(_01136_ ) );
OAI21_X1 _21793_ ( .A(_01135_ ), .B1(_01136_ ), .B2(_01112_ ), .ZN(\exu.io_out_bits_csr_wdata [29] ) );
NAND3_X1 _21794_ ( .A1(_01117_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [11] ), .ZN(_01137_ ) );
AOI21_X1 _21795_ ( .A(\exu.add.io_rs1_data [11] ), .B1(_01106_ ), .B2(\exu.csrrs.io_csr_rdata [11] ), .ZN(_01138_ ) );
OAI21_X1 _21796_ ( .A(_01137_ ), .B1(_01138_ ), .B2(_01112_ ), .ZN(\exu.io_out_bits_csr_wdata [11] ) );
AOI21_X1 _21797_ ( .A(\exu.add.io_rs1_data [10] ), .B1(_01122_ ), .B2(\exu.csrrs.io_csr_rdata [10] ), .ZN(_01139_ ) );
OAI22_X1 _21798_ ( .A1(_01139_ ), .A2(_01124_ ), .B1(_10211_ ), .B2(_01125_ ), .ZN(\exu.io_out_bits_csr_wdata [10] ) );
NAND3_X1 _21799_ ( .A1(_01117_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [9] ), .ZN(_01140_ ) );
BUF_X4 _21800_ ( .A(_01105_ ), .Z(_01141_ ) );
AOI21_X1 _21801_ ( .A(\exu.add.io_rs1_data [9] ), .B1(_01141_ ), .B2(\exu.csrrs.io_csr_rdata [9] ), .ZN(_01142_ ) );
BUF_X4 _21802_ ( .A(_01111_ ), .Z(_01143_ ) );
OAI21_X1 _21803_ ( .A(_01140_ ), .B1(_01142_ ), .B2(_01143_ ), .ZN(\exu.io_out_bits_csr_wdata [9] ) );
NAND3_X1 _21804_ ( .A1(_01117_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [8] ), .ZN(_01144_ ) );
AOI21_X1 _21805_ ( .A(\exu.add.io_rs1_data [8] ), .B1(_01141_ ), .B2(\exu.csrrs.io_csr_rdata [8] ), .ZN(_01145_ ) );
OAI21_X1 _21806_ ( .A(_01144_ ), .B1(_01145_ ), .B2(_01143_ ), .ZN(\exu.io_out_bits_csr_wdata [8] ) );
NAND3_X1 _21807_ ( .A1(_01117_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [7] ), .ZN(_01146_ ) );
AOI21_X1 _21808_ ( .A(\exu.add.io_rs1_data [7] ), .B1(_01141_ ), .B2(\exu.csrrs.io_csr_rdata [7] ), .ZN(_01147_ ) );
OAI21_X1 _21809_ ( .A(_01146_ ), .B1(_01147_ ), .B2(_01143_ ), .ZN(\exu.io_out_bits_csr_wdata [7] ) );
NAND3_X1 _21810_ ( .A1(_11892_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [6] ), .ZN(_01148_ ) );
AOI21_X1 _21811_ ( .A(\exu.add.io_rs1_data [6] ), .B1(_01141_ ), .B2(\exu.csrrs.io_csr_rdata [6] ), .ZN(_01149_ ) );
OAI21_X1 _21812_ ( .A(_01148_ ), .B1(_01149_ ), .B2(_01143_ ), .ZN(\exu.io_out_bits_csr_wdata [6] ) );
AOI21_X1 _21813_ ( .A(\exu.add.io_rs1_data [5] ), .B1(_01122_ ), .B2(\exu.csrrs.io_csr_rdata [5] ), .ZN(_01150_ ) );
OAI22_X1 _21814_ ( .A1(_01150_ ), .A2(_01124_ ), .B1(_08608_ ), .B2(_01125_ ), .ZN(\exu.io_out_bits_csr_wdata [5] ) );
NAND3_X1 _21815_ ( .A1(_11892_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [4] ), .ZN(_01151_ ) );
AOI21_X1 _21816_ ( .A(\exu.add.io_rs1_data [4] ), .B1(_01141_ ), .B2(\exu.csrrs.io_csr_rdata [4] ), .ZN(_01152_ ) );
OAI21_X1 _21817_ ( .A(_01151_ ), .B1(_01152_ ), .B2(_01143_ ), .ZN(\exu.io_out_bits_csr_wdata [4] ) );
AOI21_X1 _21818_ ( .A(\exu.add.io_rs1_data [3] ), .B1(_01122_ ), .B2(\exu.csrrs.io_csr_rdata [3] ), .ZN(_01153_ ) );
OAI22_X1 _21819_ ( .A1(_01153_ ), .A2(_01124_ ), .B1(_09196_ ), .B2(_01125_ ), .ZN(\exu.io_out_bits_csr_wdata [3] ) );
AOI21_X1 _21820_ ( .A(\exu.add.io_rs1_data [2] ), .B1(_01122_ ), .B2(\exu.csrrs.io_csr_rdata [2] ), .ZN(_01154_ ) );
OAI22_X1 _21821_ ( .A1(_01154_ ), .A2(_01124_ ), .B1(_09197_ ), .B2(_01125_ ), .ZN(\exu.io_out_bits_csr_wdata [2] ) );
NAND3_X1 _21822_ ( .A1(_11892_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [28] ), .ZN(_01155_ ) );
AOI21_X1 _21823_ ( .A(\exu.add.io_rs1_data [28] ), .B1(_01141_ ), .B2(\exu.csrrs.io_csr_rdata [28] ), .ZN(_01156_ ) );
OAI21_X1 _21824_ ( .A(_01155_ ), .B1(_01156_ ), .B2(_01143_ ), .ZN(\exu.io_out_bits_csr_wdata [28] ) );
AOI21_X1 _21825_ ( .A(\exu.add.io_rs1_data [1] ), .B1(_01122_ ), .B2(\exu.csrrs.io_csr_rdata [1] ), .ZN(_01157_ ) );
OAI22_X1 _21826_ ( .A1(_01157_ ), .A2(_01124_ ), .B1(_08591_ ), .B2(_01125_ ), .ZN(\exu.io_out_bits_csr_wdata [1] ) );
AOI21_X1 _21827_ ( .A(\exu.add.io_rs1_data [0] ), .B1(_01122_ ), .B2(\exu.csrrs.io_csr_rdata [0] ), .ZN(_01158_ ) );
OAI22_X1 _21828_ ( .A1(_01158_ ), .A2(_01124_ ), .B1(_11377_ ), .B2(_01125_ ), .ZN(\exu.io_out_bits_csr_wdata [0] ) );
NAND3_X1 _21829_ ( .A1(_11892_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [27] ), .ZN(_01159_ ) );
AOI21_X1 _21830_ ( .A(\exu.add.io_rs1_data [27] ), .B1(_01141_ ), .B2(\exu.csrrs.io_csr_rdata [27] ), .ZN(_01160_ ) );
OAI21_X1 _21831_ ( .A(_01159_ ), .B1(_01160_ ), .B2(_01143_ ), .ZN(\exu.io_out_bits_csr_wdata [27] ) );
NAND3_X1 _21832_ ( .A1(_11892_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [26] ), .ZN(_01161_ ) );
AOI21_X1 _21833_ ( .A(\exu.add.io_rs1_data [26] ), .B1(_01141_ ), .B2(\exu.csrrs.io_csr_rdata [26] ), .ZN(_01162_ ) );
OAI21_X1 _21834_ ( .A(_01161_ ), .B1(_01162_ ), .B2(_01143_ ), .ZN(\exu.io_out_bits_csr_wdata [26] ) );
NAND3_X1 _21835_ ( .A1(_11892_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [25] ), .ZN(_01163_ ) );
AOI21_X1 _21836_ ( .A(\exu.add.io_rs1_data [25] ), .B1(_01141_ ), .B2(\exu.csrrs.io_csr_rdata [25] ), .ZN(_01164_ ) );
OAI21_X1 _21837_ ( .A(_01163_ ), .B1(_01164_ ), .B2(_01143_ ), .ZN(\exu.io_out_bits_csr_wdata [25] ) );
NAND3_X1 _21838_ ( .A1(_11892_ ), .A2(\exu.ecall.io_is ), .A3(\exu.auipc.io_rs1_data [24] ), .ZN(_01165_ ) );
AOI21_X1 _21839_ ( .A(\exu.add.io_rs1_data [24] ), .B1(_01141_ ), .B2(\exu.csrrs.io_csr_rdata [24] ), .ZN(_01166_ ) );
OAI21_X1 _21840_ ( .A(_01165_ ), .B1(_01166_ ), .B2(_01143_ ), .ZN(\exu.io_out_bits_csr_wdata [24] ) );
AOI21_X1 _21841_ ( .A(\exu.add.io_rs1_data [23] ), .B1(_01105_ ), .B2(\exu.csrrs.io_csr_rdata [23] ), .ZN(_01167_ ) );
OAI22_X1 _21842_ ( .A1(_01167_ ), .A2(_01111_ ), .B1(_08668_ ), .B2(_09456_ ), .ZN(\exu.io_out_bits_csr_wdata [23] ) );
AOI21_X1 _21843_ ( .A(\exu.add.io_rs1_data [22] ), .B1(_01105_ ), .B2(\exu.csrrs.io_csr_rdata [22] ), .ZN(_01168_ ) );
OAI22_X1 _21844_ ( .A1(_01168_ ), .A2(_01111_ ), .B1(_09528_ ), .B2(_09456_ ), .ZN(\exu.io_out_bits_csr_wdata [22] ) );
INV_X1 _21845_ ( .A(\exu.io_in_bits_sltiu ), .ZN(_01169_ ) );
NAND2_X1 _21846_ ( .A1(_01169_ ), .A2(exu_io_in_bits_r_slti_$_NOT__A_Y ), .ZN(_01170_ ) );
NOR2_X1 _21847_ ( .A1(_01170_ ), .A2(\exu.addi.io_is ), .ZN(_01171_ ) );
INV_X1 _21848_ ( .A(_01171_ ), .ZN(_01172_ ) );
BUF_X4 _21849_ ( .A(_01172_ ), .Z(_01173_ ) );
INV_X1 _21850_ ( .A(\exu.io_in_bits_xori ), .ZN(_01174_ ) );
BUF_X4 _21851_ ( .A(_01174_ ), .Z(_01175_ ) );
INV_X2 _21852_ ( .A(fanout_net_5 ), .ZN(_01176_ ) );
INV_X1 _21853_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B ), .ZN(_01177_ ) );
INV_X1 _21854_ ( .A(\exu.io_in_bits_shamt [5] ), .ZN(_01178_ ) );
AND4_X1 _21855_ ( .A1(_10699_ ), .A2(_01177_ ), .A3(_01178_ ), .A4(\exu.io_in_bits_srai ), .ZN(_01179_ ) );
INV_X2 _21856_ ( .A(\exu.io_in_bits_srai ), .ZN(_01180_ ) );
BUF_X4 _21857_ ( .A(_01180_ ), .Z(_01181_ ) );
BUF_X4 _21858_ ( .A(_01181_ ), .Z(_01182_ ) );
OAI21_X1 _21859_ ( .A(_01176_ ), .B1(_01179_ ), .B2(_01182_ ), .ZN(_01183_ ) );
INV_X1 _21860_ ( .A(\exu.io_in_bits_ori ), .ZN(_01184_ ) );
NOR2_X1 _21861_ ( .A1(_01184_ ), .A2(fanout_net_26 ), .ZN(_01185_ ) );
BUF_X4 _21862_ ( .A(_01185_ ), .Z(_01186_ ) );
OAI21_X1 _21863_ ( .A(_01186_ ), .B1(\exu.add.io_rs1_data [31] ), .B2(\exu.addi.io_imm [31] ), .ZN(_01187_ ) );
INV_X1 _21864_ ( .A(\exu.io_in_bits_srli ), .ZN(_01188_ ) );
NAND2_X1 _21865_ ( .A1(_01188_ ), .A2(_01089_ ), .ZN(_01189_ ) );
BUF_X2 _21866_ ( .A(_01189_ ), .Z(_01190_ ) );
INV_X1 _21867_ ( .A(\exu.io_in_bits_shamt [0] ), .ZN(_01191_ ) );
NAND2_X1 _21868_ ( .A1(_01191_ ), .A2(\exu.io_in_bits_srli ), .ZN(_01192_ ) );
BUF_X2 _21869_ ( .A(_01192_ ), .Z(_01193_ ) );
AOI21_X1 _21870_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B ), .B1(_01190_ ), .B2(_01193_ ), .ZN(_01194_ ) );
NAND2_X1 _21871_ ( .A1(_01188_ ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_14_B_$_ANDNOT__Y_B ), .ZN(_01195_ ) );
NAND2_X1 _21872_ ( .A1(\exu.io_in_bits_srli ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__A_B ), .ZN(_01196_ ) );
NAND2_X2 _21873_ ( .A1(_01195_ ), .A2(_01196_ ), .ZN(_01197_ ) );
NAND2_X1 _21874_ ( .A1(_01188_ ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_13_B_$_ANDNOT__Y_B ), .ZN(_01198_ ) );
NAND2_X1 _21875_ ( .A1(\exu.io_in_bits_srli ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__A_B ), .ZN(_01199_ ) );
NAND2_X2 _21876_ ( .A1(_01198_ ), .A2(_01199_ ), .ZN(_01200_ ) );
AND3_X1 _21877_ ( .A1(_01194_ ), .A2(_01197_ ), .A3(_01200_ ), .ZN(_01201_ ) );
NAND2_X1 _21878_ ( .A1(_01188_ ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_12_B_$_ANDNOT__Y_B ), .ZN(_01202_ ) );
NAND2_X1 _21879_ ( .A1(\exu.io_in_bits_srli ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__A_B ), .ZN(_01203_ ) );
NAND2_X1 _21880_ ( .A1(_01202_ ), .A2(_01203_ ), .ZN(_01204_ ) );
BUF_X2 _21881_ ( .A(_01204_ ), .Z(_01205_ ) );
BUF_X2 _21882_ ( .A(_01205_ ), .Z(_01206_ ) );
BUF_X2 _21883_ ( .A(_01206_ ), .Z(_01207_ ) );
NAND2_X1 _21884_ ( .A1(_01188_ ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_11_B_$_ANDNOT__Y_B ), .ZN(_01208_ ) );
NAND2_X1 _21885_ ( .A1(\exu.io_in_bits_srli ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__A_B ), .ZN(_01209_ ) );
NAND2_X1 _21886_ ( .A1(_01208_ ), .A2(_01209_ ), .ZN(_01210_ ) );
BUF_X2 _21887_ ( .A(_01210_ ), .Z(_01211_ ) );
CLKBUF_X2 _21888_ ( .A(_01211_ ), .Z(_01212_ ) );
BUF_X2 _21889_ ( .A(_01212_ ), .Z(_01213_ ) );
BUF_X4 _21890_ ( .A(_01188_ ), .Z(_01214_ ) );
NOR2_X1 _21891_ ( .A1(_01214_ ), .A2(fanout_net_26 ), .ZN(_01215_ ) );
AND2_X1 _21892_ ( .A1(_01215_ ), .A2(_01178_ ), .ZN(_01216_ ) );
BUF_X2 _21893_ ( .A(_01216_ ), .Z(_01217_ ) );
NAND4_X1 _21894_ ( .A1(_01201_ ), .A2(_01207_ ), .A3(_01213_ ), .A4(_01217_ ), .ZN(_01218_ ) );
INV_X1 _21895_ ( .A(\exu.io_in_bits_slli ), .ZN(_01219_ ) );
NAND2_X1 _21896_ ( .A1(_01219_ ), .A2(_01089_ ), .ZN(_01220_ ) );
BUF_X2 _21897_ ( .A(_01220_ ), .Z(_01221_ ) );
NAND2_X1 _21898_ ( .A1(_01191_ ), .A2(\exu.io_in_bits_slli ), .ZN(_01222_ ) );
BUF_X2 _21899_ ( .A(_01222_ ), .Z(_01223_ ) );
AND3_X1 _21900_ ( .A1(_01221_ ), .A2(_01223_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01224_ ) );
INV_X1 _21901_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01225_ ) );
BUF_X2 _21902_ ( .A(_01220_ ), .Z(_01226_ ) );
BUF_X2 _21903_ ( .A(_01222_ ), .Z(_01227_ ) );
AOI21_X1 _21904_ ( .A(_01225_ ), .B1(_01226_ ), .B2(_01227_ ), .ZN(_01228_ ) );
OR2_X1 _21905_ ( .A1(_01224_ ), .A2(_01228_ ), .ZN(_01229_ ) );
AND2_X2 _21906_ ( .A1(_01220_ ), .A2(_01222_ ), .ZN(_01230_ ) );
MUX2_X1 _21907_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .S(_01230_ ), .Z(_01231_ ) );
NAND2_X1 _21908_ ( .A1(_01219_ ), .A2(\exu._GEN_0 [1] ), .ZN(_01232_ ) );
NAND2_X1 _21909_ ( .A1(\exu.io_in_bits_slli ), .A2(\exu.io_in_bits_shamt [1] ), .ZN(_01233_ ) );
NAND2_X1 _21910_ ( .A1(_01232_ ), .A2(_01233_ ), .ZN(_01234_ ) );
BUF_X4 _21911_ ( .A(_01234_ ), .Z(_01235_ ) );
MUX2_X1 _21912_ ( .A(_01229_ ), .B(_01231_ ), .S(_01235_ ), .Z(_01236_ ) );
NAND2_X1 _21913_ ( .A1(_01219_ ), .A2(\exu._GEN_0 [2] ), .ZN(_01237_ ) );
NAND2_X1 _21914_ ( .A1(\exu.io_in_bits_slli ), .A2(\exu.io_in_bits_shamt [2] ), .ZN(_01238_ ) );
NAND2_X1 _21915_ ( .A1(_01237_ ), .A2(_01238_ ), .ZN(_01239_ ) );
BUF_X4 _21916_ ( .A(_01239_ ), .Z(_01240_ ) );
BUF_X2 _21917_ ( .A(_01240_ ), .Z(_01241_ ) );
NAND2_X1 _21918_ ( .A1(_01236_ ), .A2(_01241_ ), .ZN(_01242_ ) );
NAND2_X1 _21919_ ( .A1(_01219_ ), .A2(\exu._GEN_0 [3] ), .ZN(_01243_ ) );
NAND2_X1 _21920_ ( .A1(\exu.io_in_bits_slli ), .A2(\exu.io_in_bits_shamt [3] ), .ZN(_01244_ ) );
NAND2_X1 _21921_ ( .A1(_01243_ ), .A2(_01244_ ), .ZN(_01245_ ) );
BUF_X4 _21922_ ( .A(_01245_ ), .Z(_01246_ ) );
AND3_X1 _21923_ ( .A1(_01220_ ), .A2(_01222_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01247_ ) );
INV_X1 _21924_ ( .A(_01234_ ), .ZN(_01248_ ) );
INV_X1 _21925_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01249_ ) );
AOI21_X1 _21926_ ( .A(_01249_ ), .B1(_01220_ ), .B2(_01222_ ), .ZN(_01250_ ) );
OR3_X1 _21927_ ( .A1(_01247_ ), .A2(_01248_ ), .A3(_01250_ ), .ZN(_01251_ ) );
INV_X2 _21928_ ( .A(_01239_ ), .ZN(_01252_ ) );
BUF_X2 _21929_ ( .A(_01235_ ), .Z(_01253_ ) );
BUF_X2 _21930_ ( .A(_01253_ ), .Z(_01254_ ) );
INV_X1 _21931_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01255_ ) );
AND3_X1 _21932_ ( .A1(_01220_ ), .A2(_01223_ ), .A3(_01255_ ), .ZN(_01256_ ) );
AOI21_X1 _21933_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01221_ ), .B2(_01223_ ), .ZN(_01257_ ) );
NOR2_X1 _21934_ ( .A1(_01256_ ), .A2(_01257_ ), .ZN(_01258_ ) );
OAI211_X1 _21935_ ( .A(_01251_ ), .B(_01252_ ), .C1(_01254_ ), .C2(_01258_ ), .ZN(_01259_ ) );
NAND3_X1 _21936_ ( .A1(_01242_ ), .A2(_01246_ ), .A3(_01259_ ), .ZN(_01260_ ) );
INV_X1 _21937_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01261_ ) );
OR2_X1 _21938_ ( .A1(_01230_ ), .A2(_01261_ ), .ZN(_01262_ ) );
INV_X1 _21939_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01263_ ) );
INV_X1 _21940_ ( .A(_01230_ ), .ZN(_01264_ ) );
OAI211_X1 _21941_ ( .A(_01262_ ), .B(_01248_ ), .C1(_01263_ ), .C2(_01264_ ), .ZN(_01265_ ) );
NAND3_X1 _21942_ ( .A1(_01226_ ), .A2(_01227_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01266_ ) );
INV_X1 _21943_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01267_ ) );
OAI211_X1 _21944_ ( .A(_01234_ ), .B(_01266_ ), .C1(_01230_ ), .C2(_01267_ ), .ZN(_01268_ ) );
NAND3_X1 _21945_ ( .A1(_01265_ ), .A2(_01241_ ), .A3(_01268_ ), .ZN(_01269_ ) );
INV_X1 _21946_ ( .A(_01245_ ), .ZN(_01270_ ) );
BUF_X4 _21947_ ( .A(_01270_ ), .Z(_01271_ ) );
NAND3_X1 _21948_ ( .A1(_01226_ ), .A2(_01227_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01272_ ) );
BUF_X4 _21949_ ( .A(_01230_ ), .Z(_01273_ ) );
INV_X1 _21950_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01274_ ) );
OAI211_X1 _21951_ ( .A(_01234_ ), .B(_01272_ ), .C1(_01273_ ), .C2(_01274_ ), .ZN(_01275_ ) );
NAND3_X1 _21952_ ( .A1(_01226_ ), .A2(_01227_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01276_ ) );
INV_X1 _21953_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01277_ ) );
OAI211_X1 _21954_ ( .A(_01248_ ), .B(_01276_ ), .C1(_01230_ ), .C2(_01277_ ), .ZN(_01278_ ) );
BUF_X2 _21955_ ( .A(_01252_ ), .Z(_01279_ ) );
NAND3_X1 _21956_ ( .A1(_01275_ ), .A2(_01278_ ), .A3(_01279_ ), .ZN(_01280_ ) );
NAND3_X1 _21957_ ( .A1(_01269_ ), .A2(_01271_ ), .A3(_01280_ ), .ZN(_01281_ ) );
NAND2_X1 _21958_ ( .A1(_01260_ ), .A2(_01281_ ), .ZN(_01282_ ) );
INV_X1 _21959_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01283_ ) );
AND3_X1 _21960_ ( .A1(_01226_ ), .A2(_01227_ ), .A3(_01283_ ), .ZN(_01284_ ) );
BUF_X2 _21961_ ( .A(_01221_ ), .Z(_01285_ ) );
BUF_X2 _21962_ ( .A(_01222_ ), .Z(_01286_ ) );
AOI21_X1 _21963_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01285_ ), .B2(_01286_ ), .ZN(_01287_ ) );
NOR2_X1 _21964_ ( .A1(_01284_ ), .A2(_01287_ ), .ZN(_01288_ ) );
NAND2_X1 _21965_ ( .A1(_01288_ ), .A2(_01253_ ), .ZN(_01289_ ) );
BUF_X4 _21966_ ( .A(_01248_ ), .Z(_01290_ ) );
BUF_X4 _21967_ ( .A(_01290_ ), .Z(_01291_ ) );
AND3_X1 _21968_ ( .A1(_01220_ ), .A2(_01222_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01292_ ) );
INV_X1 _21969_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01293_ ) );
AOI21_X1 _21970_ ( .A(_01293_ ), .B1(_01221_ ), .B2(_01223_ ), .ZN(_01294_ ) );
OAI21_X1 _21971_ ( .A(_01291_ ), .B1(_01292_ ), .B2(_01294_ ), .ZN(_01295_ ) );
AND3_X1 _21972_ ( .A1(_01289_ ), .A2(_01240_ ), .A3(_01295_ ), .ZN(_01296_ ) );
BUF_X4 _21973_ ( .A(_01273_ ), .Z(_01297_ ) );
MUX2_X1 _21974_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B ), .B(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_01297_ ), .Z(_01298_ ) );
BUF_X4 _21975_ ( .A(_01291_ ), .Z(_01299_ ) );
AND2_X1 _21976_ ( .A1(_01298_ ), .A2(_01299_ ), .ZN(_01300_ ) );
INV_X1 _21977_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01301_ ) );
AND3_X1 _21978_ ( .A1(_01221_ ), .A2(_01223_ ), .A3(_01301_ ), .ZN(_01302_ ) );
AOI21_X1 _21979_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01226_ ), .B2(_01227_ ), .ZN(_01303_ ) );
NOR2_X1 _21980_ ( .A1(_01302_ ), .A2(_01303_ ), .ZN(_01304_ ) );
AOI21_X1 _21981_ ( .A(_01300_ ), .B1(_01254_ ), .B2(_01304_ ), .ZN(_01305_ ) );
BUF_X4 _21982_ ( .A(_01252_ ), .Z(_01306_ ) );
AOI211_X1 _21983_ ( .A(_01246_ ), .B(_01296_ ), .C1(_01305_ ), .C2(_01306_ ), .ZN(_01307_ ) );
BUF_X4 _21984_ ( .A(_01246_ ), .Z(_01308_ ) );
BUF_X2 _21985_ ( .A(_01226_ ), .Z(_01309_ ) );
BUF_X2 _21986_ ( .A(_01227_ ), .Z(_01310_ ) );
NAND3_X1 _21987_ ( .A1(_01309_ ), .A2(_01310_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01311_ ) );
INV_X1 _21988_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01312_ ) );
OAI211_X1 _21989_ ( .A(_01254_ ), .B(_01311_ ), .C1(_01297_ ), .C2(_01312_ ), .ZN(_01313_ ) );
AND3_X1 _21990_ ( .A1(_01226_ ), .A2(_01227_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01314_ ) );
INV_X1 _21991_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01315_ ) );
AOI21_X1 _21992_ ( .A(_01315_ ), .B1(_01285_ ), .B2(_01286_ ), .ZN(_01316_ ) );
OR2_X1 _21993_ ( .A1(_01314_ ), .A2(_01316_ ), .ZN(_01317_ ) );
OAI211_X1 _21994_ ( .A(_01279_ ), .B(_01313_ ), .C1(_01317_ ), .C2(_01254_ ), .ZN(_01318_ ) );
NAND3_X1 _21995_ ( .A1(_01226_ ), .A2(_01227_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01319_ ) );
INV_X1 _21996_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01320_ ) );
OAI211_X1 _21997_ ( .A(_01234_ ), .B(_01319_ ), .C1(_01273_ ), .C2(_01320_ ), .ZN(_01321_ ) );
NAND3_X1 _21998_ ( .A1(_01226_ ), .A2(_01227_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01322_ ) );
INV_X1 _21999_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01323_ ) );
OAI211_X1 _22000_ ( .A(_01290_ ), .B(_01322_ ), .C1(_01273_ ), .C2(_01323_ ), .ZN(_01324_ ) );
BUF_X2 _22001_ ( .A(_01240_ ), .Z(_01325_ ) );
NAND3_X1 _22002_ ( .A1(_01321_ ), .A2(_01324_ ), .A3(_01325_ ), .ZN(_01326_ ) );
NAND2_X1 _22003_ ( .A1(_01318_ ), .A2(_01326_ ), .ZN(_01327_ ) );
AOI21_X1 _22004_ ( .A(_01307_ ), .B1(_01308_ ), .B2(_01327_ ), .ZN(_01328_ ) );
NAND2_X1 _22005_ ( .A1(_01219_ ), .A2(\exu._GEN_0 [4] ), .ZN(_01329_ ) );
NAND2_X1 _22006_ ( .A1(\exu.io_in_bits_slli ), .A2(\exu.io_in_bits_shamt [4] ), .ZN(_01330_ ) );
NAND2_X1 _22007_ ( .A1(_01329_ ), .A2(_01330_ ), .ZN(_01331_ ) );
INV_X1 _22008_ ( .A(_01331_ ), .ZN(_01332_ ) );
BUF_X2 _22009_ ( .A(_01332_ ), .Z(_01333_ ) );
MUX2_X1 _22010_ ( .A(_01282_ ), .B(_01328_ ), .S(_01333_ ), .Z(_01334_ ) );
NOR2_X1 _22011_ ( .A1(_01219_ ), .A2(fanout_net_26 ), .ZN(_01335_ ) );
AND2_X1 _22012_ ( .A1(_01335_ ), .A2(_01178_ ), .ZN(_01336_ ) );
BUF_X2 _22013_ ( .A(_01336_ ), .Z(_01337_ ) );
BUF_X4 _22014_ ( .A(_01337_ ), .Z(_01338_ ) );
NAND2_X1 _22015_ ( .A1(_01334_ ), .A2(_01338_ ), .ZN(_01339_ ) );
BUF_X4 _22016_ ( .A(_09657_ ), .Z(_01340_ ) );
BUF_X4 _22017_ ( .A(_01340_ ), .Z(_01341_ ) );
BUF_X2 _22018_ ( .A(_09999_ ), .Z(_01342_ ) );
INV_X1 _22019_ ( .A(_08762_ ), .ZN(_01343_ ) );
INV_X1 _22020_ ( .A(_08765_ ), .ZN(_01344_ ) );
INV_X1 _22021_ ( .A(_08768_ ), .ZN(_01345_ ) );
INV_X1 _22022_ ( .A(_08769_ ), .ZN(_01346_ ) );
NAND2_X1 _22023_ ( .A1(_08717_ ), .A2(_08718_ ), .ZN(_01347_ ) );
INV_X1 _22024_ ( .A(_08720_ ), .ZN(_01348_ ) );
INV_X1 _22025_ ( .A(_08723_ ), .ZN(_01349_ ) );
NOR3_X1 _22026_ ( .A1(_01347_ ), .A2(_01348_ ), .A3(_01349_ ), .ZN(_01350_ ) );
AND2_X1 _22027_ ( .A1(_08705_ ), .A2(_08708_ ), .ZN(_01351_ ) );
AND3_X1 _22028_ ( .A1(_01351_ ), .A2(_08712_ ), .A3(_08714_ ), .ZN(_01352_ ) );
INV_X1 _22029_ ( .A(_08732_ ), .ZN(_01353_ ) );
AND2_X1 _22030_ ( .A1(\exu.add.io_rs1_data [0] ), .A2(\exu._GEN_0 [0] ), .ZN(_01354_ ) );
AND2_X1 _22031_ ( .A1(_08778_ ), .A2(_01354_ ), .ZN(_01355_ ) );
AND2_X1 _22032_ ( .A1(\exu.add.io_rs1_data [1] ), .A2(\exu._GEN_0 [1] ), .ZN(_01356_ ) );
OAI21_X1 _22033_ ( .A(_08779_ ), .B1(_01355_ ), .B2(_01356_ ), .ZN(_01357_ ) );
AND2_X1 _22034_ ( .A1(\exu.add.io_rs1_data [2] ), .A2(\exu._GEN_0 [2] ), .ZN(_01358_ ) );
INV_X1 _22035_ ( .A(_01358_ ), .ZN(_01359_ ) );
AOI21_X1 _22036_ ( .A(_08739_ ), .B1(_01357_ ), .B2(_01359_ ), .ZN(_01360_ ) );
INV_X1 _22037_ ( .A(_01360_ ), .ZN(_01361_ ) );
AND2_X1 _22038_ ( .A1(\exu.add.io_rs1_data [3] ), .A2(\exu._GEN_0 [3] ), .ZN(_01362_ ) );
INV_X1 _22039_ ( .A(_01362_ ), .ZN(_01363_ ) );
AOI21_X1 _22040_ ( .A(_01353_ ), .B1(_01361_ ), .B2(_01363_ ), .ZN(_01364_ ) );
AND2_X1 _22041_ ( .A1(\exu.add.io_rs1_data [4] ), .A2(\exu._GEN_0 [4] ), .ZN(_01365_ ) );
NOR2_X1 _22042_ ( .A1(_01364_ ), .A2(_01365_ ), .ZN(_01366_ ) );
NOR2_X1 _22043_ ( .A1(_01366_ ), .A2(_08734_ ), .ZN(_01367_ ) );
AOI21_X1 _22044_ ( .A(_01367_ ), .B1(\exu.add.io_rs1_data [5] ), .B2(\exu._GEN_0 [5] ), .ZN(_01368_ ) );
INV_X1 _22045_ ( .A(_08727_ ), .ZN(_01369_ ) );
NOR2_X1 _22046_ ( .A1(_01368_ ), .A2(_01369_ ), .ZN(_01370_ ) );
AND2_X1 _22047_ ( .A1(\exu.add.io_rs1_data [6] ), .A2(\exu._GEN_0 [6] ), .ZN(_01371_ ) );
NOR2_X1 _22048_ ( .A1(_01370_ ), .A2(_01371_ ), .ZN(_01372_ ) );
NOR2_X1 _22049_ ( .A1(_01372_ ), .A2(_08729_ ), .ZN(_01373_ ) );
OAI211_X1 _22050_ ( .A(_01350_ ), .B(_01352_ ), .C1(_01373_ ), .C2(_08728_ ), .ZN(_01374_ ) );
INV_X1 _22051_ ( .A(_08707_ ), .ZN(_01375_ ) );
AND2_X1 _22052_ ( .A1(\exu.add.io_rs1_data [10] ), .A2(\exu._GEN_0 [10] ), .ZN(_01376_ ) );
AOI21_X1 _22053_ ( .A(_08706_ ), .B1(_01375_ ), .B2(_01376_ ), .ZN(_01377_ ) );
INV_X1 _22054_ ( .A(_01351_ ), .ZN(_01378_ ) );
INV_X1 _22055_ ( .A(_08711_ ), .ZN(_01379_ ) );
AND2_X1 _22056_ ( .A1(\exu.add.io_rs1_data [8] ), .A2(\exu._GEN_0 [8] ), .ZN(_01380_ ) );
AOI21_X1 _22057_ ( .A(_08710_ ), .B1(_01379_ ), .B2(_01380_ ), .ZN(_01381_ ) );
OAI21_X1 _22058_ ( .A(_01377_ ), .B1(_01378_ ), .B2(_01381_ ), .ZN(_01382_ ) );
AND2_X1 _22059_ ( .A1(_01382_ ), .A2(_01350_ ), .ZN(_01383_ ) );
AND2_X1 _22060_ ( .A1(\exu.add.io_rs1_data [15] ), .A2(\exu._GEN_0 [15] ), .ZN(_01384_ ) );
AND2_X1 _22061_ ( .A1(\exu.add.io_rs1_data [12] ), .A2(\exu._GEN_0 [12] ), .ZN(_01385_ ) );
AOI21_X1 _22062_ ( .A(_08721_ ), .B1(_08723_ ), .B2(_01385_ ), .ZN(_01386_ ) );
NOR2_X1 _22063_ ( .A1(_01347_ ), .A2(_01386_ ), .ZN(_01387_ ) );
AND2_X1 _22064_ ( .A1(\exu.add.io_rs1_data [14] ), .A2(\exu._GEN_0 [14] ), .ZN(_01388_ ) );
AND2_X1 _22065_ ( .A1(_08717_ ), .A2(_01388_ ), .ZN(_01389_ ) );
NOR4_X1 _22066_ ( .A1(_01383_ ), .A2(_01384_ ), .A3(_01387_ ), .A4(_01389_ ), .ZN(_01390_ ) );
AND2_X1 _22067_ ( .A1(_01374_ ), .A2(_01390_ ), .ZN(_01391_ ) );
INV_X1 _22068_ ( .A(_01391_ ), .ZN(_01392_ ) );
NAND2_X1 _22069_ ( .A1(_08751_ ), .A2(_08752_ ), .ZN(_01393_ ) );
INV_X1 _22070_ ( .A(_08754_ ), .ZN(_01394_ ) );
INV_X1 _22071_ ( .A(_08757_ ), .ZN(_01395_ ) );
NOR3_X1 _22072_ ( .A1(_01393_ ), .A2(_01394_ ), .A3(_01395_ ), .ZN(_01396_ ) );
AND2_X1 _22073_ ( .A1(_08743_ ), .A2(_08744_ ), .ZN(_01397_ ) );
AND3_X1 _22074_ ( .A1(_01397_ ), .A2(_08746_ ), .A3(_08748_ ), .ZN(_01398_ ) );
NAND3_X1 _22075_ ( .A1(_01392_ ), .A2(_01396_ ), .A3(_01398_ ), .ZN(_01399_ ) );
AND2_X1 _22076_ ( .A1(\exu.add.io_rs1_data [19] ), .A2(\exu._GEN_0 [19] ), .ZN(_01400_ ) );
AND2_X1 _22077_ ( .A1(\exu.add.io_rs1_data [18] ), .A2(\exu._GEN_0 [18] ), .ZN(_01401_ ) );
AOI21_X1 _22078_ ( .A(_01400_ ), .B1(_08743_ ), .B2(_01401_ ), .ZN(_01402_ ) );
INV_X1 _22079_ ( .A(_01397_ ), .ZN(_01403_ ) );
AND2_X1 _22080_ ( .A1(\exu.add.io_rs1_data [17] ), .A2(\exu._GEN_0 [17] ), .ZN(_01404_ ) );
AND2_X1 _22081_ ( .A1(\exu.add.io_rs1_data [16] ), .A2(\exu._GEN_0 [16] ), .ZN(_01405_ ) );
AOI21_X1 _22082_ ( .A(_01404_ ), .B1(_08746_ ), .B2(_01405_ ), .ZN(_01406_ ) );
OAI21_X1 _22083_ ( .A(_01402_ ), .B1(_01403_ ), .B2(_01406_ ), .ZN(_01407_ ) );
AND2_X1 _22084_ ( .A1(_01407_ ), .A2(_01396_ ), .ZN(_01408_ ) );
AND2_X1 _22085_ ( .A1(\exu.add.io_rs1_data [23] ), .A2(\exu._GEN_0 [23] ), .ZN(_01409_ ) );
INV_X1 _22086_ ( .A(_08756_ ), .ZN(_01410_ ) );
AND2_X1 _22087_ ( .A1(\exu.add.io_rs1_data [20] ), .A2(\exu._GEN_0 [20] ), .ZN(_01411_ ) );
AOI21_X1 _22088_ ( .A(_08755_ ), .B1(_01410_ ), .B2(_01411_ ), .ZN(_01412_ ) );
NOR2_X1 _22089_ ( .A1(_01393_ ), .A2(_01412_ ), .ZN(_01413_ ) );
AND2_X1 _22090_ ( .A1(\exu.add.io_rs1_data [22] ), .A2(\exu._GEN_0 [22] ), .ZN(_01414_ ) );
AND2_X1 _22091_ ( .A1(_08751_ ), .A2(_01414_ ), .ZN(_01415_ ) );
NOR4_X1 _22092_ ( .A1(_01408_ ), .A2(_01409_ ), .A3(_01413_ ), .A4(_01415_ ), .ZN(_01416_ ) );
AOI211_X1 _22093_ ( .A(_01345_ ), .B(_01346_ ), .C1(_01399_ ), .C2(_01416_ ), .ZN(_01417_ ) );
AND2_X1 _22094_ ( .A1(\exu.add.io_rs1_data [25] ), .A2(\exu._GEN_0 [25] ), .ZN(_01418_ ) );
AND2_X1 _22095_ ( .A1(\exu.add.io_rs1_data [24] ), .A2(\exu._GEN_0 [24] ), .ZN(_01419_ ) );
AOI21_X1 _22096_ ( .A(_01418_ ), .B1(_08768_ ), .B2(_01419_ ), .ZN(_01420_ ) );
INV_X1 _22097_ ( .A(_01420_ ), .ZN(_01421_ ) );
OAI211_X1 _22098_ ( .A(_08771_ ), .B(_08772_ ), .C1(_01417_ ), .C2(_01421_ ), .ZN(_01422_ ) );
AND2_X1 _22099_ ( .A1(\exu.add.io_rs1_data [27] ), .A2(\exu._GEN_0 [27] ), .ZN(_01423_ ) );
AND2_X1 _22100_ ( .A1(\exu.add.io_rs1_data [26] ), .A2(\exu._GEN_0 [26] ), .ZN(_01424_ ) );
AOI21_X1 _22101_ ( .A(_01423_ ), .B1(_08771_ ), .B2(_01424_ ), .ZN(_01425_ ) );
AOI21_X1 _22102_ ( .A(_01344_ ), .B1(_01422_ ), .B2(_01425_ ), .ZN(_01426_ ) );
AND2_X1 _22103_ ( .A1(\exu.add.io_rs1_data [28] ), .A2(\exu._GEN_0 [28] ), .ZN(_01427_ ) );
OAI21_X1 _22104_ ( .A(_08764_ ), .B1(_01426_ ), .B2(_01427_ ), .ZN(_01428_ ) );
AND2_X1 _22105_ ( .A1(\exu.add.io_rs1_data [29] ), .A2(\exu._GEN_0 [29] ), .ZN(_01429_ ) );
INV_X1 _22106_ ( .A(_01429_ ), .ZN(_01430_ ) );
AOI21_X1 _22107_ ( .A(_01343_ ), .B1(_01428_ ), .B2(_01430_ ), .ZN(_01431_ ) );
AND2_X1 _22108_ ( .A1(\exu.add.io_rs1_data [30] ), .A2(\exu._GEN_0 [30] ), .ZN(_01432_ ) );
OR3_X1 _22109_ ( .A1(_01431_ ), .A2(_08761_ ), .A3(_01432_ ), .ZN(_01433_ ) );
OAI21_X1 _22110_ ( .A(_08761_ ), .B1(_01431_ ), .B2(_01432_ ), .ZN(_01434_ ) );
AND2_X1 _22111_ ( .A1(_09463_ ), .A2(\exu.add.io_is ), .ZN(_01435_ ) );
BUF_X2 _22112_ ( .A(_01435_ ), .Z(_01436_ ) );
AND3_X1 _22113_ ( .A1(_01433_ ), .A2(_01434_ ), .A3(_01436_ ), .ZN(_01437_ ) );
INV_X1 _22114_ ( .A(fanout_net_12 ), .ZN(_01438_ ) );
NOR2_X1 _22115_ ( .A1(_01438_ ), .A2(fanout_net_26 ), .ZN(_01439_ ) );
BUF_X4 _22116_ ( .A(_01439_ ), .Z(_01440_ ) );
BUF_X4 _22117_ ( .A(_01440_ ), .Z(_01441_ ) );
NAND2_X1 _22118_ ( .A1(_01334_ ), .A2(_01441_ ), .ZN(_01442_ ) );
INV_X2 _22119_ ( .A(\exu.io_in_bits_sra ), .ZN(_01443_ ) );
NOR2_X1 _22120_ ( .A1(_01443_ ), .A2(fanout_net_26 ), .ZN(_01444_ ) );
CLKBUF_X2 _22121_ ( .A(_01444_ ), .Z(_01445_ ) );
INV_X1 _22122_ ( .A(\exu.io_in_bits_or ), .ZN(_01446_ ) );
NOR2_X2 _22123_ ( .A1(_01446_ ), .A2(fanout_net_26 ), .ZN(_01447_ ) );
BUF_X4 _22124_ ( .A(_01447_ ), .Z(_01448_ ) );
OAI21_X1 _22125_ ( .A(_01448_ ), .B1(\exu._GEN_0 [31] ), .B2(\exu.add.io_rs1_data [31] ), .ZN(_01449_ ) );
BUF_X2 _22126_ ( .A(_01211_ ), .Z(_01450_ ) );
NAND3_X1 _22127_ ( .A1(_01201_ ), .A2(_01206_ ), .A3(_01450_ ), .ZN(_01451_ ) );
INV_X1 _22128_ ( .A(\exu.io_in_bits_srl ), .ZN(_01452_ ) );
NOR2_X1 _22129_ ( .A1(_01452_ ), .A2(fanout_net_26 ), .ZN(_01453_ ) );
INV_X1 _22130_ ( .A(_01453_ ), .ZN(_01454_ ) );
BUF_X4 _22131_ ( .A(_01454_ ), .Z(_01455_ ) );
NOR2_X1 _22132_ ( .A1(_01451_ ), .A2(_01455_ ), .ZN(_01456_ ) );
INV_X2 _22133_ ( .A(\exu.io_in_bits_sub ), .ZN(_01457_ ) );
INV_X1 _22134_ ( .A(\exu.auipc.io_is ), .ZN(_01458_ ) );
NOR2_X1 _22135_ ( .A1(_01458_ ), .A2(fanout_net_26 ), .ZN(_01459_ ) );
INV_X1 _22136_ ( .A(_01459_ ), .ZN(_01460_ ) );
AOI21_X1 _22137_ ( .A(_01460_ ), .B1(_09725_ ), .B2(_09726_ ), .ZN(_01461_ ) );
BUF_X2 _22138_ ( .A(_01458_ ), .Z(_01462_ ) );
CLKBUF_X2 _22139_ ( .A(_01462_ ), .Z(_01463_ ) );
AND2_X1 _22140_ ( .A1(_09192_ ), .A2(\exu.io_in_bits_lui ), .ZN(_01464_ ) );
BUF_X2 _22141_ ( .A(_01464_ ), .Z(_01465_ ) );
INV_X1 _22142_ ( .A(exu_io_in_bits_r_lui_$_NOT__A_Y ), .ZN(_01466_ ) );
BUF_X2 _22143_ ( .A(_01466_ ), .Z(_01467_ ) );
AND4_X1 _22144_ ( .A1(_01463_ ), .A2(_01465_ ), .A3(_01467_ ), .A4(\exu.addi.io_imm [31] ), .ZN(_01468_ ) );
OAI21_X1 _22145_ ( .A(_01457_ ), .B1(_01461_ ), .B2(_01468_ ), .ZN(_01469_ ) );
OAI21_X1 _22146_ ( .A(_08760_ ), .B1(_08840_ ), .B2(_08865_ ), .ZN(_01470_ ) );
NAND2_X1 _22147_ ( .A1(_01470_ ), .A2(_08900_ ), .ZN(_01471_ ) );
AOI21_X1 _22148_ ( .A(_08916_ ), .B1(_01471_ ), .B2(_08774_ ), .ZN(_01472_ ) );
NOR3_X1 _22149_ ( .A1(_01472_ ), .A2(_08764_ ), .A3(_08765_ ), .ZN(_01473_ ) );
OR3_X1 _22150_ ( .A1(_01473_ ), .A2(_08870_ ), .A3(_08868_ ), .ZN(_01474_ ) );
NAND2_X1 _22151_ ( .A1(_01474_ ), .A2(_01343_ ), .ZN(_01475_ ) );
AND3_X1 _22152_ ( .A1(_01475_ ), .A2(_08761_ ), .A3(_08873_ ), .ZN(_01476_ ) );
NOR2_X1 _22153_ ( .A1(_01457_ ), .A2(fanout_net_26 ), .ZN(_01477_ ) );
BUF_X2 _22154_ ( .A(_01477_ ), .Z(_01478_ ) );
OAI21_X1 _22155_ ( .A(_01478_ ), .B1(_09428_ ), .B2(_08761_ ), .ZN(_01479_ ) );
OAI21_X1 _22156_ ( .A(_01469_ ), .B1(_01476_ ), .B2(_01479_ ), .ZN(_01480_ ) );
BUF_X4 _22157_ ( .A(_01452_ ), .Z(_01481_ ) );
AOI21_X1 _22158_ ( .A(_01456_ ), .B1(_01480_ ), .B2(_01481_ ), .ZN(_01482_ ) );
OAI21_X1 _22159_ ( .A(_01449_ ), .B1(_01482_ ), .B2(\exu.io_in_bits_or ), .ZN(_01483_ ) );
AOI221_X4 _22160_ ( .A(fanout_net_4 ), .B1(_01177_ ), .B2(_01445_ ), .C1(_01483_ ), .C2(_01443_ ), .ZN(_01484_ ) );
INV_X1 _22161_ ( .A(fanout_net_4 ), .ZN(_01485_ ) );
BUF_X4 _22162_ ( .A(_01485_ ), .Z(_01486_ ) );
NOR2_X1 _22163_ ( .A1(_01486_ ), .A2(fanout_net_26 ), .ZN(_01487_ ) );
NAND3_X1 _22164_ ( .A1(_01487_ ), .A2(\exu._GEN_0 [31] ), .A3(\exu.add.io_rs1_data [31] ), .ZN(_01488_ ) );
AOI211_X1 _22165_ ( .A(\exu.io_in_bits_xor ), .B(_01484_ ), .C1(fanout_net_4 ), .C2(_01488_ ), .ZN(_01489_ ) );
INV_X1 _22166_ ( .A(\exu.io_in_bits_xor ), .ZN(_01490_ ) );
NOR2_X1 _22167_ ( .A1(_01490_ ), .A2(fanout_net_26 ), .ZN(_01491_ ) );
BUF_X4 _22168_ ( .A(_01491_ ), .Z(_01492_ ) );
BUF_X4 _22169_ ( .A(_01492_ ), .Z(_01493_ ) );
AOI21_X1 _22170_ ( .A(_01489_ ), .B1(_08761_ ), .B2(_01493_ ), .ZN(_01494_ ) );
OAI21_X1 _22171_ ( .A(_01442_ ), .B1(_01494_ ), .B2(fanout_net_12 ), .ZN(_01495_ ) );
NOR2_X1 _22172_ ( .A1(\exu.add.io_is ), .A2(\exu.io_in_bits_sltu ), .ZN(_01496_ ) );
INV_X1 _22173_ ( .A(\exu.io_in_bits_slt ), .ZN(_01497_ ) );
AND2_X2 _22174_ ( .A1(_01496_ ), .A2(_01497_ ), .ZN(_01498_ ) );
AOI21_X1 _22175_ ( .A(_01437_ ), .B1(_01495_ ), .B2(_01498_ ), .ZN(_01499_ ) );
OAI221_X1 _22176_ ( .A(_01341_ ), .B1(_09733_ ), .B2(_01342_ ), .C1(_01499_ ), .C2(\exu.io_in_bits_jal ), .ZN(_01500_ ) );
BUF_X4 _22177_ ( .A(_10820_ ), .Z(_01501_ ) );
AND3_X1 _22178_ ( .A1(_09731_ ), .A2(_09732_ ), .A3(_09460_ ), .ZN(_01502_ ) );
OAI211_X1 _22179_ ( .A(_01500_ ), .B(_01501_ ), .C1(_01341_ ), .C2(_01502_ ), .ZN(_01503_ ) );
BUF_X4 _22180_ ( .A(_01219_ ), .Z(_01504_ ) );
BUF_X4 _22181_ ( .A(_01504_ ), .Z(_01505_ ) );
MUX2_X1 _22182_ ( .A(_01339_ ), .B(_01503_ ), .S(_01505_ ), .Z(_01506_ ) );
BUF_X4 _22183_ ( .A(_01214_ ), .Z(_01507_ ) );
MUX2_X1 _22184_ ( .A(_01218_ ), .B(_01506_ ), .S(_01507_ ), .Z(_01508_ ) );
BUF_X4 _22185_ ( .A(_01184_ ), .Z(_01509_ ) );
BUF_X4 _22186_ ( .A(_01509_ ), .Z(_01510_ ) );
MUX2_X1 _22187_ ( .A(_01187_ ), .B(_01508_ ), .S(_01510_ ), .Z(_01511_ ) );
BUF_X4 _22188_ ( .A(_01181_ ), .Z(_01512_ ) );
AOI21_X1 _22189_ ( .A(_01183_ ), .B1(_01511_ ), .B2(_01512_ ), .ZN(_01513_ ) );
NAND2_X1 _22190_ ( .A1(\exu.add.io_rs1_data [31] ), .A2(\exu.addi.io_imm [31] ), .ZN(_01514_ ) );
BUF_X4 _22191_ ( .A(_01176_ ), .Z(_01515_ ) );
NOR3_X1 _22192_ ( .A1(_01514_ ), .A2(_01515_ ), .A3(fanout_net_26 ), .ZN(_01516_ ) );
OAI21_X1 _22193_ ( .A(_01175_ ), .B1(_01513_ ), .B2(_01516_ ), .ZN(_01517_ ) );
NOR2_X1 _22194_ ( .A1(_01174_ ), .A2(fanout_net_26 ), .ZN(_01518_ ) );
BUF_X4 _22195_ ( .A(_01518_ ), .Z(_01519_ ) );
NAND2_X1 _22196_ ( .A1(_09766_ ), .A2(_01519_ ), .ZN(_01520_ ) );
AOI21_X1 _22197_ ( .A(_01173_ ), .B1(_01517_ ), .B2(_01520_ ), .ZN(_01521_ ) );
INV_X1 _22198_ ( .A(\exu.addi.io_is ), .ZN(_01522_ ) );
NOR2_X1 _22199_ ( .A1(_01522_ ), .A2(fanout_net_26 ), .ZN(_01523_ ) );
AND2_X1 _22200_ ( .A1(\exu.addi._io_rd_T_4 [31] ), .A2(_01523_ ), .ZN(_01524_ ) );
OAI21_X1 _22201_ ( .A(_01108_ ), .B1(_01521_ ), .B2(_01524_ ), .ZN(_01525_ ) );
INV_X1 _22202_ ( .A(_01525_ ), .ZN(_01526_ ) );
NOR3_X1 _22203_ ( .A1(_01109_ ), .A2(fanout_net_26 ), .A3(_09741_ ), .ZN(_01527_ ) );
NOR2_X1 _22204_ ( .A1(_01526_ ), .A2(_01527_ ), .ZN(_01528_ ) );
INV_X1 _22205_ ( .A(_01528_ ), .ZN(\exu.io_out_bits_rd_wdata [31] ) );
NOR2_X1 _22206_ ( .A1(_01180_ ), .A2(fanout_net_26 ), .ZN(_01529_ ) );
AND2_X2 _22207_ ( .A1(_01529_ ), .A2(_01178_ ), .ZN(_01530_ ) );
NAND2_X1 _22208_ ( .A1(_01180_ ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_11_B_$_ANDNOT__Y_B ), .ZN(_01531_ ) );
NAND2_X1 _22209_ ( .A1(\exu.io_in_bits_srai ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__A_B ), .ZN(_01532_ ) );
NAND2_X1 _22210_ ( .A1(_01531_ ), .A2(_01532_ ), .ZN(_01533_ ) );
NOR2_X1 _22211_ ( .A1(_01533_ ), .A2(_01177_ ), .ZN(_01534_ ) );
INV_X1 _22212_ ( .A(_01534_ ), .ZN(_01535_ ) );
BUF_X2 _22213_ ( .A(_01535_ ), .Z(_01536_ ) );
BUF_X2 _22214_ ( .A(_01536_ ), .Z(_01537_ ) );
NAND2_X1 _22215_ ( .A1(_01180_ ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_12_B_$_ANDNOT__Y_B ), .ZN(_01538_ ) );
NAND2_X1 _22216_ ( .A1(\exu.io_in_bits_srai ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__A_B ), .ZN(_01539_ ) );
NAND2_X1 _22217_ ( .A1(_01538_ ), .A2(_01539_ ), .ZN(_01540_ ) );
BUF_X4 _22218_ ( .A(_01540_ ), .Z(_01541_ ) );
NOR2_X1 _22219_ ( .A1(_01541_ ), .A2(_01177_ ), .ZN(_01542_ ) );
NAND2_X1 _22220_ ( .A1(_01180_ ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_13_B_$_ANDNOT__Y_B ), .ZN(_01543_ ) );
NAND2_X1 _22221_ ( .A1(\exu.io_in_bits_srai ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__A_B ), .ZN(_01544_ ) );
NAND2_X1 _22222_ ( .A1(_01543_ ), .A2(_01544_ ), .ZN(_01545_ ) );
BUF_X4 _22223_ ( .A(_01545_ ), .Z(_01546_ ) );
BUF_X2 _22224_ ( .A(_01546_ ), .Z(_01547_ ) );
NOR2_X1 _22225_ ( .A1(_01547_ ), .A2(_01177_ ), .ZN(_01548_ ) );
INV_X1 _22226_ ( .A(_01548_ ), .ZN(_01549_ ) );
NAND2_X1 _22227_ ( .A1(_01180_ ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_14_B_$_ANDNOT__Y_B ), .ZN(_01550_ ) );
NAND2_X1 _22228_ ( .A1(\exu.io_in_bits_srai ), .A2(\exu.io_out_bits_wdata_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__A_B ), .ZN(_01551_ ) );
AND3_X1 _22229_ ( .A1(_01550_ ), .A2(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B ), .A3(_01551_ ), .ZN(_01552_ ) );
NAND2_X1 _22230_ ( .A1(_01180_ ), .A2(_01089_ ), .ZN(_01553_ ) );
NAND2_X1 _22231_ ( .A1(_01191_ ), .A2(\exu.io_in_bits_srai ), .ZN(_01554_ ) );
AND2_X1 _22232_ ( .A1(_01553_ ), .A2(_01554_ ), .ZN(_01555_ ) );
BUF_X4 _22233_ ( .A(_01555_ ), .Z(_01556_ ) );
MUX2_X1 _22234_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B ), .S(_01556_ ), .Z(_01557_ ) );
NAND2_X1 _22235_ ( .A1(_01550_ ), .A2(_01551_ ), .ZN(_01558_ ) );
BUF_X4 _22236_ ( .A(_01558_ ), .Z(_01559_ ) );
AOI21_X1 _22237_ ( .A(_01552_ ), .B1(_01557_ ), .B2(_01559_ ), .ZN(_01560_ ) );
INV_X1 _22238_ ( .A(_01545_ ), .ZN(_01561_ ) );
BUF_X4 _22239_ ( .A(_01561_ ), .Z(_01562_ ) );
OAI21_X1 _22240_ ( .A(_01549_ ), .B1(_01560_ ), .B2(_01562_ ), .ZN(_01563_ ) );
BUF_X4 _22241_ ( .A(_01541_ ), .Z(_01564_ ) );
AOI21_X1 _22242_ ( .A(_01542_ ), .B1(_01563_ ), .B2(_01564_ ), .ZN(_01565_ ) );
INV_X1 _22243_ ( .A(_01533_ ), .ZN(_01566_ ) );
BUF_X4 _22244_ ( .A(_01566_ ), .Z(_01567_ ) );
BUF_X4 _22245_ ( .A(_01567_ ), .Z(_01568_ ) );
OAI211_X1 _22246_ ( .A(_01530_ ), .B(_01537_ ), .C1(_01565_ ), .C2(_01568_ ), .ZN(_01569_ ) );
AND2_X1 _22247_ ( .A1(_01501_ ), .A2(_01505_ ), .ZN(_01570_ ) );
BUF_X4 _22248_ ( .A(_09410_ ), .Z(_01571_ ) );
INV_X1 _22249_ ( .A(_01498_ ), .ZN(_01572_ ) );
BUF_X4 _22250_ ( .A(_01572_ ), .Z(_01573_ ) );
BUF_X4 _22251_ ( .A(_01573_ ), .Z(_01574_ ) );
BUF_X2 _22252_ ( .A(_10698_ ), .Z(_01575_ ) );
NAND3_X1 _22253_ ( .A1(_01432_ ), .A2(_01575_ ), .A3(fanout_net_4 ), .ZN(_01576_ ) );
OAI21_X1 _22254_ ( .A(_01537_ ), .B1(_01565_ ), .B2(_01568_ ), .ZN(_01577_ ) );
INV_X1 _22255_ ( .A(_01444_ ), .ZN(_01578_ ) );
BUF_X4 _22256_ ( .A(_01578_ ), .Z(_01579_ ) );
NOR2_X1 _22257_ ( .A1(_01577_ ), .A2(_01579_ ), .ZN(_01580_ ) );
BUF_X4 _22258_ ( .A(_01448_ ), .Z(_01581_ ) );
OAI21_X1 _22259_ ( .A(_01581_ ), .B1(\exu.add.io_rs1_data [30] ), .B2(\exu._GEN_0 [30] ), .ZN(_01582_ ) );
AND2_X2 _22260_ ( .A1(_01189_ ), .A2(_01192_ ), .ZN(_01583_ ) );
MUX2_X1 _22261_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B ), .S(_01583_ ), .Z(_01584_ ) );
INV_X1 _22262_ ( .A(_01197_ ), .ZN(_01585_ ) );
BUF_X4 _22263_ ( .A(_01585_ ), .Z(_01586_ ) );
BUF_X4 _22264_ ( .A(_01586_ ), .Z(_01587_ ) );
NOR2_X1 _22265_ ( .A1(_01584_ ), .A2(_01587_ ), .ZN(_01588_ ) );
BUF_X4 _22266_ ( .A(_01200_ ), .Z(_01589_ ) );
BUF_X4 _22267_ ( .A(_01589_ ), .Z(_01590_ ) );
BUF_X2 _22268_ ( .A(_01204_ ), .Z(_01591_ ) );
AND3_X1 _22269_ ( .A1(_01588_ ), .A2(_01590_ ), .A3(_01591_ ), .ZN(_01592_ ) );
BUF_X2 _22270_ ( .A(_01453_ ), .Z(_01593_ ) );
CLKBUF_X2 _22271_ ( .A(_01593_ ), .Z(_01594_ ) );
AND3_X1 _22272_ ( .A1(_01592_ ), .A2(_01212_ ), .A3(_01594_ ), .ZN(_01595_ ) );
INV_X1 _22273_ ( .A(_01477_ ), .ZN(_01596_ ) );
BUF_X2 _22274_ ( .A(_01596_ ), .Z(_01597_ ) );
AOI21_X1 _22275_ ( .A(_01597_ ), .B1(_01474_ ), .B2(_01343_ ), .ZN(_01598_ ) );
OAI21_X1 _22276_ ( .A(_01598_ ), .B1(_01343_ ), .B2(_01474_ ), .ZN(_01599_ ) );
CLKBUF_X2 _22277_ ( .A(_01465_ ), .Z(_01600_ ) );
CLKBUF_X2 _22278_ ( .A(_01600_ ), .Z(_01601_ ) );
CLKBUF_X2 _22279_ ( .A(_01462_ ), .Z(_01602_ ) );
CLKBUF_X2 _22280_ ( .A(_01467_ ), .Z(_01603_ ) );
CLKBUF_X2 _22281_ ( .A(_01603_ ), .Z(_01604_ ) );
AND4_X1 _22282_ ( .A1(\exu.addi.io_imm [30] ), .A2(_01601_ ), .A3(_01602_ ), .A4(_01604_ ), .ZN(_01605_ ) );
BUF_X4 _22283_ ( .A(_01459_ ), .Z(_01606_ ) );
BUF_X4 _22284_ ( .A(_01606_ ), .Z(_01607_ ) );
AOI21_X1 _22285_ ( .A(_01605_ ), .B1(_09665_ ), .B2(_01607_ ), .ZN(_01608_ ) );
OAI21_X1 _22286_ ( .A(_01599_ ), .B1(_01608_ ), .B2(\exu.io_in_bits_sub ), .ZN(_01609_ ) );
BUF_X4 _22287_ ( .A(_01481_ ), .Z(_01610_ ) );
AOI21_X1 _22288_ ( .A(_01595_ ), .B1(_01609_ ), .B2(_01610_ ), .ZN(_01611_ ) );
OAI21_X1 _22289_ ( .A(_01582_ ), .B1(_01611_ ), .B2(\exu.io_in_bits_or ), .ZN(_01612_ ) );
BUF_X4 _22290_ ( .A(_01443_ ), .Z(_01613_ ) );
BUF_X4 _22291_ ( .A(_01613_ ), .Z(_01614_ ) );
AOI21_X1 _22292_ ( .A(_01580_ ), .B1(_01612_ ), .B2(_01614_ ), .ZN(_01615_ ) );
OAI21_X1 _22293_ ( .A(_01576_ ), .B1(_01615_ ), .B2(fanout_net_4 ), .ZN(_01616_ ) );
BUF_X4 _22294_ ( .A(_01490_ ), .Z(_01617_ ) );
BUF_X4 _22295_ ( .A(_01617_ ), .Z(_01618_ ) );
AOI221_X4 _22296_ ( .A(fanout_net_12 ), .B1(_08762_ ), .B2(_01493_ ), .C1(_01616_ ), .C2(_01618_ ), .ZN(_01619_ ) );
NAND2_X1 _22297_ ( .A1(_01264_ ), .A2(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01620_ ) );
NAND3_X1 _22298_ ( .A1(_01285_ ), .A2(_01286_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01621_ ) );
NAND2_X1 _22299_ ( .A1(_01620_ ), .A2(_01621_ ), .ZN(_01622_ ) );
NAND2_X1 _22300_ ( .A1(_01622_ ), .A2(_01235_ ), .ZN(_01623_ ) );
AND3_X1 _22301_ ( .A1(_01285_ ), .A2(_01286_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01624_ ) );
AOI21_X1 _22302_ ( .A(_01255_ ), .B1(_01285_ ), .B2(_01286_ ), .ZN(_01625_ ) );
OAI21_X1 _22303_ ( .A(_01290_ ), .B1(_01624_ ), .B2(_01625_ ), .ZN(_01626_ ) );
NAND2_X1 _22304_ ( .A1(_01623_ ), .A2(_01626_ ), .ZN(_01627_ ) );
NAND2_X1 _22305_ ( .A1(_01627_ ), .A2(_01306_ ), .ZN(_01628_ ) );
INV_X1 _22306_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01629_ ) );
AND3_X1 _22307_ ( .A1(_01285_ ), .A2(_01286_ ), .A3(_01629_ ), .ZN(_01630_ ) );
AOI21_X1 _22308_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B1(_01285_ ), .B2(_01286_ ), .ZN(_01631_ ) );
NOR2_X1 _22309_ ( .A1(_01630_ ), .A2(_01631_ ), .ZN(_01632_ ) );
NAND2_X1 _22310_ ( .A1(_01632_ ), .A2(_01291_ ), .ZN(_01633_ ) );
AOI21_X1 _22311_ ( .A(_08821_ ), .B1(_01309_ ), .B2(_01310_ ), .ZN(_01634_ ) );
OAI21_X1 _22312_ ( .A(_01633_ ), .B1(_01291_ ), .B2(_01634_ ), .ZN(_01635_ ) );
NAND2_X1 _22313_ ( .A1(_01635_ ), .A2(_01325_ ), .ZN(_01636_ ) );
NAND3_X1 _22314_ ( .A1(_01628_ ), .A2(_01246_ ), .A3(_01636_ ), .ZN(_01637_ ) );
INV_X1 _22315_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01638_ ) );
OR2_X1 _22316_ ( .A1(_01230_ ), .A2(_01638_ ), .ZN(_01639_ ) );
OAI211_X1 _22317_ ( .A(_01639_ ), .B(_01248_ ), .C1(_01274_ ), .C2(_01264_ ), .ZN(_01640_ ) );
NAND3_X1 _22318_ ( .A1(_01221_ ), .A2(_01223_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01641_ ) );
INV_X1 _22319_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01642_ ) );
OAI211_X1 _22320_ ( .A(_01234_ ), .B(_01641_ ), .C1(_01230_ ), .C2(_01642_ ), .ZN(_01643_ ) );
NAND3_X1 _22321_ ( .A1(_01640_ ), .A2(_01306_ ), .A3(_01643_ ), .ZN(_01644_ ) );
NAND3_X1 _22322_ ( .A1(_01285_ ), .A2(_01286_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01645_ ) );
OAI211_X1 _22323_ ( .A(_01290_ ), .B(_01645_ ), .C1(_01273_ ), .C2(_01263_ ), .ZN(_01646_ ) );
AND3_X1 _22324_ ( .A1(_01285_ ), .A2(_01286_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01647_ ) );
INV_X1 _22325_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01648_ ) );
AOI21_X1 _22326_ ( .A(_01648_ ), .B1(_01285_ ), .B2(_01286_ ), .ZN(_01649_ ) );
OR2_X1 _22327_ ( .A1(_01647_ ), .A2(_01649_ ), .ZN(_01650_ ) );
OAI211_X1 _22328_ ( .A(_01241_ ), .B(_01646_ ), .C1(_01650_ ), .C2(_01299_ ), .ZN(_01651_ ) );
NAND3_X1 _22329_ ( .A1(_01644_ ), .A2(_01271_ ), .A3(_01651_ ), .ZN(_01652_ ) );
NAND2_X1 _22330_ ( .A1(_01637_ ), .A2(_01652_ ), .ZN(_01653_ ) );
BUF_X2 _22331_ ( .A(_01331_ ), .Z(_01654_ ) );
NAND2_X1 _22332_ ( .A1(_01653_ ), .A2(_01654_ ), .ZN(_01655_ ) );
AND3_X1 _22333_ ( .A1(_01221_ ), .A2(_01223_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01656_ ) );
INV_X1 _22334_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01657_ ) );
AOI21_X1 _22335_ ( .A(_01657_ ), .B1(_01221_ ), .B2(_01223_ ), .ZN(_01658_ ) );
OAI21_X1 _22336_ ( .A(_01290_ ), .B1(_01656_ ), .B2(_01658_ ), .ZN(_01659_ ) );
AND3_X1 _22337_ ( .A1(_01221_ ), .A2(_01223_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01660_ ) );
INV_X1 _22338_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01661_ ) );
AOI21_X1 _22339_ ( .A(_01661_ ), .B1(_01221_ ), .B2(_01223_ ), .ZN(_01662_ ) );
OAI21_X1 _22340_ ( .A(_01234_ ), .B1(_01660_ ), .B2(_01662_ ), .ZN(_01663_ ) );
AND3_X1 _22341_ ( .A1(_01659_ ), .A2(_01663_ ), .A3(_01325_ ), .ZN(_01664_ ) );
NAND3_X1 _22342_ ( .A1(_01309_ ), .A2(_01310_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01665_ ) );
INV_X1 _22343_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01666_ ) );
OAI211_X1 _22344_ ( .A(_01299_ ), .B(_01665_ ), .C1(_01297_ ), .C2(_01666_ ), .ZN(_01667_ ) );
AND3_X1 _22345_ ( .A1(_01309_ ), .A2(_01310_ ), .A3(_01323_ ), .ZN(_01668_ ) );
AOI21_X1 _22346_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_01309_ ), .B2(_01310_ ), .ZN(_01669_ ) );
OAI21_X1 _22347_ ( .A(_01254_ ), .B1(_01668_ ), .B2(_01669_ ), .ZN(_01670_ ) );
AOI21_X1 _22348_ ( .A(_01325_ ), .B1(_01667_ ), .B2(_01670_ ), .ZN(_01671_ ) );
NOR2_X1 _22349_ ( .A1(_01664_ ), .A2(_01671_ ), .ZN(_01672_ ) );
NAND3_X1 _22350_ ( .A1(_01309_ ), .A2(_01310_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01673_ ) );
OAI211_X1 _22351_ ( .A(_01254_ ), .B(_01673_ ), .C1(_01297_ ), .C2(_01283_ ), .ZN(_01674_ ) );
INV_X1 _22352_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01675_ ) );
AND3_X1 _22353_ ( .A1(_01309_ ), .A2(_01310_ ), .A3(_01675_ ), .ZN(_01676_ ) );
AOI21_X1 _22354_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B1(_01309_ ), .B2(_01310_ ), .ZN(_01677_ ) );
OAI21_X1 _22355_ ( .A(_01299_ ), .B1(_01676_ ), .B2(_01677_ ), .ZN(_01678_ ) );
AND2_X1 _22356_ ( .A1(_01674_ ), .A2(_01678_ ), .ZN(_01679_ ) );
AND3_X1 _22357_ ( .A1(_01309_ ), .A2(_01310_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01680_ ) );
AOI21_X1 _22358_ ( .A(_01301_ ), .B1(_01309_ ), .B2(_01310_ ), .ZN(_01681_ ) );
OR2_X1 _22359_ ( .A1(_01680_ ), .A2(_01681_ ), .ZN(_01682_ ) );
MUX2_X1 _22360_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(_01297_ ), .Z(_01683_ ) );
MUX2_X1 _22361_ ( .A(_01682_ ), .B(_01683_ ), .S(_01299_ ), .Z(_01684_ ) );
MUX2_X1 _22362_ ( .A(_01679_ ), .B(_01684_ ), .S(_01306_ ), .Z(_01685_ ) );
BUF_X4 _22363_ ( .A(_01271_ ), .Z(_01686_ ) );
MUX2_X1 _22364_ ( .A(_01672_ ), .B(_01685_ ), .S(_01686_ ), .Z(_01687_ ) );
OAI21_X1 _22365_ ( .A(_01655_ ), .B1(_01687_ ), .B2(_01654_ ), .ZN(_01688_ ) );
BUF_X4 _22366_ ( .A(_01441_ ), .Z(_01689_ ) );
NAND2_X1 _22367_ ( .A1(_01688_ ), .A2(_01689_ ), .ZN(_01690_ ) );
AOI211_X1 _22368_ ( .A(_01574_ ), .B(_01619_ ), .C1(fanout_net_12 ), .C2(_01690_ ), .ZN(_01691_ ) );
AND3_X1 _22369_ ( .A1(_01428_ ), .A2(_01343_ ), .A3(_01430_ ), .ZN(_01692_ ) );
INV_X1 _22370_ ( .A(_01436_ ), .ZN(_01693_ ) );
BUF_X4 _22371_ ( .A(_01693_ ), .Z(_01694_ ) );
NOR3_X1 _22372_ ( .A1(_01692_ ), .A2(_01431_ ), .A3(_01694_ ), .ZN(_01695_ ) );
OAI21_X1 _22373_ ( .A(_01571_ ), .B1(_01691_ ), .B2(_01695_ ), .ZN(_01696_ ) );
NAND2_X1 _22374_ ( .A1(_09672_ ), .A2(_09452_ ), .ZN(_01697_ ) );
AOI21_X1 _22375_ ( .A(\exu.io_in_bits_jalr ), .B1(_01696_ ), .B2(_01697_ ), .ZN(_01698_ ) );
CLKBUF_X2 _22376_ ( .A(_09460_ ), .Z(_01699_ ) );
AND2_X1 _22377_ ( .A1(_09672_ ), .A2(_01699_ ), .ZN(_01700_ ) );
OAI21_X1 _22378_ ( .A(_01570_ ), .B1(_01698_ ), .B2(_01700_ ), .ZN(_01701_ ) );
BUF_X4 _22379_ ( .A(_01338_ ), .Z(_01702_ ) );
NAND2_X1 _22380_ ( .A1(_01688_ ), .A2(_01702_ ), .ZN(_01703_ ) );
NAND3_X1 _22381_ ( .A1(_01701_ ), .A2(_01507_ ), .A3(_01703_ ), .ZN(_01704_ ) );
BUF_X4 _22382_ ( .A(_01507_ ), .Z(_01705_ ) );
AND3_X1 _22383_ ( .A1(_01592_ ), .A2(_01213_ ), .A3(_01217_ ), .ZN(_01706_ ) );
OAI211_X1 _22384_ ( .A(_01704_ ), .B(_01510_ ), .C1(_01705_ ), .C2(_01706_ ), .ZN(_01707_ ) );
OAI21_X1 _22385_ ( .A(_01186_ ), .B1(\exu.add.io_rs1_data [30] ), .B2(\exu.addi.io_imm [30] ), .ZN(_01708_ ) );
AND2_X1 _22386_ ( .A1(_01708_ ), .A2(_01181_ ), .ZN(_01709_ ) );
AOI221_X4 _22387_ ( .A(fanout_net_5 ), .B1(\exu.io_in_bits_srai ), .B2(_01569_ ), .C1(_01707_ ), .C2(_01709_ ), .ZN(_01710_ ) );
AND3_X1 _22388_ ( .A1(_09707_ ), .A2(_10843_ ), .A3(fanout_net_5 ), .ZN(_01711_ ) );
OAI21_X1 _22389_ ( .A(_01175_ ), .B1(_01710_ ), .B2(_01711_ ), .ZN(_01712_ ) );
NAND2_X1 _22390_ ( .A1(_09709_ ), .A2(_01519_ ), .ZN(_01713_ ) );
AOI21_X1 _22391_ ( .A(_01173_ ), .B1(_01712_ ), .B2(_01713_ ), .ZN(_01714_ ) );
AND2_X1 _22392_ ( .A1(\exu.addi._io_rd_T_4 [30] ), .A2(_01523_ ), .ZN(_01715_ ) );
OAI21_X1 _22393_ ( .A(_01108_ ), .B1(_01714_ ), .B2(_01715_ ), .ZN(_01716_ ) );
INV_X1 _22394_ ( .A(_01716_ ), .ZN(_01717_ ) );
INV_X1 _22395_ ( .A(_01108_ ), .ZN(_01718_ ) );
AND3_X1 _22396_ ( .A1(_01718_ ), .A2(_10844_ ), .A3(\exu.csrrs.io_csr_rdata [30] ), .ZN(_01719_ ) );
NOR2_X1 _22397_ ( .A1(_01717_ ), .A2(_01719_ ), .ZN(_01720_ ) );
INV_X1 _22398_ ( .A(_01720_ ), .ZN(\exu.io_out_bits_rd_wdata [30] ) );
BUF_X4 _22399_ ( .A(_01108_ ), .Z(_01721_ ) );
BUF_X4 _22400_ ( .A(_01172_ ), .Z(_01722_ ) );
BUF_X4 _22401_ ( .A(_01175_ ), .Z(_01723_ ) );
INV_X1 _22402_ ( .A(_01558_ ), .ZN(_01724_ ) );
BUF_X4 _22403_ ( .A(_01724_ ), .Z(_01725_ ) );
BUF_X2 _22404_ ( .A(_01553_ ), .Z(_01726_ ) );
BUF_X2 _22405_ ( .A(_01554_ ), .Z(_01727_ ) );
NAND3_X1 _22406_ ( .A1(_01726_ ), .A2(_01727_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01728_ ) );
BUF_X4 _22407_ ( .A(_01556_ ), .Z(_01729_ ) );
OAI211_X1 _22408_ ( .A(_01725_ ), .B(_01728_ ), .C1(_01729_ ), .C2(_01315_ ), .ZN(_01730_ ) );
NAND3_X1 _22409_ ( .A1(_01553_ ), .A2(_01554_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01731_ ) );
OAI211_X1 _22410_ ( .A(_01559_ ), .B(_01731_ ), .C1(_01729_ ), .C2(_01312_ ), .ZN(_01732_ ) );
AND3_X1 _22411_ ( .A1(_01730_ ), .A2(_01732_ ), .A3(_01547_ ), .ZN(_01733_ ) );
BUF_X4 _22412_ ( .A(_01546_ ), .Z(_01734_ ) );
INV_X1 _22413_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01735_ ) );
NAND3_X1 _22414_ ( .A1(_01726_ ), .A2(_01727_ ), .A3(_01735_ ), .ZN(_01736_ ) );
OAI211_X1 _22415_ ( .A(_01559_ ), .B(_01736_ ), .C1(_01729_ ), .C2(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01737_ ) );
AND3_X1 _22416_ ( .A1(_01553_ ), .A2(_01554_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01738_ ) );
AOI21_X1 _22417_ ( .A(_01293_ ), .B1(_01553_ ), .B2(_01554_ ), .ZN(_01739_ ) );
OAI21_X1 _22418_ ( .A(_01725_ ), .B1(_01738_ ), .B2(_01739_ ), .ZN(_01740_ ) );
AOI21_X1 _22419_ ( .A(_01734_ ), .B1(_01737_ ), .B2(_01740_ ), .ZN(_01741_ ) );
NOR2_X1 _22420_ ( .A1(_01733_ ), .A2(_01741_ ), .ZN(_01742_ ) );
MUX2_X1 _22421_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .S(_01556_ ), .Z(_01743_ ) );
AOI21_X1 _22422_ ( .A(_01552_ ), .B1(_01743_ ), .B2(_01558_ ), .ZN(_01744_ ) );
MUX2_X1 _22423_ ( .A(_01177_ ), .B(_01744_ ), .S(_01545_ ), .Z(_01745_ ) );
INV_X1 _22424_ ( .A(_01540_ ), .ZN(_01746_ ) );
BUF_X4 _22425_ ( .A(_01746_ ), .Z(_01747_ ) );
BUF_X2 _22426_ ( .A(_01747_ ), .Z(_01748_ ) );
MUX2_X1 _22427_ ( .A(_01742_ ), .B(_01745_ ), .S(_01748_ ), .Z(_01749_ ) );
OAI21_X1 _22428_ ( .A(_01537_ ), .B1(_01749_ ), .B2(_01568_ ), .ZN(_01750_ ) );
INV_X1 _22429_ ( .A(_01530_ ), .ZN(_01751_ ) );
BUF_X4 _22430_ ( .A(_01751_ ), .Z(_01752_ ) );
NOR2_X1 _22431_ ( .A1(_01750_ ), .A2(_01752_ ), .ZN(_01753_ ) );
OAI21_X1 _22432_ ( .A(_01515_ ), .B1(_01753_ ), .B2(_01512_ ), .ZN(_01754_ ) );
BUF_X4 _22433_ ( .A(_01186_ ), .Z(_01755_ ) );
OAI21_X1 _22434_ ( .A(_01755_ ), .B1(\exu.add.io_rs1_data [21] ), .B2(\exu.addi.io_imm [21] ), .ZN(_01756_ ) );
AND3_X1 _22435_ ( .A1(_01189_ ), .A2(_01192_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01757_ ) );
BUF_X2 _22436_ ( .A(_01189_ ), .Z(_01758_ ) );
BUF_X2 _22437_ ( .A(_01192_ ), .Z(_01759_ ) );
AOI21_X1 _22438_ ( .A(_01315_ ), .B1(_01758_ ), .B2(_01759_ ), .ZN(_01760_ ) );
BUF_X4 _22439_ ( .A(_01197_ ), .Z(_01761_ ) );
OR3_X1 _22440_ ( .A1(_01757_ ), .A2(_01760_ ), .A3(_01761_ ), .ZN(_01762_ ) );
BUF_X4 _22441_ ( .A(_01761_ ), .Z(_01763_ ) );
BUF_X2 _22442_ ( .A(_01758_ ), .Z(_01764_ ) );
BUF_X2 _22443_ ( .A(_01759_ ), .Z(_01765_ ) );
NAND3_X1 _22444_ ( .A1(_01764_ ), .A2(_01765_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01766_ ) );
BUF_X4 _22445_ ( .A(_01583_ ), .Z(_01767_ ) );
OAI211_X1 _22446_ ( .A(_01763_ ), .B(_01766_ ), .C1(_01767_ ), .C2(_01312_ ), .ZN(_01768_ ) );
NAND3_X1 _22447_ ( .A1(_01762_ ), .A2(_01590_ ), .A3(_01768_ ), .ZN(_01769_ ) );
INV_X2 _22448_ ( .A(_01200_ ), .ZN(_01770_ ) );
BUF_X4 _22449_ ( .A(_01770_ ), .Z(_01771_ ) );
AND3_X1 _22450_ ( .A1(_01189_ ), .A2(_01192_ ), .A3(_01735_ ), .ZN(_01772_ ) );
AOI21_X1 _22451_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01189_ ), .B2(_01192_ ), .ZN(_01773_ ) );
OAI21_X1 _22452_ ( .A(_01763_ ), .B1(_01772_ ), .B2(_01773_ ), .ZN(_01774_ ) );
AND3_X1 _22453_ ( .A1(_01758_ ), .A2(_01759_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01775_ ) );
AOI21_X1 _22454_ ( .A(_01293_ ), .B1(_01758_ ), .B2(_01759_ ), .ZN(_01776_ ) );
OR2_X1 _22455_ ( .A1(_01775_ ), .A2(_01776_ ), .ZN(_01777_ ) );
BUF_X4 _22456_ ( .A(_01761_ ), .Z(_01778_ ) );
OAI211_X1 _22457_ ( .A(_01771_ ), .B(_01774_ ), .C1(_01777_ ), .C2(_01778_ ), .ZN(_01779_ ) );
NAND3_X1 _22458_ ( .A1(_01769_ ), .A2(_01779_ ), .A3(_01206_ ), .ZN(_01780_ ) );
BUF_X2 _22459_ ( .A(_01586_ ), .Z(_01781_ ) );
NAND2_X1 _22460_ ( .A1(_01781_ ), .A2(_01194_ ), .ZN(_01782_ ) );
INV_X1 _22461_ ( .A(_01583_ ), .ZN(_01783_ ) );
NAND2_X1 _22462_ ( .A1(_01783_ ), .A2(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01784_ ) );
NAND3_X1 _22463_ ( .A1(_01758_ ), .A2(_01759_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01785_ ) );
NAND2_X1 _22464_ ( .A1(_01784_ ), .A2(_01785_ ), .ZN(_01786_ ) );
OAI21_X1 _22465_ ( .A(_01782_ ), .B1(_01786_ ), .B2(_01781_ ), .ZN(_01787_ ) );
BUF_X4 _22466_ ( .A(_01590_ ), .Z(_01788_ ) );
INV_X1 _22467_ ( .A(_01204_ ), .ZN(_01789_ ) );
BUF_X4 _22468_ ( .A(_01789_ ), .Z(_01790_ ) );
NAND3_X1 _22469_ ( .A1(_01787_ ), .A2(_01788_ ), .A3(_01790_ ), .ZN(_01791_ ) );
AND2_X1 _22470_ ( .A1(_01780_ ), .A2(_01791_ ), .ZN(_01792_ ) );
INV_X1 _22471_ ( .A(_01210_ ), .ZN(_01793_ ) );
BUF_X4 _22472_ ( .A(_01793_ ), .Z(_01794_ ) );
BUF_X2 _22473_ ( .A(_01794_ ), .Z(_01795_ ) );
INV_X1 _22474_ ( .A(_01216_ ), .ZN(_01796_ ) );
BUF_X2 _22475_ ( .A(_01796_ ), .Z(_01797_ ) );
OR3_X1 _22476_ ( .A1(_01792_ ), .A2(_01795_ ), .A3(_01797_ ), .ZN(_01798_ ) );
OR3_X1 _22477_ ( .A1(_01231_ ), .A2(_01252_ ), .A3(_01235_ ), .ZN(_01799_ ) );
OAI21_X1 _22478_ ( .A(_01290_ ), .B1(_01247_ ), .B2(_01250_ ), .ZN(_01800_ ) );
OAI21_X1 _22479_ ( .A(_01235_ ), .B1(_01224_ ), .B2(_01228_ ), .ZN(_01801_ ) );
NAND2_X1 _22480_ ( .A1(_01800_ ), .A2(_01801_ ), .ZN(_01802_ ) );
OAI21_X1 _22481_ ( .A(_01799_ ), .B1(_01240_ ), .B2(_01802_ ), .ZN(_01803_ ) );
BUF_X2 _22482_ ( .A(_01331_ ), .Z(_01804_ ) );
NAND3_X1 _22483_ ( .A1(_01803_ ), .A2(_01804_ ), .A3(_01686_ ), .ZN(_01805_ ) );
OAI211_X1 _22484_ ( .A(_01253_ ), .B(_01322_ ), .C1(_01297_ ), .C2(_01323_ ), .ZN(_01806_ ) );
OAI211_X1 _22485_ ( .A(_01291_ ), .B(_01311_ ), .C1(_01273_ ), .C2(_01312_ ), .ZN(_01807_ ) );
NAND3_X1 _22486_ ( .A1(_01806_ ), .A2(_01807_ ), .A3(_01252_ ), .ZN(_01808_ ) );
OAI211_X1 _22487_ ( .A(_01235_ ), .B(_01276_ ), .C1(_01273_ ), .C2(_01277_ ), .ZN(_01809_ ) );
OAI211_X1 _22488_ ( .A(_01290_ ), .B(_01319_ ), .C1(_01273_ ), .C2(_01320_ ), .ZN(_01810_ ) );
NAND3_X1 _22489_ ( .A1(_01809_ ), .A2(_01810_ ), .A3(_01240_ ), .ZN(_01811_ ) );
NAND2_X1 _22490_ ( .A1(_01808_ ), .A2(_01811_ ), .ZN(_01812_ ) );
OAI211_X1 _22491_ ( .A(_01262_ ), .B(_01235_ ), .C1(_01263_ ), .C2(_01264_ ), .ZN(_01813_ ) );
OAI211_X1 _22492_ ( .A(_01291_ ), .B(_01272_ ), .C1(_01273_ ), .C2(_01274_ ), .ZN(_01814_ ) );
AOI21_X1 _22493_ ( .A(_01240_ ), .B1(_01813_ ), .B2(_01814_ ), .ZN(_01815_ ) );
OAI211_X1 _22494_ ( .A(_01290_ ), .B(_01266_ ), .C1(_01273_ ), .C2(_01267_ ), .ZN(_01816_ ) );
OAI21_X1 _22495_ ( .A(_01235_ ), .B1(_01256_ ), .B2(_01257_ ), .ZN(_01817_ ) );
AOI21_X1 _22496_ ( .A(_01252_ ), .B1(_01816_ ), .B2(_01817_ ), .ZN(_01818_ ) );
NOR2_X1 _22497_ ( .A1(_01815_ ), .A2(_01818_ ), .ZN(_01819_ ) );
MUX2_X1 _22498_ ( .A(_01812_ ), .B(_01819_ ), .S(_01308_ ), .Z(_01820_ ) );
OAI21_X1 _22499_ ( .A(_01805_ ), .B1(_01820_ ), .B2(_01804_ ), .ZN(_01821_ ) );
NAND2_X1 _22500_ ( .A1(_01821_ ), .A2(_01338_ ), .ZN(_01822_ ) );
BUF_X2 _22501_ ( .A(_01342_ ), .Z(_01823_ ) );
NAND2_X1 _22502_ ( .A1(_01392_ ), .A2(_01398_ ), .ZN(_01824_ ) );
INV_X1 _22503_ ( .A(_01407_ ), .ZN(_01825_ ) );
AOI21_X1 _22504_ ( .A(_01394_ ), .B1(_01824_ ), .B2(_01825_ ), .ZN(_01826_ ) );
OR3_X1 _22505_ ( .A1(_01826_ ), .A2(_08757_ ), .A3(_01411_ ), .ZN(_01827_ ) );
BUF_X2 _22506_ ( .A(_01436_ ), .Z(_01828_ ) );
OAI21_X1 _22507_ ( .A(_08757_ ), .B1(_01826_ ), .B2(_01411_ ), .ZN(_01829_ ) );
AND3_X1 _22508_ ( .A1(_01827_ ), .A2(_01828_ ), .A3(_01829_ ), .ZN(_01830_ ) );
NAND2_X1 _22509_ ( .A1(_01821_ ), .A2(_01441_ ), .ZN(_01831_ ) );
INV_X1 _22510_ ( .A(_01447_ ), .ZN(_01832_ ) );
NOR3_X1 _22511_ ( .A1(_01792_ ), .A2(_01795_ ), .A3(_01455_ ), .ZN(_01833_ ) );
NOR2_X1 _22512_ ( .A1(_08840_ ), .A2(_08865_ ), .ZN(_01834_ ) );
NOR4_X1 _22513_ ( .A1(_01834_ ), .A2(_08746_ ), .A3(_08748_ ), .A4(_08881_ ), .ZN(_01835_ ) );
OR3_X1 _22514_ ( .A1(_01835_ ), .A2(_08885_ ), .A3(_08883_ ), .ZN(_01836_ ) );
AND2_X1 _22515_ ( .A1(_01836_ ), .A2(_01394_ ), .ZN(_01837_ ) );
OR3_X1 _22516_ ( .A1(_01837_ ), .A2(_01395_ ), .A3(_08892_ ), .ZN(_01838_ ) );
OAI21_X1 _22517_ ( .A(_01395_ ), .B1(_01837_ ), .B2(_08892_ ), .ZN(_01839_ ) );
NAND3_X1 _22518_ ( .A1(_01838_ ), .A2(_01478_ ), .A3(_01839_ ), .ZN(_01840_ ) );
AND4_X1 _22519_ ( .A1(\exu.addi.io_imm [21] ), .A2(_01601_ ), .A3(_01602_ ), .A4(_01604_ ), .ZN(_01841_ ) );
AOI21_X1 _22520_ ( .A(_01841_ ), .B1(_09570_ ), .B2(_01607_ ), .ZN(_01842_ ) );
OAI21_X1 _22521_ ( .A(_01840_ ), .B1(_01842_ ), .B2(\exu.io_in_bits_sub ), .ZN(_01843_ ) );
AOI21_X1 _22522_ ( .A(_01833_ ), .B1(_01843_ ), .B2(_01610_ ), .ZN(_01844_ ) );
OAI221_X1 _22523_ ( .A(_01614_ ), .B1(_08756_ ), .B2(_01832_ ), .C1(_01844_ ), .C2(\exu.io_in_bits_or ), .ZN(_01845_ ) );
NOR2_X1 _22524_ ( .A1(_01750_ ), .A2(_01579_ ), .ZN(_01846_ ) );
OAI211_X1 _22525_ ( .A(_01845_ ), .B(_01486_ ), .C1(_01614_ ), .C2(_01846_ ), .ZN(_01847_ ) );
NAND3_X1 _22526_ ( .A1(_08755_ ), .A2(_10699_ ), .A3(fanout_net_4 ), .ZN(_01848_ ) );
AOI21_X1 _22527_ ( .A(\exu.io_in_bits_xor ), .B1(_01847_ ), .B2(_01848_ ), .ZN(_01849_ ) );
AOI21_X1 _22528_ ( .A(_01849_ ), .B1(_08757_ ), .B2(_01493_ ), .ZN(_01850_ ) );
OAI21_X1 _22529_ ( .A(_01831_ ), .B1(_01850_ ), .B2(fanout_net_12 ), .ZN(_01851_ ) );
AOI21_X1 _22530_ ( .A(_01830_ ), .B1(_01851_ ), .B2(_01498_ ), .ZN(_01852_ ) );
OAI221_X1 _22531_ ( .A(_01341_ ), .B1(_01823_ ), .B2(_09576_ ), .C1(_01852_ ), .C2(\exu.io_in_bits_jal ), .ZN(_01853_ ) );
BUF_X4 _22532_ ( .A(_01341_ ), .Z(_01854_ ) );
BUF_X2 _22533_ ( .A(_09177_ ), .Z(_01855_ ) );
NOR2_X1 _22534_ ( .A1(_09576_ ), .A2(_01855_ ), .ZN(_01856_ ) );
OAI211_X1 _22535_ ( .A(_01853_ ), .B(_01501_ ), .C1(_01854_ ), .C2(_01856_ ), .ZN(_01857_ ) );
MUX2_X1 _22536_ ( .A(_01822_ ), .B(_01857_ ), .S(_01505_ ), .Z(_01858_ ) );
MUX2_X1 _22537_ ( .A(_01798_ ), .B(_01858_ ), .S(_01705_ ), .Z(_01859_ ) );
BUF_X4 _22538_ ( .A(_01510_ ), .Z(_01860_ ) );
MUX2_X1 _22539_ ( .A(_01756_ ), .B(_01859_ ), .S(_01860_ ), .Z(_01861_ ) );
BUF_X4 _22540_ ( .A(_01182_ ), .Z(_01862_ ) );
AOI21_X1 _22541_ ( .A(_01754_ ), .B1(_01861_ ), .B2(_01862_ ), .ZN(_01863_ ) );
CLKBUF_X2 _22542_ ( .A(_10842_ ), .Z(_01864_ ) );
AND3_X1 _22543_ ( .A1(_09145_ ), .A2(_01864_ ), .A3(fanout_net_5 ), .ZN(_01865_ ) );
OAI21_X1 _22544_ ( .A(_01723_ ), .B1(_01863_ ), .B2(_01865_ ), .ZN(_01866_ ) );
BUF_X4 _22545_ ( .A(_01518_ ), .Z(_01867_ ) );
NAND2_X1 _22546_ ( .A1(_09147_ ), .A2(_01867_ ), .ZN(_01868_ ) );
AOI21_X1 _22547_ ( .A(_01722_ ), .B1(_01866_ ), .B2(_01868_ ), .ZN(_01869_ ) );
CLKBUF_X2 _22548_ ( .A(_01523_ ), .Z(_01870_ ) );
AND2_X1 _22549_ ( .A1(\exu.addi._io_rd_T_4 [21] ), .A2(_01870_ ), .ZN(_01871_ ) );
OAI21_X1 _22550_ ( .A(_01721_ ), .B1(_01869_ ), .B2(_01871_ ), .ZN(_01872_ ) );
BUF_X2 _22551_ ( .A(_10844_ ), .Z(_01873_ ) );
OAI211_X1 _22552_ ( .A(_01873_ ), .B(\exu.csrrs.io_csr_rdata [21] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_01874_ ) );
NAND2_X1 _22553_ ( .A1(_01872_ ), .A2(_01874_ ), .ZN(\exu.io_out_bits_rd_wdata [21] ) );
BUF_X4 _22554_ ( .A(_01109_ ), .Z(_01875_ ) );
BUF_X4 _22555_ ( .A(_01173_ ), .Z(_01876_ ) );
BUF_X4 _22556_ ( .A(_01175_ ), .Z(_01877_ ) );
BUF_X4 _22557_ ( .A(_01176_ ), .Z(_01878_ ) );
BUF_X4 _22558_ ( .A(_01533_ ), .Z(_01879_ ) );
BUF_X4 _22559_ ( .A(_01879_ ), .Z(_01880_ ) );
BUF_X4 _22560_ ( .A(_01564_ ), .Z(_01881_ ) );
BUF_X2 _22561_ ( .A(_01562_ ), .Z(_01882_ ) );
OR2_X1 _22562_ ( .A1(_01556_ ), .A2(_01666_ ), .ZN(_01883_ ) );
BUF_X4 _22563_ ( .A(_01725_ ), .Z(_01884_ ) );
INV_X1 _22564_ ( .A(_01556_ ), .ZN(_01885_ ) );
OAI211_X1 _22565_ ( .A(_01883_ ), .B(_01884_ ), .C1(_01315_ ), .C2(_01885_ ), .ZN(_01886_ ) );
BUF_X4 _22566_ ( .A(_01559_ ), .Z(_01887_ ) );
BUF_X4 _22567_ ( .A(_01887_ ), .Z(_01888_ ) );
NAND3_X1 _22568_ ( .A1(_01726_ ), .A2(_01727_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01889_ ) );
BUF_X4 _22569_ ( .A(_01729_ ), .Z(_01890_ ) );
BUF_X4 _22570_ ( .A(_01890_ ), .Z(_01891_ ) );
INV_X1 _22571_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01892_ ) );
OAI211_X1 _22572_ ( .A(_01888_ ), .B(_01889_ ), .C1(_01891_ ), .C2(_01892_ ), .ZN(_01893_ ) );
AOI21_X1 _22573_ ( .A(_01882_ ), .B1(_01886_ ), .B2(_01893_ ), .ZN(_01894_ ) );
AND3_X1 _22574_ ( .A1(_01726_ ), .A2(_01727_ ), .A3(_01675_ ), .ZN(_01895_ ) );
AOI21_X1 _22575_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_01726_ ), .B2(_01727_ ), .ZN(_01896_ ) );
NOR2_X1 _22576_ ( .A1(_01895_ ), .A2(_01896_ ), .ZN(_01897_ ) );
NAND2_X1 _22577_ ( .A1(_01897_ ), .A2(_01888_ ), .ZN(_01898_ ) );
BUF_X4 _22578_ ( .A(_01725_ ), .Z(_01899_ ) );
BUF_X2 _22579_ ( .A(_01553_ ), .Z(_01900_ ) );
BUF_X2 _22580_ ( .A(_01900_ ), .Z(_01901_ ) );
BUF_X2 _22581_ ( .A(_01554_ ), .Z(_01902_ ) );
BUF_X2 _22582_ ( .A(_01902_ ), .Z(_01903_ ) );
NAND3_X1 _22583_ ( .A1(_01901_ ), .A2(_01903_ ), .A3(_01293_ ), .ZN(_01904_ ) );
OAI211_X1 _22584_ ( .A(_01899_ ), .B(_01904_ ), .C1(_01891_ ), .C2(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01905_ ) );
AND3_X1 _22585_ ( .A1(_01898_ ), .A2(_01882_ ), .A3(_01905_ ), .ZN(_01906_ ) );
OAI21_X1 _22586_ ( .A(_01881_ ), .B1(_01894_ ), .B2(_01906_ ), .ZN(_01907_ ) );
OR2_X1 _22587_ ( .A1(_01729_ ), .A2(_01301_ ), .ZN(_01908_ ) );
NAND3_X1 _22588_ ( .A1(_01726_ ), .A2(_01727_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01909_ ) );
NAND2_X1 _22589_ ( .A1(_01908_ ), .A2(_01909_ ), .ZN(_01910_ ) );
MUX2_X1 _22590_ ( .A(_01910_ ), .B(_01557_ ), .S(_01899_ ), .Z(_01911_ ) );
MUX2_X1 _22591_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B ), .B(_01911_ ), .S(_01734_ ), .Z(_01912_ ) );
OAI211_X1 _22592_ ( .A(_01880_ ), .B(_01907_ ), .C1(_01912_ ), .C2(_01881_ ), .ZN(_01913_ ) );
BUF_X2 _22593_ ( .A(_01530_ ), .Z(_01914_ ) );
AND3_X1 _22594_ ( .A1(_01913_ ), .A2(_01914_ ), .A3(_01537_ ), .ZN(_01915_ ) );
OAI21_X1 _22595_ ( .A(_01878_ ), .B1(_01915_ ), .B2(_01512_ ), .ZN(_01916_ ) );
OAI21_X1 _22596_ ( .A(_01755_ ), .B1(\exu.add.io_rs1_data [20] ), .B2(\exu.addi.io_imm [20] ), .ZN(_01917_ ) );
AND3_X1 _22597_ ( .A1(_01190_ ), .A2(_01193_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01918_ ) );
AOI21_X1 _22598_ ( .A(_01735_ ), .B1(_01764_ ), .B2(_01765_ ), .ZN(_01919_ ) );
OR3_X1 _22599_ ( .A1(_01918_ ), .A2(_01919_ ), .A3(_01761_ ), .ZN(_01920_ ) );
AND3_X1 _22600_ ( .A1(_01764_ ), .A2(_01765_ ), .A3(_01675_ ), .ZN(_01921_ ) );
BUF_X2 _22601_ ( .A(_01190_ ), .Z(_01922_ ) );
BUF_X2 _22602_ ( .A(_01193_ ), .Z(_01923_ ) );
AOI21_X1 _22603_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_01922_ ), .B2(_01923_ ), .ZN(_01924_ ) );
OAI21_X1 _22604_ ( .A(_01761_ ), .B1(_01921_ ), .B2(_01924_ ), .ZN(_01925_ ) );
AOI21_X1 _22605_ ( .A(_01788_ ), .B1(_01920_ ), .B2(_01925_ ), .ZN(_01926_ ) );
BUF_X2 _22606_ ( .A(_01771_ ), .Z(_01927_ ) );
AND3_X1 _22607_ ( .A1(_01922_ ), .A2(_01923_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01928_ ) );
AOI21_X1 _22608_ ( .A(_01666_ ), .B1(_01922_ ), .B2(_01923_ ), .ZN(_01929_ ) );
OR3_X1 _22609_ ( .A1(_01928_ ), .A2(_01929_ ), .A3(_01761_ ), .ZN(_01930_ ) );
NAND3_X1 _22610_ ( .A1(_01922_ ), .A2(_01923_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01931_ ) );
OAI211_X1 _22611_ ( .A(_01763_ ), .B(_01931_ ), .C1(_01767_ ), .C2(_01892_ ), .ZN(_01932_ ) );
AOI21_X1 _22612_ ( .A(_01927_ ), .B1(_01930_ ), .B2(_01932_ ), .ZN(_01933_ ) );
NOR2_X1 _22613_ ( .A1(_01926_ ), .A2(_01933_ ), .ZN(_01934_ ) );
BUF_X4 _22614_ ( .A(_01790_ ), .Z(_01935_ ) );
NOR2_X1 _22615_ ( .A1(_01934_ ), .A2(_01935_ ), .ZN(_01936_ ) );
AND3_X1 _22616_ ( .A1(_01190_ ), .A2(_01193_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01937_ ) );
AOI21_X1 _22617_ ( .A(_01301_ ), .B1(_01764_ ), .B2(_01765_ ), .ZN(_01938_ ) );
OR2_X1 _22618_ ( .A1(_01937_ ), .A2(_01938_ ), .ZN(_01939_ ) );
MUX2_X1 _22619_ ( .A(_01939_ ), .B(_01584_ ), .S(_01586_ ), .Z(_01940_ ) );
NOR2_X1 _22620_ ( .A1(_01940_ ), .A2(_01927_ ), .ZN(_01941_ ) );
AOI21_X1 _22621_ ( .A(_01936_ ), .B1(_01941_ ), .B2(_01935_ ), .ZN(_01942_ ) );
OR3_X1 _22622_ ( .A1(_01942_ ), .A2(_01795_ ), .A3(_01797_ ), .ZN(_01943_ ) );
AND2_X1 _22623_ ( .A1(_01291_ ), .A2(_01634_ ), .ZN(_01944_ ) );
INV_X1 _22624_ ( .A(_01944_ ), .ZN(_01945_ ) );
NAND2_X1 _22625_ ( .A1(_01622_ ), .A2(_01299_ ), .ZN(_01946_ ) );
NAND2_X1 _22626_ ( .A1(_01632_ ), .A2(_01253_ ), .ZN(_01947_ ) );
NAND2_X1 _22627_ ( .A1(_01946_ ), .A2(_01947_ ), .ZN(_01948_ ) );
MUX2_X1 _22628_ ( .A(_01945_ ), .B(_01948_ ), .S(_01279_ ), .Z(_01949_ ) );
OR3_X1 _22629_ ( .A1(_01949_ ), .A2(_01333_ ), .A3(_01308_ ), .ZN(_01950_ ) );
OAI21_X1 _22630_ ( .A(_01299_ ), .B1(_01647_ ), .B2(_01649_ ), .ZN(_01951_ ) );
OAI21_X1 _22631_ ( .A(_01254_ ), .B1(_01624_ ), .B2(_01625_ ), .ZN(_01952_ ) );
AND3_X1 _22632_ ( .A1(_01951_ ), .A2(_01952_ ), .A3(_01241_ ), .ZN(_01953_ ) );
OAI211_X1 _22633_ ( .A(_01253_ ), .B(_01645_ ), .C1(_01297_ ), .C2(_01263_ ), .ZN(_01954_ ) );
OAI211_X1 _22634_ ( .A(_01291_ ), .B(_01641_ ), .C1(_01297_ ), .C2(_01642_ ), .ZN(_01955_ ) );
AOI21_X1 _22635_ ( .A(_01241_ ), .B1(_01954_ ), .B2(_01955_ ), .ZN(_01956_ ) );
NOR2_X1 _22636_ ( .A1(_01953_ ), .A2(_01956_ ), .ZN(_01957_ ) );
OAI211_X1 _22637_ ( .A(_01639_ ), .B(_01253_ ), .C1(_01274_ ), .C2(_01264_ ), .ZN(_01958_ ) );
OR3_X1 _22638_ ( .A1(_01660_ ), .A2(_01662_ ), .A3(_01253_ ), .ZN(_01959_ ) );
AOI21_X1 _22639_ ( .A(_01306_ ), .B1(_01958_ ), .B2(_01959_ ), .ZN(_01960_ ) );
OR3_X1 _22640_ ( .A1(_01668_ ), .A2(_01669_ ), .A3(_01253_ ), .ZN(_01961_ ) );
OAI21_X1 _22641_ ( .A(_01253_ ), .B1(_01656_ ), .B2(_01658_ ), .ZN(_01962_ ) );
AND3_X1 _22642_ ( .A1(_01961_ ), .A2(_01962_ ), .A3(_01279_ ), .ZN(_01963_ ) );
NOR2_X1 _22643_ ( .A1(_01960_ ), .A2(_01963_ ), .ZN(_01964_ ) );
MUX2_X1 _22644_ ( .A(_01957_ ), .B(_01964_ ), .S(_01686_ ), .Z(_01965_ ) );
OAI21_X1 _22645_ ( .A(_01950_ ), .B1(_01965_ ), .B2(_01654_ ), .ZN(_01966_ ) );
NAND2_X1 _22646_ ( .A1(_01966_ ), .A2(_01702_ ), .ZN(_01967_ ) );
BUF_X4 _22647_ ( .A(_01492_ ), .Z(_01968_ ) );
NAND3_X1 _22648_ ( .A1(_01411_ ), .A2(_01575_ ), .A3(fanout_net_4 ), .ZN(_01969_ ) );
AND3_X1 _22649_ ( .A1(_01913_ ), .A2(_01445_ ), .A3(_01536_ ), .ZN(_01970_ ) );
OAI21_X1 _22650_ ( .A(_01581_ ), .B1(\exu.add.io_rs1_data [20] ), .B2(\exu._GEN_0 [20] ), .ZN(_01971_ ) );
NOR3_X1 _22651_ ( .A1(_01942_ ), .A2(_01794_ ), .A3(_01455_ ), .ZN(_01972_ ) );
AOI21_X1 _22652_ ( .A(_01597_ ), .B1(_01836_ ), .B2(_01394_ ), .ZN(_01973_ ) );
OAI21_X1 _22653_ ( .A(_01973_ ), .B1(_01394_ ), .B2(_01836_ ), .ZN(_01974_ ) );
AND4_X1 _22654_ ( .A1(\exu.addi.io_imm [20] ), .A2(_01600_ ), .A3(_01463_ ), .A4(_01603_ ), .ZN(_01975_ ) );
AOI21_X1 _22655_ ( .A(_01975_ ), .B1(_10018_ ), .B2(_01607_ ), .ZN(_01976_ ) );
OAI21_X1 _22656_ ( .A(_01974_ ), .B1(_01976_ ), .B2(\exu.io_in_bits_sub ), .ZN(_01977_ ) );
AOI21_X1 _22657_ ( .A(_01972_ ), .B1(_01977_ ), .B2(_01610_ ), .ZN(_01978_ ) );
OAI21_X1 _22658_ ( .A(_01971_ ), .B1(_01978_ ), .B2(\exu.io_in_bits_or ), .ZN(_01979_ ) );
AOI21_X1 _22659_ ( .A(_01970_ ), .B1(_01979_ ), .B2(_01614_ ), .ZN(_01980_ ) );
OAI21_X1 _22660_ ( .A(_01969_ ), .B1(_01980_ ), .B2(fanout_net_4 ), .ZN(_01981_ ) );
AOI221_X4 _22661_ ( .A(fanout_net_12 ), .B1(_08754_ ), .B2(_01968_ ), .C1(_01981_ ), .C2(_01618_ ), .ZN(_01982_ ) );
NAND2_X1 _22662_ ( .A1(_01966_ ), .A2(_01689_ ), .ZN(_01983_ ) );
AOI211_X1 _22663_ ( .A(_01574_ ), .B(_01982_ ), .C1(fanout_net_12 ), .C2(_01983_ ), .ZN(_01984_ ) );
NAND3_X1 _22664_ ( .A1(_01824_ ), .A2(_01394_ ), .A3(_01825_ ), .ZN(_01985_ ) );
NOR2_X1 _22665_ ( .A1(_01826_ ), .A2(_01694_ ), .ZN(_01986_ ) );
AOI21_X1 _22666_ ( .A(_01984_ ), .B1(_01985_ ), .B2(_01986_ ), .ZN(_01987_ ) );
OAI221_X1 _22667_ ( .A(_01341_ ), .B1(_01823_ ), .B2(_10031_ ), .C1(_01987_ ), .C2(\exu.io_in_bits_jal ), .ZN(_01988_ ) );
BUF_X4 _22668_ ( .A(_01501_ ), .Z(_01989_ ) );
AND2_X1 _22669_ ( .A1(_10020_ ), .A2(_01699_ ), .ZN(_01990_ ) );
OAI211_X1 _22670_ ( .A(_01988_ ), .B(_01989_ ), .C1(_01854_ ), .C2(_01990_ ), .ZN(_01991_ ) );
BUF_X4 _22671_ ( .A(_01505_ ), .Z(_01992_ ) );
MUX2_X1 _22672_ ( .A(_01967_ ), .B(_01991_ ), .S(_01992_ ), .Z(_01993_ ) );
BUF_X4 _22673_ ( .A(_01507_ ), .Z(_01994_ ) );
MUX2_X1 _22674_ ( .A(_01943_ ), .B(_01993_ ), .S(_01994_ ), .Z(_01995_ ) );
MUX2_X1 _22675_ ( .A(_01917_ ), .B(_01995_ ), .S(_01860_ ), .Z(_01996_ ) );
AOI21_X1 _22676_ ( .A(_01916_ ), .B1(_01996_ ), .B2(_01862_ ), .ZN(_01997_ ) );
AND3_X1 _22677_ ( .A1(_09148_ ), .A2(_10844_ ), .A3(fanout_net_5 ), .ZN(_01998_ ) );
OAI21_X1 _22678_ ( .A(_01877_ ), .B1(_01997_ ), .B2(_01998_ ), .ZN(_01999_ ) );
BUF_X4 _22679_ ( .A(_01519_ ), .Z(_02000_ ) );
NAND2_X1 _22680_ ( .A1(_09150_ ), .A2(_02000_ ), .ZN(_02001_ ) );
AOI21_X1 _22681_ ( .A(_01876_ ), .B1(_01999_ ), .B2(_02001_ ), .ZN(_02002_ ) );
CLKBUF_X2 _22682_ ( .A(_01523_ ), .Z(_02003_ ) );
AND2_X1 _22683_ ( .A1(\exu.addi._io_rd_T_4 [20] ), .A2(_02003_ ), .ZN(_02004_ ) );
OAI21_X1 _22684_ ( .A(_01875_ ), .B1(_02002_ ), .B2(_02004_ ), .ZN(_02005_ ) );
OAI211_X1 _22685_ ( .A(_01058_ ), .B(\exu.csrrs.io_csr_rdata [20] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_02006_ ) );
NAND2_X1 _22686_ ( .A1(_02005_ ), .A2(_02006_ ), .ZN(\exu.io_out_bits_rd_wdata [20] ) );
AND3_X1 _22687_ ( .A1(_09043_ ), .A2(_10842_ ), .A3(fanout_net_5 ), .ZN(_02007_ ) );
NAND3_X1 _22688_ ( .A1(_01726_ ), .A2(_01727_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02008_ ) );
OAI211_X1 _22689_ ( .A(_01725_ ), .B(_02008_ ), .C1(_01556_ ), .C2(_01675_ ), .ZN(_02009_ ) );
OAI211_X1 _22690_ ( .A(_01558_ ), .B(_01728_ ), .C1(_01556_ ), .C2(_01315_ ), .ZN(_02010_ ) );
AOI21_X1 _22691_ ( .A(_01545_ ), .B1(_02009_ ), .B2(_02010_ ), .ZN(_02011_ ) );
OAI211_X1 _22692_ ( .A(_01724_ ), .B(_01731_ ), .C1(_01556_ ), .C2(_01312_ ), .ZN(_02012_ ) );
NAND3_X1 _22693_ ( .A1(_01553_ ), .A2(_01554_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02013_ ) );
OAI211_X1 _22694_ ( .A(_01558_ ), .B(_02013_ ), .C1(_01556_ ), .C2(_01323_ ), .ZN(_02014_ ) );
AOI21_X1 _22695_ ( .A(_01561_ ), .B1(_02012_ ), .B2(_02014_ ), .ZN(_02015_ ) );
NOR2_X1 _22696_ ( .A1(_02011_ ), .A2(_02015_ ), .ZN(_02016_ ) );
OR2_X1 _22697_ ( .A1(_01738_ ), .A2(_01739_ ), .ZN(_02017_ ) );
MUX2_X1 _22698_ ( .A(_02017_ ), .B(_01743_ ), .S(_01724_ ), .Z(_02018_ ) );
MUX2_X1 _22699_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B ), .B(_02018_ ), .S(_01545_ ), .Z(_02019_ ) );
MUX2_X1 _22700_ ( .A(_02016_ ), .B(_02019_ ), .S(_01746_ ), .Z(_02020_ ) );
BUF_X4 _22701_ ( .A(_01880_ ), .Z(_02021_ ) );
AOI211_X1 _22702_ ( .A(_01751_ ), .B(_01534_ ), .C1(_02020_ ), .C2(_02021_ ), .ZN(_02022_ ) );
BUF_X4 _22703_ ( .A(_01184_ ), .Z(_02023_ ) );
NOR3_X1 _22704_ ( .A1(_09044_ ), .A2(fanout_net_26 ), .A3(_02023_ ), .ZN(_02024_ ) );
OAI211_X1 _22705_ ( .A(_01586_ ), .B(_01766_ ), .C1(_01583_ ), .C2(_01312_ ), .ZN(_02025_ ) );
AND3_X1 _22706_ ( .A1(_01190_ ), .A2(_01193_ ), .A3(_01892_ ), .ZN(_02026_ ) );
AOI21_X1 _22707_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_01190_ ), .B2(_01193_ ), .ZN(_02027_ ) );
OAI21_X1 _22708_ ( .A(_01197_ ), .B1(_02026_ ), .B2(_02027_ ), .ZN(_02028_ ) );
NAND2_X1 _22709_ ( .A1(_02025_ ), .A2(_02028_ ), .ZN(_02029_ ) );
NAND2_X1 _22710_ ( .A1(_02029_ ), .A2(_01200_ ), .ZN(_02030_ ) );
NOR2_X1 _22711_ ( .A1(_01772_ ), .A2(_01773_ ), .ZN(_02031_ ) );
NAND2_X1 _22712_ ( .A1(_02031_ ), .A2(_01585_ ), .ZN(_02032_ ) );
OAI21_X1 _22713_ ( .A(_01197_ ), .B1(_01757_ ), .B2(_01760_ ), .ZN(_02033_ ) );
NAND3_X1 _22714_ ( .A1(_02032_ ), .A2(_01770_ ), .A3(_02033_ ), .ZN(_02034_ ) );
AOI21_X1 _22715_ ( .A(_01789_ ), .B1(_02030_ ), .B2(_02034_ ), .ZN(_02035_ ) );
NAND3_X1 _22716_ ( .A1(_01770_ ), .A2(_01194_ ), .A3(_01763_ ), .ZN(_02036_ ) );
NAND2_X1 _22717_ ( .A1(_01786_ ), .A2(_01585_ ), .ZN(_02037_ ) );
OAI21_X1 _22718_ ( .A(_01197_ ), .B1(_01775_ ), .B2(_01776_ ), .ZN(_02038_ ) );
NAND2_X1 _22719_ ( .A1(_02037_ ), .A2(_02038_ ), .ZN(_02039_ ) );
OAI21_X1 _22720_ ( .A(_02036_ ), .B1(_02039_ ), .B2(_01770_ ), .ZN(_02040_ ) );
AOI21_X1 _22721_ ( .A(_02035_ ), .B1(_02040_ ), .B2(_01789_ ), .ZN(_02041_ ) );
NOR3_X1 _22722_ ( .A1(_02041_ ), .A2(_01795_ ), .A3(_01796_ ), .ZN(_02042_ ) );
NOR3_X1 _22723_ ( .A1(_01236_ ), .A2(_01245_ ), .A3(_01240_ ), .ZN(_02043_ ) );
NAND3_X1 _22724_ ( .A1(_01321_ ), .A2(_01324_ ), .A3(_01252_ ), .ZN(_02044_ ) );
NAND3_X1 _22725_ ( .A1(_01275_ ), .A2(_01278_ ), .A3(_01240_ ), .ZN(_02045_ ) );
AND2_X1 _22726_ ( .A1(_02044_ ), .A2(_02045_ ), .ZN(_02046_ ) );
AOI21_X1 _22727_ ( .A(_01239_ ), .B1(_01265_ ), .B2(_01268_ ), .ZN(_02047_ ) );
OAI21_X1 _22728_ ( .A(_01290_ ), .B1(_01256_ ), .B2(_01257_ ), .ZN(_02048_ ) );
AOI21_X1 _22729_ ( .A(_01252_ ), .B1(_01251_ ), .B2(_02048_ ), .ZN(_02049_ ) );
OR2_X1 _22730_ ( .A1(_02047_ ), .A2(_02049_ ), .ZN(_02050_ ) );
MUX2_X1 _22731_ ( .A(_02046_ ), .B(_02050_ ), .S(_01245_ ), .Z(_02051_ ) );
MUX2_X1 _22732_ ( .A(_02043_ ), .B(_02051_ ), .S(_01332_ ), .Z(_02052_ ) );
AND2_X1 _22733_ ( .A1(_02052_ ), .A2(_01337_ ), .ZN(_02053_ ) );
NAND3_X1 _22734_ ( .A1(_01400_ ), .A2(_09462_ ), .A3(fanout_net_4 ), .ZN(_02054_ ) );
NAND2_X1 _22735_ ( .A1(_02020_ ), .A2(_01533_ ), .ZN(_02055_ ) );
AND3_X1 _22736_ ( .A1(_02055_ ), .A2(_01444_ ), .A3(_01535_ ), .ZN(_02056_ ) );
OAI21_X1 _22737_ ( .A(_01447_ ), .B1(\exu.add.io_rs1_data [19] ), .B2(\exu._GEN_0 [19] ), .ZN(_02057_ ) );
NOR3_X1 _22738_ ( .A1(_02041_ ), .A2(_01793_ ), .A3(_01454_ ), .ZN(_02058_ ) );
AND2_X1 _22739_ ( .A1(_09926_ ), .A2(_01459_ ), .ZN(_02059_ ) );
AND4_X1 _22740_ ( .A1(\exu.addi.io_imm [19] ), .A2(_01464_ ), .A3(_01458_ ), .A4(_01466_ ), .ZN(_02060_ ) );
OAI21_X1 _22741_ ( .A(_01457_ ), .B1(_02059_ ), .B2(_02060_ ), .ZN(_02061_ ) );
NOR2_X1 _22742_ ( .A1(_01834_ ), .A2(_08748_ ), .ZN(_02062_ ) );
AND2_X1 _22743_ ( .A1(_02062_ ), .A2(_08747_ ), .ZN(_02063_ ) );
INV_X1 _22744_ ( .A(_02063_ ), .ZN(_02064_ ) );
AOI21_X1 _22745_ ( .A(_08744_ ), .B1(_02064_ ), .B2(_08880_ ), .ZN(_02065_ ) );
AOI21_X1 _22746_ ( .A(_02065_ ), .B1(\exu.add.io_rs1_data [18] ), .B2(_01083_ ), .ZN(_02066_ ) );
XNOR2_X1 _22747_ ( .A(_02066_ ), .B(_08743_ ), .ZN(_02067_ ) );
OAI21_X1 _22748_ ( .A(_02061_ ), .B1(_01596_ ), .B2(_02067_ ), .ZN(_02068_ ) );
AOI21_X1 _22749_ ( .A(_02058_ ), .B1(_02068_ ), .B2(_01452_ ), .ZN(_02069_ ) );
OAI21_X1 _22750_ ( .A(_02057_ ), .B1(_02069_ ), .B2(\exu.io_in_bits_or ), .ZN(_02070_ ) );
AOI21_X1 _22751_ ( .A(_02056_ ), .B1(_02070_ ), .B2(_01443_ ), .ZN(_02071_ ) );
OAI21_X1 _22752_ ( .A(_02054_ ), .B1(_02071_ ), .B2(fanout_net_4 ), .ZN(_02072_ ) );
AOI221_X4 _22753_ ( .A(fanout_net_12 ), .B1(_08743_ ), .B2(_01491_ ), .C1(_02072_ ), .C2(_01490_ ), .ZN(_02073_ ) );
NAND2_X1 _22754_ ( .A1(_02052_ ), .A2(_01439_ ), .ZN(_02074_ ) );
AOI211_X1 _22755_ ( .A(_01572_ ), .B(_02073_ ), .C1(fanout_net_12 ), .C2(_02074_ ), .ZN(_02075_ ) );
INV_X1 _22756_ ( .A(_01401_ ), .ZN(_02076_ ) );
OR2_X1 _22757_ ( .A1(_01391_ ), .A2(_08749_ ), .ZN(_02077_ ) );
INV_X1 _22758_ ( .A(_01405_ ), .ZN(_02078_ ) );
AOI21_X1 _22759_ ( .A(_08747_ ), .B1(_02077_ ), .B2(_02078_ ), .ZN(_02079_ ) );
NOR2_X1 _22760_ ( .A1(_02079_ ), .A2(_01404_ ), .ZN(_02080_ ) );
INV_X1 _22761_ ( .A(_08744_ ), .ZN(_02081_ ) );
OAI21_X1 _22762_ ( .A(_02076_ ), .B1(_02080_ ), .B2(_02081_ ), .ZN(_02082_ ) );
XOR2_X1 _22763_ ( .A(_02082_ ), .B(_08743_ ), .Z(_02083_ ) );
AOI21_X1 _22764_ ( .A(_02075_ ), .B1(_01436_ ), .B2(_02083_ ), .ZN(_02084_ ) );
OR2_X1 _22765_ ( .A1(_02084_ ), .A2(\exu.io_in_bits_jal ), .ZN(_02085_ ) );
OAI21_X1 _22766_ ( .A(_02085_ ), .B1(_09999_ ), .B2(_09929_ ), .ZN(_02086_ ) );
NAND2_X1 _22767_ ( .A1(_02086_ ), .A2(_01340_ ), .ZN(_02087_ ) );
OR2_X1 _22768_ ( .A1(_09929_ ), .A2(_09177_ ), .ZN(_02088_ ) );
AOI21_X1 _22769_ ( .A(_10821_ ), .B1(_02087_ ), .B2(_02088_ ), .ZN(_02089_ ) );
MUX2_X1 _22770_ ( .A(_02053_ ), .B(_02089_ ), .S(_01504_ ), .Z(_02090_ ) );
MUX2_X1 _22771_ ( .A(_02042_ ), .B(_02090_ ), .S(_01214_ ), .Z(_02091_ ) );
MUX2_X1 _22772_ ( .A(_02024_ ), .B(_02091_ ), .S(_02023_ ), .Z(_02092_ ) );
MUX2_X1 _22773_ ( .A(_02022_ ), .B(_02092_ ), .S(_01181_ ), .Z(_02093_ ) );
MUX2_X1 _22774_ ( .A(_02007_ ), .B(_02093_ ), .S(_01515_ ), .Z(_02094_ ) );
AND2_X1 _22775_ ( .A1(_02094_ ), .A2(_01175_ ), .ZN(_02095_ ) );
INV_X1 _22776_ ( .A(_01518_ ), .ZN(_02096_ ) );
NOR3_X1 _22777_ ( .A1(_02096_ ), .A2(_09043_ ), .A3(_09044_ ), .ZN(_02097_ ) );
OAI21_X1 _22778_ ( .A(_01171_ ), .B1(_02095_ ), .B2(_02097_ ), .ZN(_02098_ ) );
NAND2_X1 _22779_ ( .A1(\exu.addi._io_rd_T_4 [19] ), .A2(_02003_ ), .ZN(_02099_ ) );
AOI21_X1 _22780_ ( .A(_01718_ ), .B1(_02098_ ), .B2(_02099_ ), .ZN(_02100_ ) );
AND3_X1 _22781_ ( .A1(_01718_ ), .A2(_01873_ ), .A3(\exu.csrrs.io_csr_rdata [19] ), .ZN(_02101_ ) );
OR2_X1 _22782_ ( .A1(_02100_ ), .A2(_02101_ ), .ZN(\exu.io_out_bits_rd_wdata [19] ) );
AND3_X1 _22783_ ( .A1(_09046_ ), .A2(_10699_ ), .A3(fanout_net_5 ), .ZN(_02102_ ) );
OAI211_X1 _22784_ ( .A(_01883_ ), .B(_01559_ ), .C1(_01315_ ), .C2(_01885_ ), .ZN(_02103_ ) );
OAI211_X1 _22785_ ( .A(_01561_ ), .B(_02103_ ), .C1(_01897_ ), .C2(_01559_ ), .ZN(_02104_ ) );
OAI211_X1 _22786_ ( .A(_01725_ ), .B(_01889_ ), .C1(_01729_ ), .C2(_01892_ ), .ZN(_02105_ ) );
AND3_X1 _22787_ ( .A1(_01553_ ), .A2(_01554_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02106_ ) );
AOI21_X1 _22788_ ( .A(_01657_ ), .B1(_01553_ ), .B2(_01554_ ), .ZN(_02107_ ) );
OR2_X1 _22789_ ( .A1(_02106_ ), .A2(_02107_ ), .ZN(_02108_ ) );
OAI211_X1 _22790_ ( .A(_01545_ ), .B(_02105_ ), .C1(_02108_ ), .C2(_01725_ ), .ZN(_02109_ ) );
NAND2_X1 _22791_ ( .A1(_02104_ ), .A2(_02109_ ), .ZN(_02110_ ) );
OAI211_X1 _22792_ ( .A(_01725_ ), .B(_01909_ ), .C1(_01729_ ), .C2(_01301_ ), .ZN(_02111_ ) );
NAND3_X1 _22793_ ( .A1(_01726_ ), .A2(_01727_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02112_ ) );
OAI211_X1 _22794_ ( .A(_01559_ ), .B(_02112_ ), .C1(_01729_ ), .C2(_01735_ ), .ZN(_02113_ ) );
NAND3_X1 _22795_ ( .A1(_02111_ ), .A2(_02113_ ), .A3(_01546_ ), .ZN(_02114_ ) );
OAI21_X1 _22796_ ( .A(_02114_ ), .B1(_01560_ ), .B2(_01546_ ), .ZN(_02115_ ) );
MUX2_X1 _22797_ ( .A(_02110_ ), .B(_02115_ ), .S(_01746_ ), .Z(_02116_ ) );
AOI211_X1 _22798_ ( .A(_01751_ ), .B(_01534_ ), .C1(_02116_ ), .C2(_02021_ ), .ZN(_02117_ ) );
NOR3_X1 _22799_ ( .A1(_09047_ ), .A2(fanout_net_26 ), .A3(_01184_ ), .ZN(_02118_ ) );
AND3_X1 _22800_ ( .A1(_01764_ ), .A2(_01765_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02119_ ) );
AOI21_X1 _22801_ ( .A(_01657_ ), .B1(_01764_ ), .B2(_01765_ ), .ZN(_02120_ ) );
OR3_X1 _22802_ ( .A1(_02119_ ), .A2(_01586_ ), .A3(_02120_ ), .ZN(_02121_ ) );
OAI211_X1 _22803_ ( .A(_01586_ ), .B(_01931_ ), .C1(_01767_ ), .C2(_01892_ ), .ZN(_02122_ ) );
AND3_X1 _22804_ ( .A1(_02121_ ), .A2(_01589_ ), .A3(_02122_ ), .ZN(_02123_ ) );
OR3_X1 _22805_ ( .A1(_01921_ ), .A2(_01924_ ), .A3(_01761_ ), .ZN(_02124_ ) );
OAI21_X1 _22806_ ( .A(_01761_ ), .B1(_01928_ ), .B2(_01929_ ), .ZN(_02125_ ) );
AOI21_X1 _22807_ ( .A(_01589_ ), .B1(_02124_ ), .B2(_02125_ ), .ZN(_02126_ ) );
OAI21_X1 _22808_ ( .A(_01591_ ), .B1(_02123_ ), .B2(_02126_ ), .ZN(_02127_ ) );
OR3_X1 _22809_ ( .A1(_01584_ ), .A2(_01781_ ), .A3(_01200_ ), .ZN(_02128_ ) );
OAI21_X1 _22810_ ( .A(_01781_ ), .B1(_01937_ ), .B2(_01938_ ), .ZN(_02129_ ) );
OAI21_X1 _22811_ ( .A(_01761_ ), .B1(_01918_ ), .B2(_01919_ ), .ZN(_02130_ ) );
NAND3_X1 _22812_ ( .A1(_02129_ ), .A2(_02130_ ), .A3(_01589_ ), .ZN(_02131_ ) );
NAND2_X1 _22813_ ( .A1(_02128_ ), .A2(_02131_ ), .ZN(_02132_ ) );
OAI21_X1 _22814_ ( .A(_02127_ ), .B1(_02132_ ), .B2(_01591_ ), .ZN(_02133_ ) );
NOR3_X1 _22815_ ( .A1(_02133_ ), .A2(_01795_ ), .A3(_01796_ ), .ZN(_02134_ ) );
NOR3_X1 _22816_ ( .A1(_01635_ ), .A2(_01245_ ), .A3(_01240_ ), .ZN(_02135_ ) );
AND3_X1 _22817_ ( .A1(_01640_ ), .A2(_01239_ ), .A3(_01643_ ), .ZN(_02136_ ) );
AOI21_X1 _22818_ ( .A(_01239_ ), .B1(_01659_ ), .B2(_01663_ ), .ZN(_02137_ ) );
OR2_X1 _22819_ ( .A1(_02136_ ), .A2(_02137_ ), .ZN(_02138_ ) );
AND2_X1 _22820_ ( .A1(_02138_ ), .A2(_01270_ ), .ZN(_02139_ ) );
NAND2_X1 _22821_ ( .A1(_01627_ ), .A2(_01240_ ), .ZN(_02140_ ) );
OAI211_X1 _22822_ ( .A(_01252_ ), .B(_01646_ ), .C1(_01650_ ), .C2(_01291_ ), .ZN(_02141_ ) );
NAND2_X1 _22823_ ( .A1(_02140_ ), .A2(_02141_ ), .ZN(_02142_ ) );
AOI21_X1 _22824_ ( .A(_02139_ ), .B1(_01245_ ), .B2(_02142_ ), .ZN(_02143_ ) );
MUX2_X1 _22825_ ( .A(_02135_ ), .B(_02143_ ), .S(_01332_ ), .Z(_02144_ ) );
AND2_X1 _22826_ ( .A1(_02144_ ), .A2(_01336_ ), .ZN(_02145_ ) );
NAND3_X1 _22827_ ( .A1(_01401_ ), .A2(_09462_ ), .A3(fanout_net_4 ), .ZN(_02146_ ) );
NAND2_X1 _22828_ ( .A1(_02116_ ), .A2(_01533_ ), .ZN(_02147_ ) );
AND3_X1 _22829_ ( .A1(_02147_ ), .A2(_01444_ ), .A3(_01535_ ), .ZN(_02148_ ) );
OAI21_X1 _22830_ ( .A(_01447_ ), .B1(\exu.add.io_rs1_data [18] ), .B2(\exu._GEN_0 [18] ), .ZN(_02149_ ) );
NOR3_X1 _22831_ ( .A1(_02133_ ), .A2(_01793_ ), .A3(_01454_ ), .ZN(_02150_ ) );
AND3_X1 _22832_ ( .A1(_02064_ ), .A2(_08744_ ), .A3(_08880_ ), .ZN(_02151_ ) );
OR3_X1 _22833_ ( .A1(_02151_ ), .A2(_02065_ ), .A3(_01596_ ), .ZN(_02152_ ) );
AND4_X1 _22834_ ( .A1(\exu.addi.io_imm [18] ), .A2(_01464_ ), .A3(_01458_ ), .A4(_01466_ ), .ZN(_02153_ ) );
AOI21_X1 _22835_ ( .A(_02153_ ), .B1(_09972_ ), .B2(_01459_ ), .ZN(_02154_ ) );
OAI21_X1 _22836_ ( .A(_02152_ ), .B1(_02154_ ), .B2(\exu.io_in_bits_sub ), .ZN(_02155_ ) );
AOI21_X1 _22837_ ( .A(_02150_ ), .B1(_02155_ ), .B2(_01452_ ), .ZN(_02156_ ) );
OAI21_X1 _22838_ ( .A(_02149_ ), .B1(_02156_ ), .B2(\exu.io_in_bits_or ), .ZN(_02157_ ) );
AOI21_X1 _22839_ ( .A(_02148_ ), .B1(_02157_ ), .B2(_01443_ ), .ZN(_02158_ ) );
OAI21_X1 _22840_ ( .A(_02146_ ), .B1(_02158_ ), .B2(fanout_net_4 ), .ZN(_02159_ ) );
AOI221_X4 _22841_ ( .A(fanout_net_12 ), .B1(_08744_ ), .B2(_01491_ ), .C1(_02159_ ), .C2(_01490_ ), .ZN(_02160_ ) );
NAND2_X1 _22842_ ( .A1(_02144_ ), .A2(_01439_ ), .ZN(_02161_ ) );
AOI211_X1 _22843_ ( .A(_01572_ ), .B(_02160_ ), .C1(fanout_net_12 ), .C2(_02161_ ), .ZN(_02162_ ) );
OAI21_X1 _22844_ ( .A(_01435_ ), .B1(_02080_ ), .B2(_02081_ ), .ZN(_02163_ ) );
AOI21_X1 _22845_ ( .A(_02163_ ), .B1(_02081_ ), .B2(_02080_ ), .ZN(_02164_ ) );
OAI21_X1 _22846_ ( .A(_09410_ ), .B1(_02162_ ), .B2(_02164_ ), .ZN(_02165_ ) );
OAI21_X1 _22847_ ( .A(_02165_ ), .B1(_09999_ ), .B2(_09976_ ), .ZN(_02166_ ) );
NAND2_X1 _22848_ ( .A1(_02166_ ), .A2(_09657_ ), .ZN(_02167_ ) );
NAND2_X1 _22849_ ( .A1(_09975_ ), .A2(_09460_ ), .ZN(_02168_ ) );
AOI21_X1 _22850_ ( .A(_10821_ ), .B1(_02167_ ), .B2(_02168_ ), .ZN(_02169_ ) );
MUX2_X1 _22851_ ( .A(_02145_ ), .B(_02169_ ), .S(_01504_ ), .Z(_02170_ ) );
MUX2_X1 _22852_ ( .A(_02134_ ), .B(_02170_ ), .S(_01214_ ), .Z(_02171_ ) );
MUX2_X1 _22853_ ( .A(_02118_ ), .B(_02171_ ), .S(_02023_ ), .Z(_02172_ ) );
MUX2_X1 _22854_ ( .A(_02117_ ), .B(_02172_ ), .S(_01180_ ), .Z(_02173_ ) );
MUX2_X1 _22855_ ( .A(_02102_ ), .B(_02173_ ), .S(_01176_ ), .Z(_02174_ ) );
AND2_X1 _22856_ ( .A1(_02174_ ), .A2(_01175_ ), .ZN(_02175_ ) );
NOR3_X1 _22857_ ( .A1(_02096_ ), .A2(_09046_ ), .A3(_09047_ ), .ZN(_02176_ ) );
OAI21_X1 _22858_ ( .A(_01171_ ), .B1(_02175_ ), .B2(_02176_ ), .ZN(_02177_ ) );
NAND2_X1 _22859_ ( .A1(\exu.addi._io_rd_T_4 [18] ), .A2(_01870_ ), .ZN(_02178_ ) );
AOI21_X1 _22860_ ( .A(_01718_ ), .B1(_02177_ ), .B2(_02178_ ), .ZN(_02179_ ) );
AND3_X1 _22861_ ( .A1(_01718_ ), .A2(_10844_ ), .A3(\exu.csrrs.io_csr_rdata [18] ), .ZN(_02180_ ) );
OR2_X1 _22862_ ( .A1(_02179_ ), .A2(_02180_ ), .ZN(\exu.io_out_bits_rd_wdata [18] ) );
AND3_X1 _22863_ ( .A1(_01730_ ), .A2(_01732_ ), .A3(_01561_ ), .ZN(_02181_ ) );
NAND3_X1 _22864_ ( .A1(_01900_ ), .A2(_01902_ ), .A3(_01892_ ), .ZN(_02182_ ) );
OAI211_X1 _22865_ ( .A(_01725_ ), .B(_02182_ ), .C1(_01729_ ), .C2(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02183_ ) );
AND3_X1 _22866_ ( .A1(_01726_ ), .A2(_01727_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02184_ ) );
AOI21_X1 _22867_ ( .A(_01320_ ), .B1(_01726_ ), .B2(_01727_ ), .ZN(_02185_ ) );
OAI21_X1 _22868_ ( .A(_01559_ ), .B1(_02184_ ), .B2(_02185_ ), .ZN(_02186_ ) );
AOI21_X1 _22869_ ( .A(_01561_ ), .B1(_02183_ ), .B2(_02186_ ), .ZN(_02187_ ) );
OR2_X1 _22870_ ( .A1(_02181_ ), .A2(_02187_ ), .ZN(_02188_ ) );
AND3_X1 _22871_ ( .A1(_01737_ ), .A2(_01740_ ), .A3(_01546_ ), .ZN(_02189_ ) );
AOI21_X1 _22872_ ( .A(_02189_ ), .B1(_01744_ ), .B2(_01562_ ), .ZN(_02190_ ) );
MUX2_X1 _22873_ ( .A(_02188_ ), .B(_02190_ ), .S(_01746_ ), .Z(_02191_ ) );
NAND2_X1 _22874_ ( .A1(_02191_ ), .A2(_01880_ ), .ZN(_02192_ ) );
NAND3_X1 _22875_ ( .A1(_02192_ ), .A2(_01914_ ), .A3(_01537_ ), .ZN(_02193_ ) );
NAND3_X1 _22876_ ( .A1(_01404_ ), .A2(_10699_ ), .A3(fanout_net_4 ), .ZN(_02194_ ) );
AND3_X1 _22877_ ( .A1(_02192_ ), .A2(_01445_ ), .A3(_01537_ ), .ZN(_02195_ ) );
OAI21_X1 _22878_ ( .A(_01581_ ), .B1(\exu.add.io_rs1_data [17] ), .B2(\exu._GEN_0 [17] ), .ZN(_02196_ ) );
OAI211_X1 _22879_ ( .A(_01771_ ), .B(_01782_ ), .C1(_01786_ ), .C2(_01587_ ), .ZN(_02197_ ) );
OAI211_X1 _22880_ ( .A(_01589_ ), .B(_01774_ ), .C1(_01777_ ), .C2(_01778_ ), .ZN(_02198_ ) );
NAND3_X1 _22881_ ( .A1(_02197_ ), .A2(_01790_ ), .A3(_02198_ ), .ZN(_02199_ ) );
NAND3_X1 _22882_ ( .A1(_01762_ ), .A2(_01770_ ), .A3(_01768_ ), .ZN(_02200_ ) );
OAI21_X1 _22883_ ( .A(_01781_ ), .B1(_02026_ ), .B2(_02027_ ), .ZN(_02201_ ) );
AND3_X1 _22884_ ( .A1(_01189_ ), .A2(_01192_ ), .A3(_01657_ ), .ZN(_02202_ ) );
AOI21_X1 _22885_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01758_ ), .B2(_01759_ ), .ZN(_02203_ ) );
OAI21_X1 _22886_ ( .A(_01763_ ), .B1(_02202_ ), .B2(_02203_ ), .ZN(_02204_ ) );
NAND3_X1 _22887_ ( .A1(_02201_ ), .A2(_02204_ ), .A3(_01589_ ), .ZN(_02205_ ) );
NAND3_X1 _22888_ ( .A1(_02200_ ), .A2(_01591_ ), .A3(_02205_ ), .ZN(_02206_ ) );
NAND2_X1 _22889_ ( .A1(_02199_ ), .A2(_02206_ ), .ZN(_02207_ ) );
AND3_X1 _22890_ ( .A1(_02207_ ), .A2(_01212_ ), .A3(_01594_ ), .ZN(_02208_ ) );
AOI211_X1 _22891_ ( .A(_08878_ ), .B(_01597_ ), .C1(_02062_ ), .C2(_08747_ ), .ZN(_02209_ ) );
OAI21_X1 _22892_ ( .A(_08746_ ), .B1(_08877_ ), .B2(\exu._GEN_0 [16] ), .ZN(_02210_ ) );
OAI21_X1 _22893_ ( .A(_02209_ ), .B1(_02062_ ), .B2(_02210_ ), .ZN(_02211_ ) );
AND4_X1 _22894_ ( .A1(\exu.addi.io_imm [17] ), .A2(_01601_ ), .A3(_01602_ ), .A4(_01604_ ), .ZN(_02212_ ) );
AOI21_X1 _22895_ ( .A(_02212_ ), .B1(_10072_ ), .B2(_01607_ ), .ZN(_02213_ ) );
OAI21_X1 _22896_ ( .A(_02211_ ), .B1(_02213_ ), .B2(\exu.io_in_bits_sub ), .ZN(_02214_ ) );
AOI21_X1 _22897_ ( .A(_02208_ ), .B1(_02214_ ), .B2(_01610_ ), .ZN(_02215_ ) );
OAI21_X1 _22898_ ( .A(_02196_ ), .B1(_02215_ ), .B2(\exu.io_in_bits_or ), .ZN(_02216_ ) );
AOI21_X1 _22899_ ( .A(_02195_ ), .B1(_02216_ ), .B2(_01614_ ), .ZN(_02217_ ) );
OAI21_X1 _22900_ ( .A(_02194_ ), .B1(_02217_ ), .B2(fanout_net_4 ), .ZN(_02218_ ) );
AOI221_X4 _22901_ ( .A(fanout_net_12 ), .B1(_08746_ ), .B2(_01493_ ), .C1(_02218_ ), .C2(_01618_ ), .ZN(_02219_ ) );
NOR3_X1 _22902_ ( .A1(_01231_ ), .A2(_01241_ ), .A3(_01254_ ), .ZN(_02220_ ) );
NAND3_X1 _22903_ ( .A1(_02220_ ), .A2(_01654_ ), .A3(_01686_ ), .ZN(_02221_ ) );
NAND2_X1 _22904_ ( .A1(_01802_ ), .A2(_01325_ ), .ZN(_02222_ ) );
NAND3_X1 _22905_ ( .A1(_01816_ ), .A2(_01817_ ), .A3(_01279_ ), .ZN(_02223_ ) );
NAND2_X1 _22906_ ( .A1(_02222_ ), .A2(_02223_ ), .ZN(_02224_ ) );
AOI21_X1 _22907_ ( .A(_01306_ ), .B1(_01813_ ), .B2(_01814_ ), .ZN(_02225_ ) );
AOI21_X1 _22908_ ( .A(_01325_ ), .B1(_01809_ ), .B2(_01810_ ), .ZN(_02226_ ) );
NOR2_X1 _22909_ ( .A1(_02225_ ), .A2(_02226_ ), .ZN(_02227_ ) );
MUX2_X1 _22910_ ( .A(_02224_ ), .B(_02227_ ), .S(_01686_ ), .Z(_02228_ ) );
OAI21_X1 _22911_ ( .A(_02221_ ), .B1(_02228_ ), .B2(_01654_ ), .ZN(_02229_ ) );
NAND2_X1 _22912_ ( .A1(_02229_ ), .A2(_01689_ ), .ZN(_02230_ ) );
AOI211_X1 _22913_ ( .A(_01574_ ), .B(_02219_ ), .C1(fanout_net_12 ), .C2(_02230_ ), .ZN(_02231_ ) );
AND3_X1 _22914_ ( .A1(_02077_ ), .A2(_08747_ ), .A3(_02078_ ), .ZN(_02232_ ) );
NOR3_X1 _22915_ ( .A1(_02232_ ), .A2(_02079_ ), .A3(_01694_ ), .ZN(_02233_ ) );
OAI21_X1 _22916_ ( .A(_01571_ ), .B1(_02231_ ), .B2(_02233_ ), .ZN(_02234_ ) );
OR2_X1 _22917_ ( .A1(_10066_ ), .A2(_01823_ ), .ZN(_02235_ ) );
AOI21_X1 _22918_ ( .A(\exu.io_in_bits_jalr ), .B1(_02234_ ), .B2(_02235_ ), .ZN(_02236_ ) );
NOR2_X1 _22919_ ( .A1(_10066_ ), .A2(_01855_ ), .ZN(_02237_ ) );
OAI21_X1 _22920_ ( .A(_01570_ ), .B1(_02236_ ), .B2(_02237_ ), .ZN(_02238_ ) );
NAND2_X1 _22921_ ( .A1(_02229_ ), .A2(_01702_ ), .ZN(_02239_ ) );
NAND3_X1 _22922_ ( .A1(_02238_ ), .A2(_01507_ ), .A3(_02239_ ), .ZN(_02240_ ) );
AOI211_X1 _22923_ ( .A(_01795_ ), .B(_01797_ ), .C1(_02199_ ), .C2(_02206_ ), .ZN(_02241_ ) );
OAI211_X1 _22924_ ( .A(_02240_ ), .B(_01510_ ), .C1(_01705_ ), .C2(_02241_ ), .ZN(_02242_ ) );
AOI21_X1 _22925_ ( .A(\exu.io_in_bits_srai ), .B1(_09131_ ), .B2(_01186_ ), .ZN(_02243_ ) );
AOI221_X4 _22926_ ( .A(fanout_net_5 ), .B1(\exu.io_in_bits_srai ), .B2(_02193_ ), .C1(_02242_ ), .C2(_02243_ ), .ZN(_02244_ ) );
AND3_X1 _22927_ ( .A1(_09127_ ), .A2(_10843_ ), .A3(fanout_net_5 ), .ZN(_02245_ ) );
OAI21_X1 _22928_ ( .A(_01175_ ), .B1(_02244_ ), .B2(_02245_ ), .ZN(_02246_ ) );
NAND2_X1 _22929_ ( .A1(_09129_ ), .A2(_01519_ ), .ZN(_02247_ ) );
AOI21_X1 _22930_ ( .A(_01173_ ), .B1(_02246_ ), .B2(_02247_ ), .ZN(_02248_ ) );
INV_X1 _22931_ ( .A(_01523_ ), .ZN(_02249_ ) );
NOR2_X1 _22932_ ( .A1(_10093_ ), .A2(_02249_ ), .ZN(_02250_ ) );
OAI21_X1 _22933_ ( .A(_01108_ ), .B1(_02248_ ), .B2(_02250_ ), .ZN(_02251_ ) );
INV_X1 _22934_ ( .A(_02251_ ), .ZN(_02252_ ) );
AND3_X1 _22935_ ( .A1(_01718_ ), .A2(_01873_ ), .A3(\exu.csrrs.io_csr_rdata [17] ), .ZN(_02253_ ) );
NOR2_X1 _22936_ ( .A1(_02252_ ), .A2(_02253_ ), .ZN(_02254_ ) );
INV_X1 _22937_ ( .A(_02254_ ), .ZN(\exu.io_out_bits_rd_wdata [17] ) );
NAND3_X1 _22938_ ( .A1(_01886_ ), .A2(_01893_ ), .A3(_01562_ ), .ZN(_02255_ ) );
OAI21_X1 _22939_ ( .A(_01899_ ), .B1(_02106_ ), .B2(_02107_ ), .ZN(_02256_ ) );
BUF_X2 _22940_ ( .A(_01900_ ), .Z(_02257_ ) );
BUF_X2 _22941_ ( .A(_01902_ ), .Z(_02258_ ) );
AND3_X1 _22942_ ( .A1(_02257_ ), .A2(_02258_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02259_ ) );
AOI21_X1 _22943_ ( .A(_01661_ ), .B1(_02257_ ), .B2(_02258_ ), .ZN(_02260_ ) );
OAI21_X1 _22944_ ( .A(_01887_ ), .B1(_02259_ ), .B2(_02260_ ), .ZN(_02261_ ) );
NAND2_X1 _22945_ ( .A1(_02256_ ), .A2(_02261_ ), .ZN(_02262_ ) );
NAND2_X1 _22946_ ( .A1(_02262_ ), .A2(_01547_ ), .ZN(_02263_ ) );
AOI21_X1 _22947_ ( .A(_01747_ ), .B1(_02255_ ), .B2(_02263_ ), .ZN(_02264_ ) );
NAND2_X1 _22948_ ( .A1(_01898_ ), .A2(_01905_ ), .ZN(_02265_ ) );
MUX2_X1 _22949_ ( .A(_02265_ ), .B(_01911_ ), .S(_01562_ ), .Z(_02266_ ) );
AOI21_X1 _22950_ ( .A(_02264_ ), .B1(_02266_ ), .B2(_01747_ ), .ZN(_02267_ ) );
OAI21_X1 _22951_ ( .A(_01536_ ), .B1(_02267_ ), .B2(_01568_ ), .ZN(_02268_ ) );
NOR2_X1 _22952_ ( .A1(_02268_ ), .A2(_01752_ ), .ZN(_02269_ ) );
OAI21_X1 _22953_ ( .A(_01878_ ), .B1(_02269_ ), .B2(_01512_ ), .ZN(_02270_ ) );
OAI21_X1 _22954_ ( .A(_01755_ ), .B1(\exu.add.io_rs1_data [16] ), .B2(\exu.addi.io_imm [16] ), .ZN(_02271_ ) );
AND3_X1 _22955_ ( .A1(_01920_ ), .A2(_01200_ ), .A3(_01925_ ), .ZN(_02272_ ) );
AOI21_X1 _22956_ ( .A(_02272_ ), .B1(_01940_ ), .B2(_01771_ ), .ZN(_02273_ ) );
NOR2_X1 _22957_ ( .A1(_02273_ ), .A2(_01591_ ), .ZN(_02274_ ) );
AND3_X1 _22958_ ( .A1(_01930_ ), .A2(_01770_ ), .A3(_01932_ ), .ZN(_02275_ ) );
OAI21_X1 _22959_ ( .A(_01587_ ), .B1(_02119_ ), .B2(_02120_ ), .ZN(_02276_ ) );
AND3_X1 _22960_ ( .A1(_01922_ ), .A2(_01923_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02277_ ) );
AOI21_X1 _22961_ ( .A(_01661_ ), .B1(_01922_ ), .B2(_01923_ ), .ZN(_02278_ ) );
OAI21_X1 _22962_ ( .A(_01763_ ), .B1(_02277_ ), .B2(_02278_ ), .ZN(_02279_ ) );
AOI21_X1 _22963_ ( .A(_01771_ ), .B1(_02276_ ), .B2(_02279_ ), .ZN(_02280_ ) );
OR2_X1 _22964_ ( .A1(_02275_ ), .A2(_02280_ ), .ZN(_02281_ ) );
AOI21_X1 _22965_ ( .A(_02274_ ), .B1(_01205_ ), .B2(_02281_ ), .ZN(_02282_ ) );
BUF_X2 _22966_ ( .A(_01217_ ), .Z(_02283_ ) );
NAND3_X1 _22967_ ( .A1(_02282_ ), .A2(_01213_ ), .A3(_02283_ ), .ZN(_02284_ ) );
NAND4_X1 _22968_ ( .A1(_01944_ ), .A2(_01804_ ), .A3(_01686_ ), .A4(_01306_ ), .ZN(_02285_ ) );
NAND2_X1 _22969_ ( .A1(_01948_ ), .A2(_01241_ ), .ZN(_02286_ ) );
OR3_X1 _22970_ ( .A1(_01624_ ), .A2(_01291_ ), .A3(_01625_ ), .ZN(_02287_ ) );
OAI211_X1 _22971_ ( .A(_02287_ ), .B(_01279_ ), .C1(_01254_ ), .C2(_01650_ ), .ZN(_02288_ ) );
NAND2_X1 _22972_ ( .A1(_02286_ ), .A2(_02288_ ), .ZN(_02289_ ) );
AND3_X1 _22973_ ( .A1(_01958_ ), .A2(_01279_ ), .A3(_01959_ ), .ZN(_02290_ ) );
AND3_X1 _22974_ ( .A1(_01954_ ), .A2(_01955_ ), .A3(_01241_ ), .ZN(_02291_ ) );
OR2_X1 _22975_ ( .A1(_02290_ ), .A2(_02291_ ), .ZN(_02292_ ) );
MUX2_X1 _22976_ ( .A(_02289_ ), .B(_02292_ ), .S(_01271_ ), .Z(_02293_ ) );
OAI21_X1 _22977_ ( .A(_02285_ ), .B1(_02293_ ), .B2(_01804_ ), .ZN(_02294_ ) );
NAND2_X1 _22978_ ( .A1(_02294_ ), .A2(_01702_ ), .ZN(_02295_ ) );
NAND3_X1 _22979_ ( .A1(_01405_ ), .A2(_01575_ ), .A3(fanout_net_4 ), .ZN(_02296_ ) );
NOR2_X1 _22980_ ( .A1(_02268_ ), .A2(_01579_ ), .ZN(_02297_ ) );
OAI21_X1 _22981_ ( .A(_01581_ ), .B1(\exu.add.io_rs1_data [16] ), .B2(\exu._GEN_0 [16] ), .ZN(_02298_ ) );
AND3_X1 _22982_ ( .A1(_02282_ ), .A2(_01212_ ), .A3(_01594_ ), .ZN(_02299_ ) );
NOR3_X1 _22983_ ( .A1(_08840_ ), .A2(_08749_ ), .A3(_08865_ ), .ZN(_02300_ ) );
OR3_X1 _22984_ ( .A1(_02062_ ), .A2(_01597_ ), .A3(_02300_ ), .ZN(_02301_ ) );
AND4_X1 _22985_ ( .A1(\exu.addi.io_imm [16] ), .A2(_01600_ ), .A3(_01463_ ), .A4(_01603_ ), .ZN(_02302_ ) );
AOI21_X1 _22986_ ( .A(_02302_ ), .B1(_09876_ ), .B2(_01607_ ), .ZN(_02303_ ) );
OAI21_X1 _22987_ ( .A(_02301_ ), .B1(_02303_ ), .B2(\exu.io_in_bits_sub ), .ZN(_02304_ ) );
AOI21_X1 _22988_ ( .A(_02299_ ), .B1(_02304_ ), .B2(_01610_ ), .ZN(_02305_ ) );
OAI21_X1 _22989_ ( .A(_02298_ ), .B1(_02305_ ), .B2(\exu.io_in_bits_or ), .ZN(_02306_ ) );
AOI21_X1 _22990_ ( .A(_02297_ ), .B1(_02306_ ), .B2(_01613_ ), .ZN(_02307_ ) );
OAI21_X1 _22991_ ( .A(_02296_ ), .B1(_02307_ ), .B2(fanout_net_4 ), .ZN(_02308_ ) );
AOI221_X4 _22992_ ( .A(fanout_net_12 ), .B1(_08748_ ), .B2(_01968_ ), .C1(_02308_ ), .C2(_01618_ ), .ZN(_02309_ ) );
NAND2_X1 _22993_ ( .A1(_02294_ ), .A2(_01689_ ), .ZN(_02310_ ) );
AOI211_X1 _22994_ ( .A(_01574_ ), .B(_02309_ ), .C1(fanout_net_12 ), .C2(_02310_ ), .ZN(_02311_ ) );
XNOR2_X1 _22995_ ( .A(_01391_ ), .B(_08748_ ), .ZN(_02312_ ) );
AOI21_X1 _22996_ ( .A(_02311_ ), .B1(_01828_ ), .B2(_02312_ ), .ZN(_02313_ ) );
OAI221_X1 _22997_ ( .A(_01341_ ), .B1(_01823_ ), .B2(_09881_ ), .C1(_02313_ ), .C2(\exu.io_in_bits_jal ), .ZN(_02314_ ) );
AND2_X1 _22998_ ( .A1(_09880_ ), .A2(_01699_ ), .ZN(_02315_ ) );
OAI211_X1 _22999_ ( .A(_02314_ ), .B(_01989_ ), .C1(_01854_ ), .C2(_02315_ ), .ZN(_02316_ ) );
MUX2_X1 _23000_ ( .A(_02295_ ), .B(_02316_ ), .S(_01992_ ), .Z(_02317_ ) );
MUX2_X1 _23001_ ( .A(_02284_ ), .B(_02317_ ), .S(_01994_ ), .Z(_02318_ ) );
MUX2_X1 _23002_ ( .A(_02271_ ), .B(_02318_ ), .S(_01860_ ), .Z(_02319_ ) );
AOI21_X1 _23003_ ( .A(_02270_ ), .B1(_02319_ ), .B2(_01862_ ), .ZN(_02320_ ) );
AND3_X1 _23004_ ( .A1(_09124_ ), .A2(_10844_ ), .A3(fanout_net_5 ), .ZN(_02321_ ) );
OAI21_X1 _23005_ ( .A(_01877_ ), .B1(_02320_ ), .B2(_02321_ ), .ZN(_02322_ ) );
NAND2_X1 _23006_ ( .A1(_09126_ ), .A2(_02000_ ), .ZN(_02323_ ) );
AOI21_X1 _23007_ ( .A(_01876_ ), .B1(_02322_ ), .B2(_02323_ ), .ZN(_02324_ ) );
AND2_X1 _23008_ ( .A1(\exu.addi._io_rd_T_4 [16] ), .A2(_02003_ ), .ZN(_02325_ ) );
OAI21_X1 _23009_ ( .A(_01875_ ), .B1(_02324_ ), .B2(_02325_ ), .ZN(_02326_ ) );
OAI211_X1 _23010_ ( .A(_01058_ ), .B(\exu.csrrs.io_csr_rdata [16] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_02327_ ) );
NAND2_X1 _23011_ ( .A1(_02326_ ), .A2(_02327_ ), .ZN(\exu.io_out_bits_rd_wdata [16] ) );
AND3_X1 _23012_ ( .A1(_09103_ ), .A2(_10843_ ), .A3(fanout_net_5 ), .ZN(_02328_ ) );
OR3_X1 _23013_ ( .A1(_02184_ ), .A2(_02185_ ), .A3(_01559_ ), .ZN(_02329_ ) );
NAND3_X1 _23014_ ( .A1(_02257_ ), .A2(_02258_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02330_ ) );
OAI211_X1 _23015_ ( .A(_01887_ ), .B(_02330_ ), .C1(_01890_ ), .C2(_01277_ ), .ZN(_02331_ ) );
NAND3_X1 _23016_ ( .A1(_02329_ ), .A2(_01546_ ), .A3(_02331_ ), .ZN(_02332_ ) );
NAND3_X1 _23017_ ( .A1(_02012_ ), .A2(_02014_ ), .A3(_01562_ ), .ZN(_02333_ ) );
NAND2_X1 _23018_ ( .A1(_02332_ ), .A2(_02333_ ), .ZN(_02334_ ) );
AND2_X1 _23019_ ( .A1(_02009_ ), .A2(_02010_ ), .ZN(_02335_ ) );
MUX2_X1 _23020_ ( .A(_02335_ ), .B(_02018_ ), .S(_01561_ ), .Z(_02336_ ) );
MUX2_X1 _23021_ ( .A(_02334_ ), .B(_02336_ ), .S(_01747_ ), .Z(_02337_ ) );
AOI211_X1 _23022_ ( .A(_01751_ ), .B(_01534_ ), .C1(_02337_ ), .C2(_02021_ ), .ZN(_02338_ ) );
NOR3_X1 _23023_ ( .A1(_09104_ ), .A2(fanout_net_27 ), .A3(_02023_ ), .ZN(_02339_ ) );
OR3_X1 _23024_ ( .A1(_02202_ ), .A2(_02203_ ), .A3(_01197_ ), .ZN(_02340_ ) );
AND3_X1 _23025_ ( .A1(_01758_ ), .A2(_01759_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02341_ ) );
AOI21_X1 _23026_ ( .A(_01277_ ), .B1(_01190_ ), .B2(_01193_ ), .ZN(_02342_ ) );
OAI21_X1 _23027_ ( .A(_01197_ ), .B1(_02341_ ), .B2(_02342_ ), .ZN(_02343_ ) );
AND3_X1 _23028_ ( .A1(_02340_ ), .A2(_01200_ ), .A3(_02343_ ), .ZN(_02344_ ) );
AOI21_X1 _23029_ ( .A(_01200_ ), .B1(_02025_ ), .B2(_02028_ ), .ZN(_02345_ ) );
OAI21_X1 _23030_ ( .A(_01205_ ), .B1(_02344_ ), .B2(_02345_ ), .ZN(_02346_ ) );
AOI21_X1 _23031_ ( .A(_01200_ ), .B1(_02037_ ), .B2(_02038_ ), .ZN(_02347_ ) );
AOI21_X1 _23032_ ( .A(_01770_ ), .B1(_02032_ ), .B2(_02033_ ), .ZN(_02348_ ) );
OR2_X1 _23033_ ( .A1(_02347_ ), .A2(_02348_ ), .ZN(_02349_ ) );
OAI211_X1 _23034_ ( .A(_01211_ ), .B(_02346_ ), .C1(_02349_ ), .C2(_01205_ ), .ZN(_02350_ ) );
INV_X1 _23035_ ( .A(_01201_ ), .ZN(_02351_ ) );
OAI21_X1 _23036_ ( .A(_01793_ ), .B1(_02351_ ), .B2(_01790_ ), .ZN(_02352_ ) );
AND3_X1 _23037_ ( .A1(_02350_ ), .A2(_01217_ ), .A3(_02352_ ), .ZN(_02353_ ) );
BUF_X2 _23038_ ( .A(_01332_ ), .Z(_02354_ ) );
CLKBUF_X2 _23039_ ( .A(_02354_ ), .Z(_02355_ ) );
AND3_X1 _23040_ ( .A1(_01282_ ), .A2(_02355_ ), .A3(_01337_ ), .ZN(_02356_ ) );
NAND3_X1 _23041_ ( .A1(_01384_ ), .A2(_09463_ ), .A3(fanout_net_4 ), .ZN(_02357_ ) );
NAND2_X1 _23042_ ( .A1(_02337_ ), .A2(_01879_ ), .ZN(_02358_ ) );
AND3_X1 _23043_ ( .A1(_02358_ ), .A2(_01444_ ), .A3(_01536_ ), .ZN(_02359_ ) );
OAI21_X1 _23044_ ( .A(_01447_ ), .B1(\exu.add.io_rs1_data [15] ), .B2(\exu._GEN_0 [15] ), .ZN(_02360_ ) );
AND3_X1 _23045_ ( .A1(_02350_ ), .A2(_01593_ ), .A3(_02352_ ), .ZN(_02361_ ) );
AND4_X1 _23046_ ( .A1(\exu.addi.io_imm [15] ), .A2(_01464_ ), .A3(_01458_ ), .A4(_01466_ ), .ZN(_02362_ ) );
AOI21_X1 _23047_ ( .A(_02362_ ), .B1(_09837_ ), .B2(_01459_ ), .ZN(_02363_ ) );
OR2_X1 _23048_ ( .A1(_02363_ ), .A2(\exu.io_in_bits_sub ), .ZN(_02364_ ) );
AND2_X1 _23049_ ( .A1(_08830_ ), .A2(_08839_ ), .ZN(_02365_ ) );
NOR2_X1 _23050_ ( .A1(_02365_ ), .A2(_08714_ ), .ZN(_02366_ ) );
AND2_X1 _23051_ ( .A1(_02366_ ), .A2(_08713_ ), .ZN(_02367_ ) );
INV_X1 _23052_ ( .A(_02367_ ), .ZN(_02368_ ) );
OAI21_X1 _23053_ ( .A(_08852_ ), .B1(_02368_ ), .B2(_08847_ ), .ZN(_02369_ ) );
NAND2_X1 _23054_ ( .A1(_02369_ ), .A2(_08724_ ), .ZN(_02370_ ) );
AOI21_X1 _23055_ ( .A(_08718_ ), .B1(_02370_ ), .B2(_08858_ ), .ZN(_02371_ ) );
INV_X1 _23056_ ( .A(_02371_ ), .ZN(_02372_ ) );
OAI21_X1 _23057_ ( .A(_02372_ ), .B1(_08860_ ), .B2(\exu._GEN_0 [14] ), .ZN(_02373_ ) );
XOR2_X1 _23058_ ( .A(_02373_ ), .B(_08717_ ), .Z(_02374_ ) );
OAI21_X1 _23059_ ( .A(_02364_ ), .B1(_01596_ ), .B2(_02374_ ), .ZN(_02375_ ) );
AOI21_X1 _23060_ ( .A(_02361_ ), .B1(_02375_ ), .B2(_01481_ ), .ZN(_02376_ ) );
OAI21_X1 _23061_ ( .A(_02360_ ), .B1(_02376_ ), .B2(\exu.io_in_bits_or ), .ZN(_02377_ ) );
AOI21_X1 _23062_ ( .A(_02359_ ), .B1(_02377_ ), .B2(_01443_ ), .ZN(_02378_ ) );
OAI21_X1 _23063_ ( .A(_02357_ ), .B1(_02378_ ), .B2(fanout_net_4 ), .ZN(_02379_ ) );
AOI221_X4 _23064_ ( .A(fanout_net_12 ), .B1(_08717_ ), .B2(_01492_ ), .C1(_02379_ ), .C2(_01617_ ), .ZN(_02380_ ) );
NAND3_X1 _23065_ ( .A1(_01282_ ), .A2(_01333_ ), .A3(_01440_ ), .ZN(_02381_ ) );
AOI211_X1 _23066_ ( .A(_01573_ ), .B(_02380_ ), .C1(fanout_net_12 ), .C2(_02381_ ), .ZN(_02382_ ) );
INV_X1 _23067_ ( .A(_08718_ ), .ZN(_02383_ ) );
NOR2_X1 _23068_ ( .A1(_01373_ ), .A2(_08728_ ), .ZN(_02384_ ) );
NOR4_X1 _23069_ ( .A1(_02384_ ), .A2(_08713_ ), .A3(_08715_ ), .A4(_01378_ ), .ZN(_02385_ ) );
OAI211_X1 _23070_ ( .A(_08723_ ), .B(_08720_ ), .C1(_02385_ ), .C2(_01382_ ), .ZN(_02386_ ) );
AOI21_X1 _23071_ ( .A(_02383_ ), .B1(_02386_ ), .B2(_01386_ ), .ZN(_02387_ ) );
OR3_X1 _23072_ ( .A1(_02387_ ), .A2(_08717_ ), .A3(_01388_ ), .ZN(_02388_ ) );
OAI21_X1 _23073_ ( .A(_08717_ ), .B1(_02387_ ), .B2(_01388_ ), .ZN(_02389_ ) );
AND3_X1 _23074_ ( .A1(_02388_ ), .A2(_01436_ ), .A3(_02389_ ), .ZN(_02390_ ) );
OAI21_X1 _23075_ ( .A(_09410_ ), .B1(_02382_ ), .B2(_02390_ ), .ZN(_02391_ ) );
OAI21_X1 _23076_ ( .A(_02391_ ), .B1(_01342_ ), .B2(_09835_ ), .ZN(_02392_ ) );
NAND2_X1 _23077_ ( .A1(_02392_ ), .A2(_01340_ ), .ZN(_02393_ ) );
OR2_X1 _23078_ ( .A1(_09835_ ), .A2(_01855_ ), .ZN(_02394_ ) );
AOI21_X1 _23079_ ( .A(\exu.io_out_bits_ren ), .B1(_02393_ ), .B2(_02394_ ), .ZN(_02395_ ) );
MUX2_X1 _23080_ ( .A(_02356_ ), .B(_02395_ ), .S(_01504_ ), .Z(_02396_ ) );
MUX2_X1 _23081_ ( .A(_02353_ ), .B(_02396_ ), .S(_01507_ ), .Z(_02397_ ) );
MUX2_X1 _23082_ ( .A(_02339_ ), .B(_02397_ ), .S(_01509_ ), .Z(_02398_ ) );
MUX2_X1 _23083_ ( .A(_02338_ ), .B(_02398_ ), .S(_01182_ ), .Z(_02399_ ) );
MUX2_X1 _23084_ ( .A(_02328_ ), .B(_02399_ ), .S(_01878_ ), .Z(_02400_ ) );
NAND2_X1 _23085_ ( .A1(_02400_ ), .A2(_01877_ ), .ZN(_02401_ ) );
NAND2_X1 _23086_ ( .A1(_09105_ ), .A2(_02000_ ), .ZN(_02402_ ) );
AOI21_X1 _23087_ ( .A(_01876_ ), .B1(_02401_ ), .B2(_02402_ ), .ZN(_02403_ ) );
AND2_X1 _23088_ ( .A1(\exu.addi._io_rd_T_4 [15] ), .A2(_01870_ ), .ZN(_02404_ ) );
OAI21_X1 _23089_ ( .A(_01721_ ), .B1(_02403_ ), .B2(_02404_ ), .ZN(_02405_ ) );
OAI211_X1 _23090_ ( .A(_10845_ ), .B(\exu.csrrs.io_csr_rdata [15] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_02406_ ) );
NAND2_X1 _23091_ ( .A1(_02405_ ), .A2(_02406_ ), .ZN(\exu.io_out_bits_rd_wdata [15] ) );
AND3_X1 _23092_ ( .A1(_09106_ ), .A2(_10843_ ), .A3(fanout_net_5 ), .ZN(_02407_ ) );
OAI21_X1 _23093_ ( .A(_01899_ ), .B1(_01895_ ), .B2(_01896_ ), .ZN(_02408_ ) );
AND3_X1 _23094_ ( .A1(_02103_ ), .A2(_01546_ ), .A3(_02408_ ), .ZN(_02409_ ) );
AND3_X1 _23095_ ( .A1(_02111_ ), .A2(_02113_ ), .A3(_01561_ ), .ZN(_02410_ ) );
OR3_X1 _23096_ ( .A1(_02409_ ), .A2(_01541_ ), .A3(_02410_ ), .ZN(_02411_ ) );
OAI21_X1 _23097_ ( .A(_01899_ ), .B1(_02259_ ), .B2(_02260_ ), .ZN(_02412_ ) );
AND3_X1 _23098_ ( .A1(_01900_ ), .A2(_01902_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02413_ ) );
AOI21_X1 _23099_ ( .A(_01638_ ), .B1(_01900_ ), .B2(_01902_ ), .ZN(_02414_ ) );
OAI21_X1 _23100_ ( .A(_01887_ ), .B1(_02413_ ), .B2(_02414_ ), .ZN(_02415_ ) );
NAND2_X1 _23101_ ( .A1(_02412_ ), .A2(_02415_ ), .ZN(_02416_ ) );
NAND2_X1 _23102_ ( .A1(_02416_ ), .A2(_01734_ ), .ZN(_02417_ ) );
OAI211_X1 _23103_ ( .A(_01562_ ), .B(_02105_ ), .C1(_02108_ ), .C2(_01884_ ), .ZN(_02418_ ) );
NAND2_X1 _23104_ ( .A1(_02417_ ), .A2(_02418_ ), .ZN(_02419_ ) );
OAI211_X1 _23105_ ( .A(_02411_ ), .B(_01879_ ), .C1(_01748_ ), .C2(_02419_ ), .ZN(_02420_ ) );
OAI21_X1 _23106_ ( .A(_02420_ ), .B1(_01879_ ), .B2(_01565_ ), .ZN(_02421_ ) );
NOR2_X1 _23107_ ( .A1(_02421_ ), .A2(_01752_ ), .ZN(_02422_ ) );
NOR3_X1 _23108_ ( .A1(_09107_ ), .A2(fanout_net_27 ), .A3(_01509_ ), .ZN(_02423_ ) );
OR2_X1 _23109_ ( .A1(_01592_ ), .A2(_01211_ ), .ZN(_02424_ ) );
AND3_X1 _23110_ ( .A1(_01764_ ), .A2(_01765_ ), .A3(_01277_ ), .ZN(_02425_ ) );
AOI21_X1 _23111_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B1(_01764_ ), .B2(_01765_ ), .ZN(_02426_ ) );
OR3_X1 _23112_ ( .A1(_02425_ ), .A2(_01586_ ), .A3(_02426_ ), .ZN(_02427_ ) );
OAI21_X1 _23113_ ( .A(_01781_ ), .B1(_02277_ ), .B2(_02278_ ), .ZN(_02428_ ) );
NAND2_X1 _23114_ ( .A1(_02427_ ), .A2(_02428_ ), .ZN(_02429_ ) );
NAND2_X1 _23115_ ( .A1(_02429_ ), .A2(_01590_ ), .ZN(_02430_ ) );
NAND3_X1 _23116_ ( .A1(_02121_ ), .A2(_01771_ ), .A3(_02122_ ), .ZN(_02431_ ) );
NAND3_X1 _23117_ ( .A1(_02430_ ), .A2(_01205_ ), .A3(_02431_ ), .ZN(_02432_ ) );
NAND3_X1 _23118_ ( .A1(_02124_ ), .A2(_01590_ ), .A3(_02125_ ), .ZN(_02433_ ) );
NAND3_X1 _23119_ ( .A1(_02129_ ), .A2(_02130_ ), .A3(_01771_ ), .ZN(_02434_ ) );
AND2_X1 _23120_ ( .A1(_02433_ ), .A2(_02434_ ), .ZN(_02435_ ) );
OAI211_X1 _23121_ ( .A(_02432_ ), .B(_01211_ ), .C1(_01205_ ), .C2(_02435_ ), .ZN(_02436_ ) );
AND3_X1 _23122_ ( .A1(_02424_ ), .A2(_01217_ ), .A3(_02436_ ), .ZN(_02437_ ) );
AND3_X1 _23123_ ( .A1(_01653_ ), .A2(_02355_ ), .A3(_01337_ ), .ZN(_02438_ ) );
NAND3_X1 _23124_ ( .A1(_01388_ ), .A2(_09463_ ), .A3(fanout_net_4 ), .ZN(_02439_ ) );
NOR2_X1 _23125_ ( .A1(_02421_ ), .A2(_01578_ ), .ZN(_02440_ ) );
OAI21_X1 _23126_ ( .A(_01448_ ), .B1(\exu.add.io_rs1_data [14] ), .B2(\exu._GEN_0 [14] ), .ZN(_02441_ ) );
AND3_X1 _23127_ ( .A1(_02424_ ), .A2(_01593_ ), .A3(_02436_ ), .ZN(_02442_ ) );
NAND3_X1 _23128_ ( .A1(_02370_ ), .A2(_08718_ ), .A3(_08858_ ), .ZN(_02443_ ) );
NAND3_X1 _23129_ ( .A1(_02372_ ), .A2(_01477_ ), .A3(_02443_ ), .ZN(_02444_ ) );
AND4_X1 _23130_ ( .A1(\exu.addi.io_imm [14] ), .A2(_01465_ ), .A3(_01462_ ), .A4(_01467_ ), .ZN(_02445_ ) );
AOI21_X1 _23131_ ( .A(_02445_ ), .B1(_10115_ ), .B2(_01606_ ), .ZN(_02446_ ) );
OAI21_X1 _23132_ ( .A(_02444_ ), .B1(_02446_ ), .B2(\exu.io_in_bits_sub ), .ZN(_02447_ ) );
AOI21_X1 _23133_ ( .A(_02442_ ), .B1(_02447_ ), .B2(_01481_ ), .ZN(_02448_ ) );
OAI21_X1 _23134_ ( .A(_02441_ ), .B1(_02448_ ), .B2(\exu.io_in_bits_or ), .ZN(_02449_ ) );
AOI21_X1 _23135_ ( .A(_02440_ ), .B1(_02449_ ), .B2(_01443_ ), .ZN(_02450_ ) );
OAI21_X1 _23136_ ( .A(_02439_ ), .B1(_02450_ ), .B2(fanout_net_4 ), .ZN(_02451_ ) );
AOI221_X4 _23137_ ( .A(fanout_net_12 ), .B1(_08718_ ), .B2(_01492_ ), .C1(_02451_ ), .C2(_01617_ ), .ZN(_02452_ ) );
NAND3_X1 _23138_ ( .A1(_01653_ ), .A2(_01333_ ), .A3(_01441_ ), .ZN(_02453_ ) );
AOI211_X1 _23139_ ( .A(_01573_ ), .B(_02452_ ), .C1(fanout_net_12 ), .C2(_02453_ ), .ZN(_02454_ ) );
AND3_X1 _23140_ ( .A1(_02386_ ), .A2(_02383_ ), .A3(_01386_ ), .ZN(_02455_ ) );
NOR3_X1 _23141_ ( .A1(_02455_ ), .A2(_02387_ ), .A3(_01694_ ), .ZN(_02456_ ) );
OAI21_X1 _23142_ ( .A(_09410_ ), .B1(_02454_ ), .B2(_02456_ ), .ZN(_02457_ ) );
OAI21_X1 _23143_ ( .A(_02457_ ), .B1(_01342_ ), .B2(_10131_ ), .ZN(_02458_ ) );
NAND2_X1 _23144_ ( .A1(_02458_ ), .A2(_01340_ ), .ZN(_02459_ ) );
NAND2_X1 _23145_ ( .A1(_10121_ ), .A2(_09460_ ), .ZN(_02460_ ) );
AOI21_X1 _23146_ ( .A(\exu.io_out_bits_ren ), .B1(_02459_ ), .B2(_02460_ ), .ZN(_02461_ ) );
MUX2_X1 _23147_ ( .A(_02438_ ), .B(_02461_ ), .S(_01505_ ), .Z(_02462_ ) );
MUX2_X1 _23148_ ( .A(_02437_ ), .B(_02462_ ), .S(_01507_ ), .Z(_02463_ ) );
MUX2_X1 _23149_ ( .A(_02423_ ), .B(_02463_ ), .S(_01509_ ), .Z(_02464_ ) );
MUX2_X1 _23150_ ( .A(_02422_ ), .B(_02464_ ), .S(_01182_ ), .Z(_02465_ ) );
MUX2_X1 _23151_ ( .A(_02407_ ), .B(_02465_ ), .S(_01878_ ), .Z(_02466_ ) );
NAND2_X1 _23152_ ( .A1(_02466_ ), .A2(_01877_ ), .ZN(_02467_ ) );
NAND2_X1 _23153_ ( .A1(_09108_ ), .A2(_02000_ ), .ZN(_02468_ ) );
AOI21_X1 _23154_ ( .A(_01876_ ), .B1(_02467_ ), .B2(_02468_ ), .ZN(_02469_ ) );
NOR3_X1 _23155_ ( .A1(_10144_ ), .A2(_09859_ ), .A3(_02249_ ), .ZN(_02470_ ) );
OAI21_X1 _23156_ ( .A(_01875_ ), .B1(_02469_ ), .B2(_02470_ ), .ZN(_02471_ ) );
OAI211_X1 _23157_ ( .A(_01058_ ), .B(\exu.csrrs.io_csr_rdata [14] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_02472_ ) );
NAND2_X1 _23158_ ( .A1(_02471_ ), .A2(_02472_ ), .ZN(\exu.io_out_bits_rd_wdata [14] ) );
AND3_X1 _23159_ ( .A1(_09109_ ), .A2(_10842_ ), .A3(fanout_net_5 ), .ZN(_02473_ ) );
OAI211_X1 _23160_ ( .A(_01899_ ), .B(_02330_ ), .C1(_01890_ ), .C2(_01277_ ), .ZN(_02474_ ) );
NAND3_X1 _23161_ ( .A1(_02257_ ), .A2(_02258_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02475_ ) );
OAI211_X1 _23162_ ( .A(_01887_ ), .B(_02475_ ), .C1(_01890_ ), .C2(_01274_ ), .ZN(_02476_ ) );
AND2_X1 _23163_ ( .A1(_02474_ ), .A2(_02476_ ), .ZN(_02477_ ) );
OR2_X1 _23164_ ( .A1(_02477_ ), .A2(_01882_ ), .ZN(_02478_ ) );
NAND3_X1 _23165_ ( .A1(_02183_ ), .A2(_02186_ ), .A3(_01882_ ), .ZN(_02479_ ) );
AOI21_X1 _23166_ ( .A(_01747_ ), .B1(_02478_ ), .B2(_02479_ ), .ZN(_02480_ ) );
NOR3_X1 _23167_ ( .A1(_01733_ ), .A2(_01741_ ), .A3(_01564_ ), .ZN(_02481_ ) );
OR3_X1 _23168_ ( .A1(_02480_ ), .A2(_01567_ ), .A3(_02481_ ), .ZN(_02482_ ) );
MUX2_X1 _23169_ ( .A(_01177_ ), .B(_01745_ ), .S(_01540_ ), .Z(_02483_ ) );
OAI21_X1 _23170_ ( .A(_02482_ ), .B1(_02483_ ), .B2(_01880_ ), .ZN(_02484_ ) );
NOR2_X1 _23171_ ( .A1(_02484_ ), .A2(_01751_ ), .ZN(_02485_ ) );
NOR3_X1 _23172_ ( .A1(_09110_ ), .A2(fanout_net_27 ), .A3(_02023_ ), .ZN(_02486_ ) );
OR3_X1 _23173_ ( .A1(_02341_ ), .A2(_02342_ ), .A3(_01761_ ), .ZN(_02487_ ) );
AND3_X1 _23174_ ( .A1(_01190_ ), .A2(_01193_ ), .A3(_01638_ ), .ZN(_02488_ ) );
AOI21_X1 _23175_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01764_ ), .B2(_01765_ ), .ZN(_02489_ ) );
OAI21_X1 _23176_ ( .A(_01763_ ), .B1(_02488_ ), .B2(_02489_ ), .ZN(_02490_ ) );
AOI21_X1 _23177_ ( .A(_01771_ ), .B1(_02487_ ), .B2(_02490_ ), .ZN(_02491_ ) );
AOI21_X1 _23178_ ( .A(_01590_ ), .B1(_02201_ ), .B2(_02204_ ), .ZN(_02492_ ) );
NOR3_X1 _23179_ ( .A1(_02491_ ), .A2(_01790_ ), .A3(_02492_ ), .ZN(_02493_ ) );
AOI21_X1 _23180_ ( .A(_01205_ ), .B1(_01769_ ), .B2(_01779_ ), .ZN(_02494_ ) );
NOR3_X1 _23181_ ( .A1(_02493_ ), .A2(_02494_ ), .A3(_01793_ ), .ZN(_02495_ ) );
AND3_X1 _23182_ ( .A1(_01787_ ), .A2(_01589_ ), .A3(_01204_ ), .ZN(_02496_ ) );
AOI21_X1 _23183_ ( .A(_02495_ ), .B1(_01794_ ), .B2(_02496_ ), .ZN(_02497_ ) );
NOR2_X1 _23184_ ( .A1(_02497_ ), .A2(_01797_ ), .ZN(_02498_ ) );
NAND2_X1 _23185_ ( .A1(_01803_ ), .A2(_01245_ ), .ZN(_02499_ ) );
OAI21_X1 _23186_ ( .A(_02499_ ), .B1(_01246_ ), .B2(_01819_ ), .ZN(_02500_ ) );
AND3_X1 _23187_ ( .A1(_02500_ ), .A2(_02355_ ), .A3(_01337_ ), .ZN(_02501_ ) );
OR2_X1 _23188_ ( .A1(_02497_ ), .A2(_01455_ ), .ZN(_02502_ ) );
AND2_X1 _23189_ ( .A1(_02369_ ), .A2(_01348_ ), .ZN(_02503_ ) );
INV_X1 _23190_ ( .A(_02503_ ), .ZN(_02504_ ) );
OAI21_X1 _23191_ ( .A(_02504_ ), .B1(_08855_ ), .B2(\exu._GEN_0 [12] ), .ZN(_02505_ ) );
OAI21_X1 _23192_ ( .A(_01477_ ), .B1(_02505_ ), .B2(_01349_ ), .ZN(_02506_ ) );
AOI21_X1 _23193_ ( .A(_02506_ ), .B1(_01349_ ), .B2(_02505_ ), .ZN(_02507_ ) );
NAND4_X1 _23194_ ( .A1(_01600_ ), .A2(\exu.addi.io_imm [13] ), .A3(_01463_ ), .A4(_01603_ ), .ZN(_02508_ ) );
OAI21_X1 _23195_ ( .A(_02508_ ), .B1(_10178_ ), .B2(_01460_ ), .ZN(_02509_ ) );
AOI21_X1 _23196_ ( .A(_02507_ ), .B1(_02509_ ), .B2(_01457_ ), .ZN(_02510_ ) );
OAI21_X1 _23197_ ( .A(_02502_ ), .B1(_02510_ ), .B2(\exu.io_in_bits_srl ), .ZN(_02511_ ) );
BUF_X2 _23198_ ( .A(_01446_ ), .Z(_02512_ ) );
AND2_X1 _23199_ ( .A1(_02511_ ), .A2(_02512_ ), .ZN(_02513_ ) );
NOR3_X1 _23200_ ( .A1(_08722_ ), .A2(fanout_net_27 ), .A3(_02512_ ), .ZN(_02514_ ) );
OAI21_X1 _23201_ ( .A(_01613_ ), .B1(_02513_ ), .B2(_02514_ ), .ZN(_02515_ ) );
OR2_X1 _23202_ ( .A1(_02484_ ), .A2(_01578_ ), .ZN(_02516_ ) );
AOI21_X1 _23203_ ( .A(fanout_net_4 ), .B1(_02515_ ), .B2(_02516_ ), .ZN(_02517_ ) );
AND3_X1 _23204_ ( .A1(_08721_ ), .A2(_10698_ ), .A3(fanout_net_4 ), .ZN(_02518_ ) );
OAI21_X1 _23205_ ( .A(_01617_ ), .B1(_02517_ ), .B2(_02518_ ), .ZN(_02519_ ) );
NAND2_X1 _23206_ ( .A1(_08723_ ), .A2(_01968_ ), .ZN(_02520_ ) );
AOI21_X1 _23207_ ( .A(fanout_net_12 ), .B1(_02519_ ), .B2(_02520_ ), .ZN(_02521_ ) );
AND3_X1 _23208_ ( .A1(_02500_ ), .A2(_01333_ ), .A3(_01440_ ), .ZN(_02522_ ) );
OAI21_X1 _23209_ ( .A(_01498_ ), .B1(_02521_ ), .B2(_02522_ ), .ZN(_02523_ ) );
OAI21_X1 _23210_ ( .A(_01352_ ), .B1(_01373_ ), .B2(_08728_ ), .ZN(_02524_ ) );
INV_X1 _23211_ ( .A(_01382_ ), .ZN(_02525_ ) );
AOI21_X1 _23212_ ( .A(_01348_ ), .B1(_02524_ ), .B2(_02525_ ), .ZN(_02526_ ) );
OR3_X1 _23213_ ( .A1(_02526_ ), .A2(_08723_ ), .A3(_01385_ ), .ZN(_02527_ ) );
OAI21_X1 _23214_ ( .A(_08723_ ), .B1(_02526_ ), .B2(_01385_ ), .ZN(_02528_ ) );
NAND3_X1 _23215_ ( .A1(_02527_ ), .A2(_01436_ ), .A3(_02528_ ), .ZN(_02529_ ) );
AOI21_X1 _23216_ ( .A(\exu.io_in_bits_jal ), .B1(_02523_ ), .B2(_02529_ ), .ZN(_02530_ ) );
NOR2_X1 _23217_ ( .A1(_10165_ ), .A2(_09999_ ), .ZN(_02531_ ) );
OAI21_X1 _23218_ ( .A(_01340_ ), .B1(_02530_ ), .B2(_02531_ ), .ZN(_02532_ ) );
OR2_X1 _23219_ ( .A1(_10165_ ), .A2(_01855_ ), .ZN(_02533_ ) );
AOI21_X1 _23220_ ( .A(\exu.io_out_bits_ren ), .B1(_02532_ ), .B2(_02533_ ), .ZN(_02534_ ) );
MUX2_X1 _23221_ ( .A(_02501_ ), .B(_02534_ ), .S(_01504_ ), .Z(_02535_ ) );
MUX2_X1 _23222_ ( .A(_02498_ ), .B(_02535_ ), .S(_01214_ ), .Z(_02536_ ) );
MUX2_X1 _23223_ ( .A(_02486_ ), .B(_02536_ ), .S(_01509_ ), .Z(_02537_ ) );
MUX2_X1 _23224_ ( .A(_02485_ ), .B(_02537_ ), .S(_01181_ ), .Z(_02538_ ) );
MUX2_X1 _23225_ ( .A(_02473_ ), .B(_02538_ ), .S(_01515_ ), .Z(_02539_ ) );
NAND2_X1 _23226_ ( .A1(_02539_ ), .A2(_01723_ ), .ZN(_02540_ ) );
NAND2_X1 _23227_ ( .A1(_09111_ ), .A2(_01867_ ), .ZN(_02541_ ) );
AOI21_X1 _23228_ ( .A(_01722_ ), .B1(_02540_ ), .B2(_02541_ ), .ZN(_02542_ ) );
AND2_X1 _23229_ ( .A1(\exu.addi._io_rd_T_4 [13] ), .A2(_01870_ ), .ZN(_02543_ ) );
OAI21_X1 _23230_ ( .A(_01721_ ), .B1(_02542_ ), .B2(_02543_ ), .ZN(_02544_ ) );
OAI211_X1 _23231_ ( .A(_01873_ ), .B(\exu.csrrs.io_csr_rdata [13] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_02545_ ) );
NAND2_X1 _23232_ ( .A1(_02544_ ), .A2(_02545_ ), .ZN(\exu.io_out_bits_rd_wdata [13] ) );
OAI21_X1 _23233_ ( .A(_01748_ ), .B1(_01894_ ), .B2(_01906_ ), .ZN(_02546_ ) );
NAND2_X1 _23234_ ( .A1(_02262_ ), .A2(_01882_ ), .ZN(_02547_ ) );
OR3_X1 _23235_ ( .A1(_02413_ ), .A2(_02414_ ), .A3(_01887_ ), .ZN(_02548_ ) );
NAND3_X1 _23236_ ( .A1(_01901_ ), .A2(_01903_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02549_ ) );
OAI211_X1 _23237_ ( .A(_01888_ ), .B(_02549_ ), .C1(_01891_ ), .C2(_01642_ ), .ZN(_02550_ ) );
NAND3_X1 _23238_ ( .A1(_02548_ ), .A2(_01734_ ), .A3(_02550_ ), .ZN(_02551_ ) );
NAND2_X1 _23239_ ( .A1(_02547_ ), .A2(_02551_ ), .ZN(_02552_ ) );
OAI211_X1 _23240_ ( .A(_02546_ ), .B(_01879_ ), .C1(_01748_ ), .C2(_02552_ ), .ZN(_02553_ ) );
AOI21_X1 _23241_ ( .A(_01542_ ), .B1(_01912_ ), .B2(_01881_ ), .ZN(_02554_ ) );
OAI21_X1 _23242_ ( .A(_02553_ ), .B1(_02554_ ), .B2(_01880_ ), .ZN(_02555_ ) );
NOR2_X1 _23243_ ( .A1(_02555_ ), .A2(_01752_ ), .ZN(_02556_ ) );
OAI21_X1 _23244_ ( .A(_01515_ ), .B1(_02556_ ), .B2(_01512_ ), .ZN(_02557_ ) );
OAI21_X1 _23245_ ( .A(_01755_ ), .B1(\exu.add.io_rs1_data [12] ), .B2(\exu.addi.io_imm [12] ), .ZN(_02558_ ) );
AND3_X1 _23246_ ( .A1(_02276_ ), .A2(_02279_ ), .A3(_01927_ ), .ZN(_02559_ ) );
OAI21_X1 _23247_ ( .A(_01587_ ), .B1(_02425_ ), .B2(_02426_ ), .ZN(_02560_ ) );
AND3_X1 _23248_ ( .A1(_01922_ ), .A2(_01923_ ), .A3(_01274_ ), .ZN(_02561_ ) );
BUF_X2 _23249_ ( .A(_01764_ ), .Z(_02562_ ) );
BUF_X2 _23250_ ( .A(_01765_ ), .Z(_02563_ ) );
AOI21_X1 _23251_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B1(_02562_ ), .B2(_02563_ ), .ZN(_02564_ ) );
OAI21_X1 _23252_ ( .A(_01778_ ), .B1(_02561_ ), .B2(_02564_ ), .ZN(_02565_ ) );
AOI21_X1 _23253_ ( .A(_01927_ ), .B1(_02560_ ), .B2(_02565_ ), .ZN(_02566_ ) );
OAI21_X1 _23254_ ( .A(_01206_ ), .B1(_02559_ ), .B2(_02566_ ), .ZN(_02567_ ) );
OAI211_X1 _23255_ ( .A(_01211_ ), .B(_02567_ ), .C1(_01934_ ), .C2(_01206_ ), .ZN(_02568_ ) );
NOR3_X1 _23256_ ( .A1(_01940_ ), .A2(_01927_ ), .A3(_01935_ ), .ZN(_02569_ ) );
OAI211_X1 _23257_ ( .A(_02283_ ), .B(_02568_ ), .C1(_02569_ ), .C2(_01213_ ), .ZN(_02570_ ) );
MUX2_X1 _23258_ ( .A(_01957_ ), .B(_01949_ ), .S(_01308_ ), .Z(_02571_ ) );
INV_X1 _23259_ ( .A(_01338_ ), .ZN(_02572_ ) );
OR3_X1 _23260_ ( .A1(_02571_ ), .A2(_01654_ ), .A3(_02572_ ), .ZN(_02573_ ) );
NAND3_X1 _23261_ ( .A1(_01385_ ), .A2(_10698_ ), .A3(fanout_net_4 ), .ZN(_02574_ ) );
NOR2_X1 _23262_ ( .A1(_02555_ ), .A2(_01579_ ), .ZN(_02575_ ) );
OAI21_X1 _23263_ ( .A(_01448_ ), .B1(\exu.add.io_rs1_data [12] ), .B2(\exu._GEN_0 [12] ), .ZN(_02576_ ) );
OAI21_X1 _23264_ ( .A(_02568_ ), .B1(_02569_ ), .B2(_01450_ ), .ZN(_02577_ ) );
NOR2_X1 _23265_ ( .A1(_02577_ ), .A2(_01455_ ), .ZN(_02578_ ) );
AOI21_X1 _23266_ ( .A(_01597_ ), .B1(_02369_ ), .B2(_01348_ ), .ZN(_02579_ ) );
OAI21_X1 _23267_ ( .A(_02579_ ), .B1(_01348_ ), .B2(_02369_ ), .ZN(_02580_ ) );
AND4_X1 _23268_ ( .A1(\exu.addi.io_imm [12] ), .A2(_01600_ ), .A3(_01463_ ), .A4(_01603_ ), .ZN(_02581_ ) );
AOI21_X1 _23269_ ( .A(_02581_ ), .B1(_10354_ ), .B2(_01606_ ), .ZN(_02582_ ) );
OAI21_X1 _23270_ ( .A(_02580_ ), .B1(_02582_ ), .B2(\exu.io_in_bits_sub ), .ZN(_02583_ ) );
AOI21_X1 _23271_ ( .A(_02578_ ), .B1(_02583_ ), .B2(_01481_ ), .ZN(_02584_ ) );
OAI21_X1 _23272_ ( .A(_02576_ ), .B1(_02584_ ), .B2(\exu.io_in_bits_or ), .ZN(_02585_ ) );
AOI21_X1 _23273_ ( .A(_02575_ ), .B1(_02585_ ), .B2(_01613_ ), .ZN(_02586_ ) );
OAI21_X1 _23274_ ( .A(_02574_ ), .B1(_02586_ ), .B2(fanout_net_4 ), .ZN(_02587_ ) );
AOI221_X4 _23275_ ( .A(fanout_net_12 ), .B1(_08720_ ), .B2(_01968_ ), .C1(_02587_ ), .C2(_01618_ ), .ZN(_02588_ ) );
INV_X1 _23276_ ( .A(_01440_ ), .ZN(_02589_ ) );
OR3_X1 _23277_ ( .A1(_02571_ ), .A2(_01804_ ), .A3(_02589_ ), .ZN(_02590_ ) );
AOI211_X1 _23278_ ( .A(_01574_ ), .B(_02588_ ), .C1(fanout_net_12 ), .C2(_02590_ ), .ZN(_02591_ ) );
AND3_X1 _23279_ ( .A1(_02524_ ), .A2(_01348_ ), .A3(_02525_ ), .ZN(_02592_ ) );
NOR3_X1 _23280_ ( .A1(_02592_ ), .A2(_02526_ ), .A3(_01694_ ), .ZN(_02593_ ) );
OAI21_X1 _23281_ ( .A(_01571_ ), .B1(_02591_ ), .B2(_02593_ ), .ZN(_02594_ ) );
NAND2_X1 _23282_ ( .A1(_10356_ ), .A2(_09452_ ), .ZN(_02595_ ) );
AOI21_X1 _23283_ ( .A(\exu.io_in_bits_jalr ), .B1(_02594_ ), .B2(_02595_ ), .ZN(_02596_ ) );
AND2_X1 _23284_ ( .A1(_10356_ ), .A2(_01699_ ), .ZN(_02597_ ) );
OAI21_X1 _23285_ ( .A(_01989_ ), .B1(_02596_ ), .B2(_02597_ ), .ZN(_02598_ ) );
MUX2_X1 _23286_ ( .A(_02573_ ), .B(_02598_ ), .S(_01505_ ), .Z(_02599_ ) );
MUX2_X1 _23287_ ( .A(_02570_ ), .B(_02599_ ), .S(_01705_ ), .Z(_02600_ ) );
MUX2_X1 _23288_ ( .A(_02558_ ), .B(_02600_ ), .S(_01860_ ), .Z(_02601_ ) );
AOI21_X1 _23289_ ( .A(_02557_ ), .B1(_02601_ ), .B2(_01862_ ), .ZN(_02602_ ) );
AND3_X1 _23290_ ( .A1(_09112_ ), .A2(_01864_ ), .A3(fanout_net_5 ), .ZN(_02603_ ) );
OAI21_X1 _23291_ ( .A(_01723_ ), .B1(_02602_ ), .B2(_02603_ ), .ZN(_02604_ ) );
NAND2_X1 _23292_ ( .A1(_09114_ ), .A2(_01867_ ), .ZN(_02605_ ) );
AOI21_X1 _23293_ ( .A(_01722_ ), .B1(_02604_ ), .B2(_02605_ ), .ZN(_02606_ ) );
AND2_X1 _23294_ ( .A1(\exu.addi._io_rd_T_4 [12] ), .A2(_01870_ ), .ZN(_02607_ ) );
OAI21_X1 _23295_ ( .A(_01721_ ), .B1(_02606_ ), .B2(_02607_ ), .ZN(_02608_ ) );
OAI211_X1 _23296_ ( .A(_01873_ ), .B(\exu.csrrs.io_csr_rdata [12] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_02609_ ) );
NAND2_X1 _23297_ ( .A1(_02608_ ), .A2(_02609_ ), .ZN(\exu.io_out_bits_rd_wdata [12] ) );
NAND3_X1 _23298_ ( .A1(_09699_ ), .A2(_10842_ ), .A3(fanout_net_5 ), .ZN(_02610_ ) );
OAI211_X1 _23299_ ( .A(_01530_ ), .B(_01537_ ), .C1(_02483_ ), .C2(_01568_ ), .ZN(_02611_ ) );
OAI21_X1 _23300_ ( .A(_01185_ ), .B1(\exu.add.io_rs1_data [29] ), .B2(\exu.addi.io_imm [29] ), .ZN(_02612_ ) );
NAND3_X1 _23301_ ( .A1(_02496_ ), .A2(_01212_ ), .A3(_01216_ ), .ZN(_02613_ ) );
NAND2_X1 _23302_ ( .A1(_02500_ ), .A2(_01331_ ), .ZN(_02614_ ) );
NAND2_X1 _23303_ ( .A1(_01288_ ), .A2(_01290_ ), .ZN(_02615_ ) );
OAI21_X1 _23304_ ( .A(_01235_ ), .B1(_01314_ ), .B2(_01316_ ), .ZN(_02616_ ) );
NAND2_X1 _23305_ ( .A1(_02615_ ), .A2(_02616_ ), .ZN(_02617_ ) );
OR2_X1 _23306_ ( .A1(_01292_ ), .A2(_01294_ ), .ZN(_02618_ ) );
MUX2_X1 _23307_ ( .A(_01304_ ), .B(_02618_ ), .S(_01235_ ), .Z(_02619_ ) );
MUX2_X1 _23308_ ( .A(_02617_ ), .B(_02619_ ), .S(_01252_ ), .Z(_02620_ ) );
MUX2_X1 _23309_ ( .A(_01812_ ), .B(_02620_ ), .S(_01270_ ), .Z(_02621_ ) );
OAI21_X1 _23310_ ( .A(_02614_ ), .B1(_01331_ ), .B2(_02621_ ), .ZN(_02622_ ) );
NAND2_X1 _23311_ ( .A1(_02622_ ), .A2(_01336_ ), .ZN(_02623_ ) );
OR3_X1 _23312_ ( .A1(_01426_ ), .A2(_08764_ ), .A3(_01427_ ), .ZN(_02624_ ) );
AND3_X1 _23313_ ( .A1(_02624_ ), .A2(_01428_ ), .A3(_01435_ ), .ZN(_02625_ ) );
NAND2_X1 _23314_ ( .A1(_02622_ ), .A2(_01440_ ), .ZN(_02626_ ) );
MUX2_X1 _23315_ ( .A(_01177_ ), .B(_02483_ ), .S(_01533_ ), .Z(_02627_ ) );
OAI21_X1 _23316_ ( .A(_01447_ ), .B1(\exu.add.io_rs1_data [29] ), .B2(\exu._GEN_0 [29] ), .ZN(_02628_ ) );
AND3_X1 _23317_ ( .A1(_02496_ ), .A2(_01211_ ), .A3(_01593_ ), .ZN(_02629_ ) );
AND4_X1 _23318_ ( .A1(\exu.addi.io_imm [29] ), .A2(_01464_ ), .A3(_01458_ ), .A4(_01466_ ), .ZN(_02630_ ) );
AOI21_X1 _23319_ ( .A(_02630_ ), .B1(_09782_ ), .B2(_01459_ ), .ZN(_02631_ ) );
OR2_X1 _23320_ ( .A1(_02631_ ), .A2(\exu.io_in_bits_sub ), .ZN(_02632_ ) );
NOR2_X1 _23321_ ( .A1(_01472_ ), .A2(_08765_ ), .ZN(_02633_ ) );
INV_X1 _23322_ ( .A(_02633_ ), .ZN(_02634_ ) );
OAI21_X1 _23323_ ( .A(_02634_ ), .B1(_08867_ ), .B2(\exu._GEN_0 [28] ), .ZN(_02635_ ) );
XOR2_X1 _23324_ ( .A(_02635_ ), .B(_08764_ ), .Z(_02636_ ) );
OAI21_X1 _23325_ ( .A(_02632_ ), .B1(_01596_ ), .B2(_02636_ ), .ZN(_02637_ ) );
AOI21_X1 _23326_ ( .A(_02629_ ), .B1(_02637_ ), .B2(_01452_ ), .ZN(_02638_ ) );
OAI21_X1 _23327_ ( .A(_02628_ ), .B1(_02638_ ), .B2(\exu.io_in_bits_or ), .ZN(_02639_ ) );
AOI221_X4 _23328_ ( .A(fanout_net_4 ), .B1(_01444_ ), .B2(_02627_ ), .C1(_02639_ ), .C2(_01443_ ), .ZN(_02640_ ) );
NAND3_X1 _23329_ ( .A1(_01429_ ), .A2(_09463_ ), .A3(fanout_net_4 ), .ZN(_02641_ ) );
AOI211_X1 _23330_ ( .A(\exu.io_in_bits_xor ), .B(_02640_ ), .C1(fanout_net_4 ), .C2(_02641_ ), .ZN(_02642_ ) );
AOI21_X1 _23331_ ( .A(_02642_ ), .B1(_08764_ ), .B2(_01492_ ), .ZN(_02643_ ) );
OAI21_X1 _23332_ ( .A(_02626_ ), .B1(_02643_ ), .B2(fanout_net_12 ), .ZN(_02644_ ) );
AOI21_X1 _23333_ ( .A(_02625_ ), .B1(_02644_ ), .B2(_01498_ ), .ZN(_02645_ ) );
OAI221_X1 _23334_ ( .A(_09657_ ), .B1(_09999_ ), .B2(_09788_ ), .C1(_02645_ ), .C2(\exu.io_in_bits_jal ), .ZN(_02646_ ) );
AND3_X1 _23335_ ( .A1(_09785_ ), .A2(_09460_ ), .A3(_09787_ ), .ZN(_02647_ ) );
OAI211_X1 _23336_ ( .A(_02646_ ), .B(_01501_ ), .C1(_09657_ ), .C2(_02647_ ), .ZN(_02648_ ) );
MUX2_X1 _23337_ ( .A(_02623_ ), .B(_02648_ ), .S(_01219_ ), .Z(_02649_ ) );
MUX2_X1 _23338_ ( .A(_02613_ ), .B(_02649_ ), .S(_01214_ ), .Z(_02650_ ) );
MUX2_X1 _23339_ ( .A(_02612_ ), .B(_02650_ ), .S(_01184_ ), .Z(_02651_ ) );
MUX2_X1 _23340_ ( .A(_02611_ ), .B(_02651_ ), .S(_01180_ ), .Z(_02652_ ) );
MUX2_X1 _23341_ ( .A(_02610_ ), .B(_02652_ ), .S(_01176_ ), .Z(_02653_ ) );
OR2_X1 _23342_ ( .A1(_02653_ ), .A2(\exu.io_in_bits_xori ), .ZN(_02654_ ) );
NAND2_X1 _23343_ ( .A1(_09701_ ), .A2(_01519_ ), .ZN(_02655_ ) );
AOI21_X1 _23344_ ( .A(_01173_ ), .B1(_02654_ ), .B2(_02655_ ), .ZN(_02656_ ) );
AOI21_X1 _23345_ ( .A(_02656_ ), .B1(\exu.addi._io_rd_T_4 [29] ), .B2(_01870_ ), .ZN(_02657_ ) );
NOR2_X1 _23346_ ( .A1(_02657_ ), .A2(_01718_ ), .ZN(_02658_ ) );
NOR3_X1 _23347_ ( .A1(_01109_ ), .A2(fanout_net_27 ), .A3(_09683_ ), .ZN(_02659_ ) );
NOR2_X1 _23348_ ( .A1(_02658_ ), .A2(_02659_ ), .ZN(_02660_ ) );
INV_X1 _23349_ ( .A(_02660_ ), .ZN(\exu.io_out_bits_rd_wdata [29] ) );
NAND3_X1 _23350_ ( .A1(_02329_ ), .A2(_01882_ ), .A3(_02331_ ), .ZN(_02661_ ) );
OAI211_X1 _23351_ ( .A(_01899_ ), .B(_02475_ ), .C1(_01890_ ), .C2(_01274_ ), .ZN(_02662_ ) );
NAND3_X1 _23352_ ( .A1(_01901_ ), .A2(_01903_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02663_ ) );
OAI211_X1 _23353_ ( .A(_01887_ ), .B(_02663_ ), .C1(_01890_ ), .C2(_01261_ ), .ZN(_02664_ ) );
NAND3_X1 _23354_ ( .A1(_02662_ ), .A2(_02664_ ), .A3(_01734_ ), .ZN(_02665_ ) );
NAND3_X1 _23355_ ( .A1(_02661_ ), .A2(_01564_ ), .A3(_02665_ ), .ZN(_02666_ ) );
OAI211_X1 _23356_ ( .A(_02666_ ), .B(_01879_ ), .C1(_02016_ ), .C2(_01564_ ), .ZN(_02667_ ) );
AOI21_X1 _23357_ ( .A(_01542_ ), .B1(_02019_ ), .B2(_01564_ ), .ZN(_02668_ ) );
OAI211_X1 _23358_ ( .A(_01530_ ), .B(_02667_ ), .C1(_02668_ ), .C2(_02021_ ), .ZN(_02669_ ) );
AND3_X1 _23359_ ( .A1(_02040_ ), .A2(_01205_ ), .A3(_01793_ ), .ZN(_02670_ ) );
NAND2_X1 _23360_ ( .A1(_02340_ ), .A2(_02343_ ), .ZN(_02671_ ) );
NAND2_X1 _23361_ ( .A1(_02671_ ), .A2(_01927_ ), .ZN(_02672_ ) );
AND3_X1 _23362_ ( .A1(_01758_ ), .A2(_01759_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02673_ ) );
AOI21_X1 _23363_ ( .A(_01261_ ), .B1(_01758_ ), .B2(_01759_ ), .ZN(_02674_ ) );
OR3_X1 _23364_ ( .A1(_02673_ ), .A2(_01586_ ), .A3(_02674_ ), .ZN(_02675_ ) );
OAI21_X1 _23365_ ( .A(_01586_ ), .B1(_02488_ ), .B2(_02489_ ), .ZN(_02676_ ) );
NAND3_X1 _23366_ ( .A1(_02675_ ), .A2(_01788_ ), .A3(_02676_ ), .ZN(_02677_ ) );
AOI21_X1 _23367_ ( .A(_01790_ ), .B1(_02672_ ), .B2(_02677_ ), .ZN(_02678_ ) );
AND3_X1 _23368_ ( .A1(_02030_ ), .A2(_02034_ ), .A3(_01790_ ), .ZN(_02679_ ) );
NOR3_X1 _23369_ ( .A1(_02678_ ), .A2(_02679_ ), .A3(_01794_ ), .ZN(_02680_ ) );
OAI21_X1 _23370_ ( .A(_01217_ ), .B1(_02670_ ), .B2(_02680_ ), .ZN(_02681_ ) );
AOI21_X1 _23371_ ( .A(\exu.io_in_bits_ori ), .B1(_02681_ ), .B2(\exu.io_in_bits_srli ), .ZN(_02682_ ) );
NOR2_X1 _23372_ ( .A1(_01236_ ), .A2(_01241_ ), .ZN(_02683_ ) );
MUX2_X1 _23373_ ( .A(_02050_ ), .B(_02683_ ), .S(_01246_ ), .Z(_02684_ ) );
AND3_X1 _23374_ ( .A1(_02684_ ), .A2(_02355_ ), .A3(_01338_ ), .ZN(_02685_ ) );
AOI21_X1 _23375_ ( .A(_08705_ ), .B1(_02368_ ), .B2(_08846_ ), .ZN(_02686_ ) );
AOI21_X1 _23376_ ( .A(_02686_ ), .B1(\exu.add.io_rs1_data [10] ), .B2(_01084_ ), .ZN(_02687_ ) );
OAI21_X1 _23377_ ( .A(_01477_ ), .B1(_02687_ ), .B2(_08708_ ), .ZN(_02688_ ) );
AOI21_X1 _23378_ ( .A(_02688_ ), .B1(_08708_ ), .B2(_02687_ ), .ZN(_02689_ ) );
NAND2_X1 _23379_ ( .A1(_10314_ ), .A2(_01606_ ), .ZN(_02690_ ) );
NAND4_X1 _23380_ ( .A1(_01465_ ), .A2(\exu.addi.io_imm [11] ), .A3(_01462_ ), .A4(_01467_ ), .ZN(_02691_ ) );
AOI21_X1 _23381_ ( .A(\exu.io_in_bits_sub ), .B1(_02690_ ), .B2(_02691_ ), .ZN(_02692_ ) );
OAI21_X1 _23382_ ( .A(_01481_ ), .B1(_02689_ ), .B2(_02692_ ), .ZN(_02693_ ) );
OAI21_X1 _23383_ ( .A(_01593_ ), .B1(_02670_ ), .B2(_02680_ ), .ZN(_02694_ ) );
AOI21_X1 _23384_ ( .A(\exu.io_in_bits_or ), .B1(_02693_ ), .B2(_02694_ ), .ZN(_02695_ ) );
AOI21_X1 _23385_ ( .A(_02695_ ), .B1(_01375_ ), .B2(_01448_ ), .ZN(_02696_ ) );
NOR2_X1 _23386_ ( .A1(_02696_ ), .A2(\exu.io_in_bits_sra ), .ZN(_02697_ ) );
OAI21_X1 _23387_ ( .A(_02667_ ), .B1(_02668_ ), .B2(_01880_ ), .ZN(_02698_ ) );
NOR2_X1 _23388_ ( .A1(_02698_ ), .A2(_01578_ ), .ZN(_02699_ ) );
OAI21_X1 _23389_ ( .A(_01486_ ), .B1(_02697_ ), .B2(_02699_ ), .ZN(_02700_ ) );
NAND3_X1 _23390_ ( .A1(_08706_ ), .A2(_10698_ ), .A3(fanout_net_4 ), .ZN(_02701_ ) );
AOI21_X1 _23391_ ( .A(\exu.io_in_bits_xor ), .B1(_02700_ ), .B2(_02701_ ), .ZN(_02702_ ) );
AOI211_X1 _23392_ ( .A(fanout_net_12 ), .B(_02702_ ), .C1(_08708_ ), .C2(_01968_ ), .ZN(_02703_ ) );
NAND3_X1 _23393_ ( .A1(_02684_ ), .A2(_01333_ ), .A3(_01441_ ), .ZN(_02704_ ) );
AOI211_X1 _23394_ ( .A(_01573_ ), .B(_02703_ ), .C1(fanout_net_12 ), .C2(_02704_ ), .ZN(_02705_ ) );
INV_X1 _23395_ ( .A(_01376_ ), .ZN(_02706_ ) );
OAI211_X1 _23396_ ( .A(_08712_ ), .B(_08714_ ), .C1(_01373_ ), .C2(_08728_ ), .ZN(_02707_ ) );
AND2_X1 _23397_ ( .A1(_02707_ ), .A2(_01381_ ), .ZN(_02708_ ) );
NOR2_X1 _23398_ ( .A1(\exu.add.io_rs1_data [10] ), .A2(\exu._GEN_0 [10] ), .ZN(_02709_ ) );
OAI21_X1 _23399_ ( .A(_02706_ ), .B1(_02708_ ), .B2(_02709_ ), .ZN(_02710_ ) );
XOR2_X1 _23400_ ( .A(_02710_ ), .B(_08708_ ), .Z(_02711_ ) );
AOI21_X1 _23401_ ( .A(_02705_ ), .B1(_01828_ ), .B2(_02711_ ), .ZN(_02712_ ) );
OR2_X1 _23402_ ( .A1(_02712_ ), .A2(\exu.io_in_bits_jal ), .ZN(_02713_ ) );
NAND3_X1 _23403_ ( .A1(_10308_ ), .A2(_09452_ ), .A3(_10310_ ), .ZN(_02714_ ) );
AOI21_X1 _23404_ ( .A(\exu.io_in_bits_jalr ), .B1(_02713_ ), .B2(_02714_ ), .ZN(_02715_ ) );
AOI21_X1 _23405_ ( .A(_02715_ ), .B1(_01699_ ), .B2(_10312_ ), .ZN(_02716_ ) );
NOR2_X1 _23406_ ( .A1(_02716_ ), .A2(\exu.io_out_bits_ren ), .ZN(_02717_ ) );
MUX2_X1 _23407_ ( .A(_02685_ ), .B(_02717_ ), .S(_01992_ ), .Z(_02718_ ) );
OAI21_X1 _23408_ ( .A(_02682_ ), .B1(_02718_ ), .B2(\exu.io_in_bits_srli ), .ZN(_02719_ ) );
AOI21_X1 _23409_ ( .A(\exu.io_in_bits_srai ), .B1(_09099_ ), .B2(_01186_ ), .ZN(_02720_ ) );
AOI221_X4 _23410_ ( .A(fanout_net_5 ), .B1(\exu.io_in_bits_srai ), .B2(_02669_ ), .C1(_02719_ ), .C2(_02720_ ), .ZN(_02721_ ) );
AND3_X1 _23411_ ( .A1(_09090_ ), .A2(_10843_ ), .A3(fanout_net_5 ), .ZN(_02722_ ) );
OAI21_X1 _23412_ ( .A(_01175_ ), .B1(_02721_ ), .B2(_02722_ ), .ZN(_02723_ ) );
NAND3_X1 _23413_ ( .A1(_09098_ ), .A2(_09099_ ), .A3(_01519_ ), .ZN(_02724_ ) );
AOI21_X1 _23414_ ( .A(_01173_ ), .B1(_02723_ ), .B2(_02724_ ), .ZN(_02725_ ) );
NOR2_X1 _23415_ ( .A1(_10343_ ), .A2(_02249_ ), .ZN(_02726_ ) );
OAI21_X1 _23416_ ( .A(_01108_ ), .B1(_02725_ ), .B2(_02726_ ), .ZN(_02727_ ) );
INV_X1 _23417_ ( .A(_02727_ ), .ZN(_02728_ ) );
NOR3_X1 _23418_ ( .A1(_01108_ ), .A2(fanout_net_27 ), .A3(_08960_ ), .ZN(_02729_ ) );
NOR2_X1 _23419_ ( .A1(_02728_ ), .A2(_02729_ ), .ZN(_02730_ ) );
INV_X1 _23420_ ( .A(_02730_ ), .ZN(\exu.io_out_bits_rd_wdata [11] ) );
AND3_X1 _23421_ ( .A1(_09087_ ), .A2(_10842_ ), .A3(fanout_net_5 ), .ZN(_02731_ ) );
MUX2_X1 _23422_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B ), .B(_02115_ ), .S(_01541_ ), .Z(_02732_ ) );
NAND2_X1 _23423_ ( .A1(_02732_ ), .A2(_01567_ ), .ZN(_02733_ ) );
NAND2_X1 _23424_ ( .A1(_02416_ ), .A2(_01562_ ), .ZN(_02734_ ) );
OAI211_X1 _23425_ ( .A(_01899_ ), .B(_02549_ ), .C1(_01891_ ), .C2(_01642_ ), .ZN(_02735_ ) );
AND3_X1 _23426_ ( .A1(_01900_ ), .A2(_01902_ ), .A3(_01261_ ), .ZN(_02736_ ) );
AOI21_X1 _23427_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B1(_01900_ ), .B2(_01902_ ), .ZN(_02737_ ) );
OAI21_X1 _23428_ ( .A(_01888_ ), .B1(_02736_ ), .B2(_02737_ ), .ZN(_02738_ ) );
NAND3_X1 _23429_ ( .A1(_02735_ ), .A2(_02738_ ), .A3(_01547_ ), .ZN(_02739_ ) );
NAND3_X1 _23430_ ( .A1(_02734_ ), .A2(_01541_ ), .A3(_02739_ ), .ZN(_02740_ ) );
OAI211_X1 _23431_ ( .A(_02740_ ), .B(_01879_ ), .C1(_02110_ ), .C2(_01564_ ), .ZN(_02741_ ) );
AND3_X1 _23432_ ( .A1(_02733_ ), .A2(_01530_ ), .A3(_02741_ ), .ZN(_02742_ ) );
NOR3_X1 _23433_ ( .A1(_09088_ ), .A2(fanout_net_27 ), .A3(_02023_ ), .ZN(_02743_ ) );
NAND2_X1 _23434_ ( .A1(_02429_ ), .A2(_01770_ ), .ZN(_02744_ ) );
OAI21_X1 _23435_ ( .A(_01781_ ), .B1(_02561_ ), .B2(_02564_ ), .ZN(_02745_ ) );
AND3_X1 _23436_ ( .A1(_01922_ ), .A2(_01923_ ), .A3(_01261_ ), .ZN(_02746_ ) );
AOI21_X1 _23437_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B1(_01922_ ), .B2(_01923_ ), .ZN(_02747_ ) );
OAI21_X1 _23438_ ( .A(_01763_ ), .B1(_02746_ ), .B2(_02747_ ), .ZN(_02748_ ) );
NAND3_X1 _23439_ ( .A1(_02745_ ), .A2(_02748_ ), .A3(_01589_ ), .ZN(_02749_ ) );
AND3_X1 _23440_ ( .A1(_02744_ ), .A2(_01204_ ), .A3(_02749_ ), .ZN(_02750_ ) );
NOR3_X1 _23441_ ( .A1(_02123_ ), .A2(_02126_ ), .A3(_01591_ ), .ZN(_02751_ ) );
OAI21_X1 _23442_ ( .A(_01211_ ), .B1(_02750_ ), .B2(_02751_ ), .ZN(_02752_ ) );
NAND3_X1 _23443_ ( .A1(_02132_ ), .A2(_01205_ ), .A3(_01793_ ), .ZN(_02753_ ) );
AOI21_X1 _23444_ ( .A(_01797_ ), .B1(_02752_ ), .B2(_02753_ ), .ZN(_02754_ ) );
OR3_X1 _23445_ ( .A1(_01635_ ), .A2(_01270_ ), .A3(_01241_ ), .ZN(_02755_ ) );
OAI21_X1 _23446_ ( .A(_02755_ ), .B1(_02142_ ), .B2(_01246_ ), .ZN(_02756_ ) );
AND3_X1 _23447_ ( .A1(_02756_ ), .A2(_02355_ ), .A3(_01337_ ), .ZN(_02757_ ) );
NAND2_X1 _23448_ ( .A1(_10209_ ), .A2(_01459_ ), .ZN(_02758_ ) );
NAND4_X1 _23449_ ( .A1(_01465_ ), .A2(\exu.addi.io_imm [10] ), .A3(_01462_ ), .A4(_01467_ ), .ZN(_02759_ ) );
AOI21_X1 _23450_ ( .A(\exu.io_in_bits_sub ), .B1(_02758_ ), .B2(_02759_ ), .ZN(_02760_ ) );
AND3_X1 _23451_ ( .A1(_02368_ ), .A2(_08705_ ), .A3(_08846_ ), .ZN(_02761_ ) );
NOR3_X1 _23452_ ( .A1(_02761_ ), .A2(_02686_ ), .A3(_01596_ ), .ZN(_02762_ ) );
OAI21_X1 _23453_ ( .A(_01452_ ), .B1(_02760_ ), .B2(_02762_ ), .ZN(_02763_ ) );
NAND2_X1 _23454_ ( .A1(_02752_ ), .A2(_02753_ ), .ZN(_02764_ ) );
NAND2_X1 _23455_ ( .A1(_02764_ ), .A2(_01593_ ), .ZN(_02765_ ) );
AOI21_X1 _23456_ ( .A(\exu.io_in_bits_or ), .B1(_02763_ ), .B2(_02765_ ), .ZN(_02766_ ) );
NOR3_X1 _23457_ ( .A1(_02709_ ), .A2(fanout_net_27 ), .A3(_02512_ ), .ZN(_02767_ ) );
OAI21_X1 _23458_ ( .A(_01443_ ), .B1(_02766_ ), .B2(_02767_ ), .ZN(_02768_ ) );
NAND3_X1 _23459_ ( .A1(_02733_ ), .A2(_01444_ ), .A3(_02741_ ), .ZN(_02769_ ) );
AOI21_X1 _23460_ ( .A(fanout_net_4 ), .B1(_02768_ ), .B2(_02769_ ), .ZN(_02770_ ) );
AND3_X1 _23461_ ( .A1(_01376_ ), .A2(_09462_ ), .A3(fanout_net_4 ), .ZN(_02771_ ) );
OR2_X1 _23462_ ( .A1(_02770_ ), .A2(_02771_ ), .ZN(_02772_ ) );
AOI221_X4 _23463_ ( .A(fanout_net_12 ), .B1(_08705_ ), .B2(_01492_ ), .C1(_02772_ ), .C2(_01617_ ), .ZN(_02773_ ) );
NAND3_X1 _23464_ ( .A1(_02756_ ), .A2(_01333_ ), .A3(_01440_ ), .ZN(_02774_ ) );
AOI211_X1 _23465_ ( .A(_01573_ ), .B(_02773_ ), .C1(fanout_net_12 ), .C2(_02774_ ), .ZN(_02775_ ) );
XNOR2_X1 _23466_ ( .A(_02708_ ), .B(_08705_ ), .ZN(_02776_ ) );
AND2_X1 _23467_ ( .A1(_02776_ ), .A2(_01436_ ), .ZN(_02777_ ) );
OAI21_X1 _23468_ ( .A(_09410_ ), .B1(_02775_ ), .B2(_02777_ ), .ZN(_02778_ ) );
OAI21_X1 _23469_ ( .A(_02778_ ), .B1(_01342_ ), .B2(_10217_ ), .ZN(_02779_ ) );
NAND2_X1 _23470_ ( .A1(_02779_ ), .A2(_01340_ ), .ZN(_02780_ ) );
NAND2_X1 _23471_ ( .A1(_10212_ ), .A2(_09460_ ), .ZN(_02781_ ) );
AOI21_X1 _23472_ ( .A(\exu.io_out_bits_ren ), .B1(_02780_ ), .B2(_02781_ ), .ZN(_02782_ ) );
MUX2_X1 _23473_ ( .A(_02757_ ), .B(_02782_ ), .S(_01504_ ), .Z(_02783_ ) );
MUX2_X1 _23474_ ( .A(_02754_ ), .B(_02783_ ), .S(_01214_ ), .Z(_02784_ ) );
MUX2_X1 _23475_ ( .A(_02743_ ), .B(_02784_ ), .S(_01509_ ), .Z(_02785_ ) );
MUX2_X1 _23476_ ( .A(_02742_ ), .B(_02785_ ), .S(_01181_ ), .Z(_02786_ ) );
MUX2_X1 _23477_ ( .A(_02731_ ), .B(_02786_ ), .S(_01515_ ), .Z(_02787_ ) );
NAND2_X1 _23478_ ( .A1(_02787_ ), .A2(_01723_ ), .ZN(_02788_ ) );
NAND2_X1 _23479_ ( .A1(_09089_ ), .A2(_01867_ ), .ZN(_02789_ ) );
AOI21_X1 _23480_ ( .A(_01722_ ), .B1(_02788_ ), .B2(_02789_ ), .ZN(_02790_ ) );
NOR3_X1 _23481_ ( .A1(_10242_ ), .A2(_10243_ ), .A3(_02249_ ), .ZN(_02791_ ) );
OAI21_X1 _23482_ ( .A(_01109_ ), .B1(_02790_ ), .B2(_02791_ ), .ZN(_02792_ ) );
OAI211_X1 _23483_ ( .A(_01873_ ), .B(\exu.csrrs.io_csr_rdata [10] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_02793_ ) );
NAND2_X1 _23484_ ( .A1(_02792_ ), .A2(_02793_ ), .ZN(\exu.io_out_bits_rd_wdata [10] ) );
NAND3_X1 _23485_ ( .A1(_02257_ ), .A2(_02258_ ), .A3(_01642_ ), .ZN(_02794_ ) );
OAI211_X1 _23486_ ( .A(_01725_ ), .B(_02794_ ), .C1(_01890_ ), .C2(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02795_ ) );
NAND3_X1 _23487_ ( .A1(_02257_ ), .A2(_02258_ ), .A3(_01263_ ), .ZN(_02796_ ) );
OAI211_X1 _23488_ ( .A(_01887_ ), .B(_02796_ ), .C1(_01890_ ), .C2(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02797_ ) );
AND3_X1 _23489_ ( .A1(_02795_ ), .A2(_02797_ ), .A3(_01546_ ), .ZN(_02798_ ) );
AOI21_X1 _23490_ ( .A(_01546_ ), .B1(_02474_ ), .B2(_02476_ ), .ZN(_02799_ ) );
NOR2_X1 _23491_ ( .A1(_02798_ ), .A2(_02799_ ), .ZN(_02800_ ) );
MUX2_X1 _23492_ ( .A(_02800_ ), .B(_02188_ ), .S(_01748_ ), .Z(_02801_ ) );
MUX2_X1 _23493_ ( .A(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B ), .B(_02190_ ), .S(_01564_ ), .Z(_02802_ ) );
MUX2_X1 _23494_ ( .A(_02801_ ), .B(_02802_ ), .S(_01567_ ), .Z(_02803_ ) );
OR2_X1 _23495_ ( .A1(_02803_ ), .A2(_01751_ ), .ZN(_02804_ ) );
INV_X1 _23496_ ( .A(_02220_ ), .ZN(_02805_ ) );
MUX2_X1 _23497_ ( .A(_02224_ ), .B(_02805_ ), .S(_01246_ ), .Z(_02806_ ) );
OR3_X1 _23498_ ( .A1(_02806_ ), .A2(_01654_ ), .A3(_02572_ ), .ZN(_02807_ ) );
NAND3_X1 _23499_ ( .A1(_02200_ ), .A2(_01935_ ), .A3(_02205_ ), .ZN(_02808_ ) );
AND3_X1 _23500_ ( .A1(_01758_ ), .A2(_01759_ ), .A3(_01263_ ), .ZN(_02809_ ) );
AOI21_X1 _23501_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_01190_ ), .B2(_01193_ ), .ZN(_02810_ ) );
NOR2_X1 _23502_ ( .A1(_02809_ ), .A2(_02810_ ), .ZN(_02811_ ) );
NAND2_X1 _23503_ ( .A1(_02811_ ), .A2(_01763_ ), .ZN(_02812_ ) );
OAI21_X1 _23504_ ( .A(_01781_ ), .B1(_02673_ ), .B2(_02674_ ), .ZN(_02813_ ) );
AND3_X1 _23505_ ( .A1(_02812_ ), .A2(_01589_ ), .A3(_02813_ ), .ZN(_02814_ ) );
AOI21_X1 _23506_ ( .A(_01589_ ), .B1(_02487_ ), .B2(_02490_ ), .ZN(_02815_ ) );
NOR2_X1 _23507_ ( .A1(_02814_ ), .A2(_02815_ ), .ZN(_02816_ ) );
OAI211_X1 _23508_ ( .A(_02808_ ), .B(_01450_ ), .C1(_02816_ ), .C2(_01935_ ), .ZN(_02817_ ) );
AND3_X1 _23509_ ( .A1(_02197_ ), .A2(_01206_ ), .A3(_02198_ ), .ZN(_02818_ ) );
OAI21_X1 _23510_ ( .A(_02817_ ), .B1(_02818_ ), .B2(_01450_ ), .ZN(_02819_ ) );
NOR2_X1 _23511_ ( .A1(_02819_ ), .A2(_01455_ ), .ZN(_02820_ ) );
AND4_X1 _23512_ ( .A1(\exu.addi.io_imm [9] ), .A2(_01465_ ), .A3(_01462_ ), .A4(_01467_ ), .ZN(_02821_ ) );
AOI21_X1 _23513_ ( .A(_02821_ ), .B1(_10257_ ), .B2(_01606_ ), .ZN(_02822_ ) );
OR2_X1 _23514_ ( .A1(_02822_ ), .A2(\exu.io_in_bits_sub ), .ZN(_02823_ ) );
OR3_X1 _23515_ ( .A1(_02366_ ), .A2(_08713_ ), .A3(_08842_ ), .ZN(_02824_ ) );
OAI211_X1 _23516_ ( .A(_02824_ ), .B(_01478_ ), .C1(_08712_ ), .C2(_08843_ ), .ZN(_02825_ ) );
OAI21_X1 _23517_ ( .A(_02823_ ), .B1(_02367_ ), .B2(_02825_ ), .ZN(_02826_ ) );
AOI21_X1 _23518_ ( .A(_02820_ ), .B1(_02826_ ), .B2(_01610_ ), .ZN(_02827_ ) );
OAI221_X1 _23519_ ( .A(_01613_ ), .B1(_08711_ ), .B2(_01832_ ), .C1(_02827_ ), .C2(\exu.io_in_bits_or ), .ZN(_02828_ ) );
NOR2_X1 _23520_ ( .A1(_02803_ ), .A2(_01579_ ), .ZN(_02829_ ) );
OAI211_X1 _23521_ ( .A(_02828_ ), .B(_01486_ ), .C1(_01614_ ), .C2(_02829_ ), .ZN(_02830_ ) );
NAND3_X1 _23522_ ( .A1(_08710_ ), .A2(_01575_ ), .A3(\exu.and_.io_is ), .ZN(_02831_ ) );
AOI21_X1 _23523_ ( .A(\exu.io_in_bits_xor ), .B1(_02830_ ), .B2(_02831_ ), .ZN(_02832_ ) );
AOI211_X1 _23524_ ( .A(fanout_net_12 ), .B(_02832_ ), .C1(_08712_ ), .C2(_01493_ ), .ZN(_02833_ ) );
OR3_X1 _23525_ ( .A1(_02806_ ), .A2(_01804_ ), .A3(_02589_ ), .ZN(_02834_ ) );
AOI211_X1 _23526_ ( .A(_01573_ ), .B(_02833_ ), .C1(fanout_net_12 ), .C2(_02834_ ), .ZN(_02835_ ) );
NOR2_X1 _23527_ ( .A1(_02384_ ), .A2(_08715_ ), .ZN(_02836_ ) );
NOR2_X1 _23528_ ( .A1(_02836_ ), .A2(_01380_ ), .ZN(_02837_ ) );
XNOR2_X1 _23529_ ( .A(_02837_ ), .B(_08712_ ), .ZN(_02838_ ) );
AOI21_X1 _23530_ ( .A(_02835_ ), .B1(_01828_ ), .B2(_02838_ ), .ZN(_02839_ ) );
OAI221_X1 _23531_ ( .A(_01341_ ), .B1(_01823_ ), .B2(_10262_ ), .C1(_02839_ ), .C2(\exu.io_in_bits_jal ), .ZN(_02840_ ) );
NOR2_X1 _23532_ ( .A1(_10262_ ), .A2(_01855_ ), .ZN(_02841_ ) );
OAI211_X1 _23533_ ( .A(_02840_ ), .B(_01501_ ), .C1(_01854_ ), .C2(_02841_ ), .ZN(_02842_ ) );
MUX2_X1 _23534_ ( .A(_02807_ ), .B(_02842_ ), .S(_01992_ ), .Z(_02843_ ) );
NAND2_X1 _23535_ ( .A1(_02843_ ), .A2(_01705_ ), .ZN(_02844_ ) );
NOR2_X1 _23536_ ( .A1(_02819_ ), .A2(_01797_ ), .ZN(_02845_ ) );
OAI211_X1 _23537_ ( .A(_02844_ ), .B(_01510_ ), .C1(_01994_ ), .C2(_02845_ ), .ZN(_02846_ ) );
AOI21_X1 _23538_ ( .A(\exu.io_in_bits_srai ), .B1(_09095_ ), .B2(_01186_ ), .ZN(_02847_ ) );
AOI221_X4 _23539_ ( .A(fanout_net_5 ), .B1(\exu.io_in_bits_srai ), .B2(_02804_ ), .C1(_02846_ ), .C2(_02847_ ), .ZN(_02848_ ) );
AND3_X1 _23540_ ( .A1(_09083_ ), .A2(_01864_ ), .A3(fanout_net_5 ), .ZN(_02849_ ) );
OAI21_X1 _23541_ ( .A(_01723_ ), .B1(_02848_ ), .B2(_02849_ ), .ZN(_02850_ ) );
NAND2_X1 _23542_ ( .A1(_09085_ ), .A2(_01867_ ), .ZN(_02851_ ) );
AOI21_X1 _23543_ ( .A(_01722_ ), .B1(_02850_ ), .B2(_02851_ ), .ZN(_02852_ ) );
AND2_X1 _23544_ ( .A1(\exu.addi._io_rd_T_4 [9] ), .A2(_01870_ ), .ZN(_02853_ ) );
OAI21_X1 _23545_ ( .A(_01109_ ), .B1(_02852_ ), .B2(_02853_ ), .ZN(_02854_ ) );
OAI211_X1 _23546_ ( .A(_01873_ ), .B(\exu.csrrs.io_csr_rdata [9] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_02855_ ) );
NAND2_X1 _23547_ ( .A1(_02854_ ), .A2(_02855_ ), .ZN(\exu.io_out_bits_rd_wdata [9] ) );
AND3_X1 _23548_ ( .A1(_09080_ ), .A2(_10843_ ), .A3(fanout_net_5 ), .ZN(_02856_ ) );
AOI21_X1 _23549_ ( .A(_01564_ ), .B1(_02255_ ), .B2(_02263_ ), .ZN(_02857_ ) );
OR3_X1 _23550_ ( .A1(_02736_ ), .A2(_02737_ ), .A3(_01559_ ), .ZN(_02858_ ) );
NAND3_X1 _23551_ ( .A1(_01901_ ), .A2(_01903_ ), .A3(_01267_ ), .ZN(_02859_ ) );
OAI211_X1 _23552_ ( .A(_01887_ ), .B(_02859_ ), .C1(_01891_ ), .C2(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02860_ ) );
AND3_X1 _23553_ ( .A1(_02858_ ), .A2(_02860_ ), .A3(_01547_ ), .ZN(_02861_ ) );
AOI21_X1 _23554_ ( .A(_01547_ ), .B1(_02548_ ), .B2(_02550_ ), .ZN(_02862_ ) );
NOR3_X1 _23555_ ( .A1(_02861_ ), .A2(_02862_ ), .A3(_01747_ ), .ZN(_02863_ ) );
OAI21_X1 _23556_ ( .A(_01879_ ), .B1(_02857_ ), .B2(_02863_ ), .ZN(_02864_ ) );
AOI21_X1 _23557_ ( .A(_01542_ ), .B1(_02266_ ), .B2(_01564_ ), .ZN(_02865_ ) );
OAI21_X1 _23558_ ( .A(_02864_ ), .B1(_02865_ ), .B2(_01879_ ), .ZN(_02866_ ) );
NOR2_X1 _23559_ ( .A1(_02866_ ), .A2(_01752_ ), .ZN(_02867_ ) );
NOR3_X1 _23560_ ( .A1(_09081_ ), .A2(fanout_net_27 ), .A3(_01509_ ), .ZN(_02868_ ) );
NAND3_X1 _23561_ ( .A1(_02273_ ), .A2(_01206_ ), .A3(_01794_ ), .ZN(_02869_ ) );
AOI21_X1 _23562_ ( .A(_01590_ ), .B1(_02560_ ), .B2(_02565_ ), .ZN(_02870_ ) );
NAND3_X1 _23563_ ( .A1(_02562_ ), .A2(_02563_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02871_ ) );
OAI211_X1 _23564_ ( .A(_01778_ ), .B(_02871_ ), .C1(_01767_ ), .C2(_01648_ ), .ZN(_02872_ ) );
OAI21_X1 _23565_ ( .A(_01587_ ), .B1(_02746_ ), .B2(_02747_ ), .ZN(_02873_ ) );
AOI21_X1 _23566_ ( .A(_01771_ ), .B1(_02872_ ), .B2(_02873_ ), .ZN(_02874_ ) );
NOR2_X1 _23567_ ( .A1(_02870_ ), .A2(_02874_ ), .ZN(_02875_ ) );
MUX2_X1 _23568_ ( .A(_02875_ ), .B(_02281_ ), .S(_01790_ ), .Z(_02876_ ) );
OAI21_X1 _23569_ ( .A(_02869_ ), .B1(_02876_ ), .B2(_01794_ ), .ZN(_02877_ ) );
AND2_X1 _23570_ ( .A1(_02877_ ), .A2(_01217_ ), .ZN(_02878_ ) );
NAND4_X1 _23571_ ( .A1(_01279_ ), .A2(_01299_ ), .A3(_01634_ ), .A4(_01246_ ), .ZN(_02879_ ) );
OAI21_X1 _23572_ ( .A(_02879_ ), .B1(_02289_ ), .B2(_01246_ ), .ZN(_02880_ ) );
AND3_X1 _23573_ ( .A1(_02880_ ), .A2(_02355_ ), .A3(_01337_ ), .ZN(_02881_ ) );
NAND3_X1 _23574_ ( .A1(_02880_ ), .A2(_01333_ ), .A3(_01440_ ), .ZN(_02882_ ) );
NAND2_X1 _23575_ ( .A1(_02877_ ), .A2(_01593_ ), .ZN(_02883_ ) );
OAI21_X1 _23576_ ( .A(_01477_ ), .B1(_02365_ ), .B2(_08714_ ), .ZN(_02884_ ) );
AOI21_X1 _23577_ ( .A(_02884_ ), .B1(_08714_ ), .B2(_02365_ ), .ZN(_02885_ ) );
NAND4_X1 _23578_ ( .A1(_01600_ ), .A2(\exu.addi.io_imm [8] ), .A3(_01463_ ), .A4(_01603_ ), .ZN(_02886_ ) );
OAI21_X1 _23579_ ( .A(_02886_ ), .B1(_10528_ ), .B2(_01460_ ), .ZN(_02887_ ) );
AOI21_X1 _23580_ ( .A(_02885_ ), .B1(_02887_ ), .B2(_01457_ ), .ZN(_02888_ ) );
OAI21_X1 _23581_ ( .A(_02883_ ), .B1(_02888_ ), .B2(\exu.io_in_bits_srl ), .ZN(_02889_ ) );
NAND2_X1 _23582_ ( .A1(_02889_ ), .A2(_02512_ ), .ZN(_02890_ ) );
OAI21_X1 _23583_ ( .A(_01448_ ), .B1(\exu.add.io_rs1_data [8] ), .B2(\exu._GEN_0 [8] ), .ZN(_02891_ ) );
AOI21_X1 _23584_ ( .A(\exu.io_in_bits_sra ), .B1(_02890_ ), .B2(_02891_ ), .ZN(_02892_ ) );
NOR2_X1 _23585_ ( .A1(_02866_ ), .A2(_01578_ ), .ZN(_02893_ ) );
OAI21_X1 _23586_ ( .A(_01486_ ), .B1(_02892_ ), .B2(_02893_ ), .ZN(_02894_ ) );
NAND3_X1 _23587_ ( .A1(_01380_ ), .A2(_10698_ ), .A3(\exu.and_.io_is ), .ZN(_02895_ ) );
AOI21_X1 _23588_ ( .A(\exu.io_in_bits_xor ), .B1(_02894_ ), .B2(_02895_ ), .ZN(_02896_ ) );
AOI21_X1 _23589_ ( .A(_02896_ ), .B1(_08714_ ), .B2(_01968_ ), .ZN(_02897_ ) );
OAI21_X1 _23590_ ( .A(_02882_ ), .B1(_02897_ ), .B2(fanout_net_12 ), .ZN(_02898_ ) );
AND2_X1 _23591_ ( .A1(_02898_ ), .A2(_01498_ ), .ZN(_02899_ ) );
OAI21_X1 _23592_ ( .A(_01436_ ), .B1(_02384_ ), .B2(_08715_ ), .ZN(_02900_ ) );
AOI21_X1 _23593_ ( .A(_02900_ ), .B1(_08715_ ), .B2(_02384_ ), .ZN(_02901_ ) );
OAI21_X1 _23594_ ( .A(_09410_ ), .B1(_02899_ ), .B2(_02901_ ), .ZN(_02902_ ) );
OAI21_X1 _23595_ ( .A(_02902_ ), .B1(_01342_ ), .B2(_10530_ ), .ZN(_02903_ ) );
NAND2_X1 _23596_ ( .A1(_02903_ ), .A2(_01340_ ), .ZN(_02904_ ) );
NAND2_X1 _23597_ ( .A1(_10525_ ), .A2(_09460_ ), .ZN(_02905_ ) );
AOI21_X1 _23598_ ( .A(\exu.io_out_bits_ren ), .B1(_02904_ ), .B2(_02905_ ), .ZN(_02906_ ) );
MUX2_X1 _23599_ ( .A(_02881_ ), .B(_02906_ ), .S(_01504_ ), .Z(_02907_ ) );
MUX2_X1 _23600_ ( .A(_02878_ ), .B(_02907_ ), .S(_01507_ ), .Z(_02908_ ) );
MUX2_X1 _23601_ ( .A(_02868_ ), .B(_02908_ ), .S(_01509_ ), .Z(_02909_ ) );
MUX2_X1 _23602_ ( .A(_02867_ ), .B(_02909_ ), .S(_01182_ ), .Z(_02910_ ) );
MUX2_X1 _23603_ ( .A(_02856_ ), .B(_02910_ ), .S(_01878_ ), .Z(_02911_ ) );
NAND2_X1 _23604_ ( .A1(_02911_ ), .A2(_01877_ ), .ZN(_02912_ ) );
NAND2_X1 _23605_ ( .A1(_09082_ ), .A2(_02000_ ), .ZN(_02913_ ) );
AOI21_X1 _23606_ ( .A(_01876_ ), .B1(_02912_ ), .B2(_02913_ ), .ZN(_02914_ ) );
AND2_X1 _23607_ ( .A1(\exu.addi._io_rd_T_4 [8] ), .A2(_02003_ ), .ZN(_02915_ ) );
OAI21_X1 _23608_ ( .A(_01875_ ), .B1(_02914_ ), .B2(_02915_ ), .ZN(_02916_ ) );
OAI211_X1 _23609_ ( .A(_01058_ ), .B(\exu.csrrs.io_csr_rdata [8] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_02917_ ) );
NAND2_X1 _23610_ ( .A1(_02916_ ), .A2(_02917_ ), .ZN(\exu.io_out_bits_rd_wdata [8] ) );
AND3_X1 _23611_ ( .A1(_09077_ ), .A2(_10842_ ), .A3(fanout_net_5 ), .ZN(_02918_ ) );
NAND3_X1 _23612_ ( .A1(_02257_ ), .A2(_02258_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02919_ ) );
OAI211_X1 _23613_ ( .A(_01899_ ), .B(_02919_ ), .C1(_01890_ ), .C2(_01267_ ), .ZN(_02920_ ) );
INV_X1 _23614_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02921_ ) );
OR2_X1 _23615_ ( .A1(_01729_ ), .A2(_02921_ ), .ZN(_02922_ ) );
NAND3_X1 _23616_ ( .A1(_02257_ ), .A2(_02258_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02923_ ) );
NAND2_X1 _23617_ ( .A1(_02922_ ), .A2(_02923_ ), .ZN(_02924_ ) );
OAI211_X1 _23618_ ( .A(_01547_ ), .B(_02920_ ), .C1(_02924_ ), .C2(_01884_ ), .ZN(_02925_ ) );
NAND3_X1 _23619_ ( .A1(_02662_ ), .A2(_02664_ ), .A3(_01562_ ), .ZN(_02926_ ) );
AOI21_X1 _23620_ ( .A(_01747_ ), .B1(_02925_ ), .B2(_02926_ ), .ZN(_02927_ ) );
AOI21_X1 _23621_ ( .A(_02927_ ), .B1(_02334_ ), .B2(_01747_ ), .ZN(_02928_ ) );
AOI21_X1 _23622_ ( .A(_01542_ ), .B1(_02336_ ), .B2(_01541_ ), .ZN(_02929_ ) );
MUX2_X1 _23623_ ( .A(_02928_ ), .B(_02929_ ), .S(_01567_ ), .Z(_02930_ ) );
AND2_X1 _23624_ ( .A1(_02930_ ), .A2(_01914_ ), .ZN(_02931_ ) );
NOR3_X1 _23625_ ( .A1(_09079_ ), .A2(fanout_net_27 ), .A3(_02023_ ), .ZN(_02932_ ) );
MUX2_X1 _23626_ ( .A(_02351_ ), .B(_02349_ ), .S(_01204_ ), .Z(_02933_ ) );
NAND3_X1 _23627_ ( .A1(_02675_ ), .A2(_01770_ ), .A3(_02676_ ), .ZN(_02934_ ) );
OAI21_X1 _23628_ ( .A(_01586_ ), .B1(_02809_ ), .B2(_02810_ ), .ZN(_02935_ ) );
NAND3_X1 _23629_ ( .A1(_01190_ ), .A2(_01193_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02936_ ) );
OAI211_X1 _23630_ ( .A(_01197_ ), .B(_02936_ ), .C1(_01583_ ), .C2(_02921_ ), .ZN(_02937_ ) );
AND2_X1 _23631_ ( .A1(_02935_ ), .A2(_02937_ ), .ZN(_02938_ ) );
INV_X1 _23632_ ( .A(_02938_ ), .ZN(_02939_ ) );
OAI211_X1 _23633_ ( .A(_01204_ ), .B(_02934_ ), .C1(_02939_ ), .C2(_01770_ ), .ZN(_02940_ ) );
OAI21_X1 _23634_ ( .A(_01789_ ), .B1(_02344_ ), .B2(_02345_ ), .ZN(_02941_ ) );
AND2_X1 _23635_ ( .A1(_02940_ ), .A2(_02941_ ), .ZN(_02942_ ) );
MUX2_X1 _23636_ ( .A(_02933_ ), .B(_02942_ ), .S(_01210_ ), .Z(_02943_ ) );
NOR2_X1 _23637_ ( .A1(_02943_ ), .A2(_01797_ ), .ZN(_02944_ ) );
AND3_X1 _23638_ ( .A1(_01242_ ), .A2(_01270_ ), .A3(_01259_ ), .ZN(_02945_ ) );
AND3_X1 _23639_ ( .A1(_02945_ ), .A2(_02354_ ), .A3(_01337_ ), .ZN(_02946_ ) );
NAND3_X1 _23640_ ( .A1(_08728_ ), .A2(_09463_ ), .A3(\exu.and_.io_is ), .ZN(_02947_ ) );
OR2_X1 _23641_ ( .A1(_02943_ ), .A2(_01454_ ), .ZN(_02948_ ) );
AOI21_X1 _23642_ ( .A(_08838_ ), .B1(_08829_ ), .B2(_08736_ ), .ZN(_02949_ ) );
NOR2_X1 _23643_ ( .A1(_02949_ ), .A2(_08727_ ), .ZN(_02950_ ) );
AOI21_X1 _23644_ ( .A(_02950_ ), .B1(\exu.add.io_rs1_data [6] ), .B2(_12841_ ), .ZN(_02951_ ) );
OAI21_X1 _23645_ ( .A(_01477_ ), .B1(_02951_ ), .B2(_08730_ ), .ZN(_02952_ ) );
AOI21_X1 _23646_ ( .A(_02952_ ), .B1(_08730_ ), .B2(_02951_ ), .ZN(_02953_ ) );
NAND4_X1 _23647_ ( .A1(_01465_ ), .A2(\exu.addi.io_imm [7] ), .A3(_01462_ ), .A4(_01467_ ), .ZN(_02954_ ) );
OAI21_X1 _23648_ ( .A(_02954_ ), .B1(_10488_ ), .B2(_01460_ ), .ZN(_02955_ ) );
AOI21_X1 _23649_ ( .A(_02953_ ), .B1(_02955_ ), .B2(_01457_ ), .ZN(_02956_ ) );
OAI21_X1 _23650_ ( .A(_02948_ ), .B1(_02956_ ), .B2(\exu.io_in_bits_srl ), .ZN(_02957_ ) );
NAND2_X1 _23651_ ( .A1(_02957_ ), .A2(_02512_ ), .ZN(_02958_ ) );
OAI21_X1 _23652_ ( .A(_01447_ ), .B1(\exu.add.io_rs1_data [7] ), .B2(\exu._GEN_0 [7] ), .ZN(_02959_ ) );
AOI21_X1 _23653_ ( .A(\exu.io_in_bits_sra ), .B1(_02958_ ), .B2(_02959_ ), .ZN(_02960_ ) );
AOI21_X1 _23654_ ( .A(_02960_ ), .B1(_01444_ ), .B2(_02930_ ), .ZN(_02961_ ) );
OAI21_X1 _23655_ ( .A(_02947_ ), .B1(_02961_ ), .B2(\exu.and_.io_is ), .ZN(_02962_ ) );
AOI221_X4 _23656_ ( .A(\exu.io_in_bits_sll ), .B1(_08730_ ), .B2(_01492_ ), .C1(_02962_ ), .C2(_01617_ ), .ZN(_02963_ ) );
NAND3_X1 _23657_ ( .A1(_02945_ ), .A2(_01333_ ), .A3(_01440_ ), .ZN(_02964_ ) );
AOI211_X1 _23658_ ( .A(_01572_ ), .B(_02963_ ), .C1(\exu.io_in_bits_sll ), .C2(_02964_ ), .ZN(_02965_ ) );
XNOR2_X1 _23659_ ( .A(_01372_ ), .B(_08730_ ), .ZN(_02966_ ) );
AND2_X1 _23660_ ( .A1(_02966_ ), .A2(_01436_ ), .ZN(_02967_ ) );
OAI21_X1 _23661_ ( .A(_09410_ ), .B1(_02965_ ), .B2(_02967_ ), .ZN(_02968_ ) );
OAI21_X1 _23662_ ( .A(_02968_ ), .B1(_01342_ ), .B2(_10480_ ), .ZN(_02969_ ) );
NAND2_X1 _23663_ ( .A1(_02969_ ), .A2(_01340_ ), .ZN(_02970_ ) );
OR2_X1 _23664_ ( .A1(_10480_ ), .A2(_01855_ ), .ZN(_02971_ ) );
AOI21_X1 _23665_ ( .A(\exu.io_out_bits_ren ), .B1(_02970_ ), .B2(_02971_ ), .ZN(_02972_ ) );
MUX2_X1 _23666_ ( .A(_02946_ ), .B(_02972_ ), .S(_01504_ ), .Z(_02973_ ) );
MUX2_X1 _23667_ ( .A(_02944_ ), .B(_02973_ ), .S(_01214_ ), .Z(_02974_ ) );
MUX2_X1 _23668_ ( .A(_02932_ ), .B(_02974_ ), .S(_02023_ ), .Z(_02975_ ) );
MUX2_X1 _23669_ ( .A(_02931_ ), .B(_02975_ ), .S(_01181_ ), .Z(_02976_ ) );
MUX2_X1 _23670_ ( .A(_02918_ ), .B(_02976_ ), .S(_01515_ ), .Z(_02977_ ) );
NAND2_X1 _23671_ ( .A1(_02977_ ), .A2(_01723_ ), .ZN(_02978_ ) );
NAND2_X1 _23672_ ( .A1(_10514_ ), .A2(_01867_ ), .ZN(_02979_ ) );
AOI21_X1 _23673_ ( .A(_01722_ ), .B1(_02978_ ), .B2(_02979_ ), .ZN(_02980_ ) );
AND2_X1 _23674_ ( .A1(\exu.addi._io_rd_T_4 [7] ), .A2(_01870_ ), .ZN(_02981_ ) );
OAI21_X1 _23675_ ( .A(_01109_ ), .B1(_02980_ ), .B2(_02981_ ), .ZN(_02982_ ) );
OAI211_X1 _23676_ ( .A(_01873_ ), .B(\exu.csrrs.io_csr_rdata [7] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_02983_ ) );
NAND2_X1 _23677_ ( .A1(_02982_ ), .A2(_02983_ ), .ZN(\exu.io_out_bits_rd_wdata [7] ) );
AND3_X1 _23678_ ( .A1(_09074_ ), .A2(_10843_ ), .A3(fanout_net_5 ), .ZN(_02984_ ) );
OR3_X1 _23679_ ( .A1(_02409_ ), .A2(_01748_ ), .A3(_02410_ ), .ZN(_02985_ ) );
OAI211_X1 _23680_ ( .A(_02985_ ), .B(_01567_ ), .C1(_01881_ ), .C2(_01563_ ), .ZN(_02986_ ) );
NAND3_X1 _23681_ ( .A1(_01901_ ), .A2(_01903_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02987_ ) );
OAI211_X1 _23682_ ( .A(_01884_ ), .B(_02987_ ), .C1(_01891_ ), .C2(_01648_ ), .ZN(_02988_ ) );
NAND3_X1 _23683_ ( .A1(_01901_ ), .A2(_01903_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02989_ ) );
OAI211_X1 _23684_ ( .A(_01888_ ), .B(_02989_ ), .C1(_01891_ ), .C2(_01255_ ), .ZN(_02990_ ) );
AOI21_X1 _23685_ ( .A(_01882_ ), .B1(_02988_ ), .B2(_02990_ ), .ZN(_02991_ ) );
AOI21_X1 _23686_ ( .A(_01734_ ), .B1(_02735_ ), .B2(_02738_ ), .ZN(_02992_ ) );
OAI21_X1 _23687_ ( .A(_01881_ ), .B1(_02991_ ), .B2(_02992_ ), .ZN(_02993_ ) );
OAI211_X1 _23688_ ( .A(_02993_ ), .B(_01880_ ), .C1(_01881_ ), .C2(_02419_ ), .ZN(_02994_ ) );
AND3_X1 _23689_ ( .A1(_02986_ ), .A2(_01914_ ), .A3(_02994_ ), .ZN(_02995_ ) );
NOR3_X1 _23690_ ( .A1(_09075_ ), .A2(fanout_net_27 ), .A3(_01509_ ), .ZN(_02996_ ) );
AOI21_X1 _23691_ ( .A(_01788_ ), .B1(_02745_ ), .B2(_02748_ ), .ZN(_02997_ ) );
OAI211_X1 _23692_ ( .A(_01587_ ), .B(_02871_ ), .C1(_01767_ ), .C2(_01648_ ), .ZN(_02998_ ) );
NAND3_X1 _23693_ ( .A1(_02562_ ), .A2(_02563_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02999_ ) );
OAI211_X1 _23694_ ( .A(_01778_ ), .B(_02999_ ), .C1(_01767_ ), .C2(_01255_ ), .ZN(_03000_ ) );
NAND2_X1 _23695_ ( .A1(_02998_ ), .A2(_03000_ ), .ZN(_03001_ ) );
AOI211_X1 _23696_ ( .A(_01790_ ), .B(_02997_ ), .C1(_03001_ ), .C2(_01788_ ), .ZN(_03002_ ) );
AOI21_X1 _23697_ ( .A(_01206_ ), .B1(_02430_ ), .B2(_02431_ ), .ZN(_03003_ ) );
OAI21_X1 _23698_ ( .A(_01450_ ), .B1(_03002_ ), .B2(_03003_ ), .ZN(_03004_ ) );
NAND3_X1 _23699_ ( .A1(_01588_ ), .A2(_01788_ ), .A3(_01935_ ), .ZN(_03005_ ) );
OAI211_X1 _23700_ ( .A(_03005_ ), .B(_01794_ ), .C1(_01935_ ), .C2(_02435_ ), .ZN(_03006_ ) );
AND3_X1 _23701_ ( .A1(_03004_ ), .A2(_01217_ ), .A3(_03006_ ), .ZN(_03007_ ) );
AND3_X1 _23702_ ( .A1(_01628_ ), .A2(_01271_ ), .A3(_01636_ ), .ZN(_03008_ ) );
AND3_X1 _23703_ ( .A1(_03008_ ), .A2(_02355_ ), .A3(_01337_ ), .ZN(_03009_ ) );
NAND3_X1 _23704_ ( .A1(_03004_ ), .A2(_01594_ ), .A3(_03006_ ), .ZN(_03010_ ) );
OAI21_X1 _23705_ ( .A(_01478_ ), .B1(_02949_ ), .B2(_08727_ ), .ZN(_03011_ ) );
AOI21_X1 _23706_ ( .A(_03011_ ), .B1(_08727_ ), .B2(_02949_ ), .ZN(_03012_ ) );
NAND4_X1 _23707_ ( .A1(_01601_ ), .A2(\exu.addi.io_imm [6] ), .A3(_01602_ ), .A4(_01604_ ), .ZN(_03013_ ) );
OAI21_X1 _23708_ ( .A(_03013_ ), .B1(_10418_ ), .B2(_01460_ ), .ZN(_03014_ ) );
AOI21_X1 _23709_ ( .A(_03012_ ), .B1(_03014_ ), .B2(_01457_ ), .ZN(_03015_ ) );
OAI21_X1 _23710_ ( .A(_03010_ ), .B1(_03015_ ), .B2(\exu.io_in_bits_srl ), .ZN(_03016_ ) );
NAND2_X1 _23711_ ( .A1(_03016_ ), .A2(_02512_ ), .ZN(_03017_ ) );
OAI21_X1 _23712_ ( .A(_01581_ ), .B1(\exu.add.io_rs1_data [6] ), .B2(\exu._GEN_0 [6] ), .ZN(_03018_ ) );
AOI21_X1 _23713_ ( .A(\exu.io_in_bits_sra ), .B1(_03017_ ), .B2(_03018_ ), .ZN(_03019_ ) );
AND3_X1 _23714_ ( .A1(_02986_ ), .A2(_01445_ ), .A3(_02994_ ), .ZN(_03020_ ) );
OAI21_X1 _23715_ ( .A(_01486_ ), .B1(_03019_ ), .B2(_03020_ ), .ZN(_03021_ ) );
NAND3_X1 _23716_ ( .A1(_01371_ ), .A2(_01575_ ), .A3(\exu.and_.io_is ), .ZN(_03022_ ) );
AOI21_X1 _23717_ ( .A(\exu.io_in_bits_xor ), .B1(_03021_ ), .B2(_03022_ ), .ZN(_03023_ ) );
AND2_X1 _23718_ ( .A1(_08727_ ), .A2(_01492_ ), .ZN(_03024_ ) );
OAI21_X1 _23719_ ( .A(_01438_ ), .B1(_03023_ ), .B2(_03024_ ), .ZN(_03025_ ) );
NAND3_X1 _23720_ ( .A1(_03008_ ), .A2(_02354_ ), .A3(_01441_ ), .ZN(_03026_ ) );
AOI21_X1 _23721_ ( .A(_01573_ ), .B1(_03025_ ), .B2(_03026_ ), .ZN(_03027_ ) );
XNOR2_X1 _23722_ ( .A(_01368_ ), .B(_08727_ ), .ZN(_03028_ ) );
AND2_X1 _23723_ ( .A1(_03028_ ), .A2(_01436_ ), .ZN(_03029_ ) );
OAI21_X1 _23724_ ( .A(_01571_ ), .B1(_03027_ ), .B2(_03029_ ), .ZN(_03030_ ) );
OAI21_X1 _23725_ ( .A(_03030_ ), .B1(_01342_ ), .B2(_10400_ ), .ZN(_03031_ ) );
NAND2_X1 _23726_ ( .A1(_03031_ ), .A2(_01340_ ), .ZN(_03032_ ) );
NAND2_X1 _23727_ ( .A1(_10398_ ), .A2(_09460_ ), .ZN(_03033_ ) );
AOI21_X1 _23728_ ( .A(\exu.io_out_bits_ren ), .B1(_03032_ ), .B2(_03033_ ), .ZN(_03034_ ) );
MUX2_X1 _23729_ ( .A(_03009_ ), .B(_03034_ ), .S(_01505_ ), .Z(_03035_ ) );
MUX2_X1 _23730_ ( .A(_03007_ ), .B(_03035_ ), .S(_01507_ ), .Z(_03036_ ) );
MUX2_X1 _23731_ ( .A(_02996_ ), .B(_03036_ ), .S(_01509_ ), .Z(_03037_ ) );
MUX2_X1 _23732_ ( .A(_02995_ ), .B(_03037_ ), .S(_01182_ ), .Z(_03038_ ) );
MUX2_X1 _23733_ ( .A(_02984_ ), .B(_03038_ ), .S(_01878_ ), .Z(_03039_ ) );
NAND2_X1 _23734_ ( .A1(_03039_ ), .A2(_01877_ ), .ZN(_03040_ ) );
NAND2_X1 _23735_ ( .A1(_10425_ ), .A2(_02000_ ), .ZN(_03041_ ) );
AOI21_X1 _23736_ ( .A(_01876_ ), .B1(_03040_ ), .B2(_03041_ ), .ZN(_03042_ ) );
AND2_X1 _23737_ ( .A1(\exu.addi._io_rd_T_4 [6] ), .A2(_02003_ ), .ZN(_03043_ ) );
OAI21_X1 _23738_ ( .A(_01875_ ), .B1(_03042_ ), .B2(_03043_ ), .ZN(_03044_ ) );
OAI211_X1 _23739_ ( .A(_01058_ ), .B(\exu.csrrs.io_csr_rdata [6] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_03045_ ) );
NAND2_X1 _23740_ ( .A1(_03044_ ), .A2(_03045_ ), .ZN(\exu.io_out_bits_rd_wdata [6] ) );
AND3_X1 _23741_ ( .A1(_02478_ ), .A2(_02479_ ), .A3(_01748_ ), .ZN(_03046_ ) );
AND3_X1 _23742_ ( .A1(_02795_ ), .A2(_02797_ ), .A3(_01882_ ), .ZN(_03047_ ) );
AND3_X1 _23743_ ( .A1(_01900_ ), .A2(_01902_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03048_ ) );
AOI21_X1 _23744_ ( .A(_01249_ ), .B1(_02257_ ), .B2(_02258_ ), .ZN(_03049_ ) );
NOR2_X1 _23745_ ( .A1(_03048_ ), .A2(_03049_ ), .ZN(_03050_ ) );
NAND2_X1 _23746_ ( .A1(_03050_ ), .A2(_01888_ ), .ZN(_03051_ ) );
OAI211_X1 _23747_ ( .A(_01899_ ), .B(_02923_ ), .C1(_01891_ ), .C2(_02921_ ), .ZN(_03052_ ) );
NAND2_X1 _23748_ ( .A1(_03051_ ), .A2(_03052_ ), .ZN(_03053_ ) );
AOI211_X1 _23749_ ( .A(_01748_ ), .B(_03047_ ), .C1(_01734_ ), .C2(_03053_ ), .ZN(_03054_ ) );
OAI21_X1 _23750_ ( .A(_01880_ ), .B1(_03046_ ), .B2(_03054_ ), .ZN(_03055_ ) );
OAI211_X1 _23751_ ( .A(_01914_ ), .B(_03055_ ), .C1(_01749_ ), .C2(_02021_ ), .ZN(_03056_ ) );
AND3_X1 _23752_ ( .A1(_01803_ ), .A2(_02354_ ), .A3(_01686_ ), .ZN(_03057_ ) );
NAND2_X1 _23753_ ( .A1(_03057_ ), .A2(_01702_ ), .ZN(_03058_ ) );
OR2_X1 _23754_ ( .A1(_01792_ ), .A2(_01450_ ), .ZN(_03059_ ) );
OR3_X1 _23755_ ( .A1(_02491_ ), .A2(_01206_ ), .A3(_02492_ ), .ZN(_03060_ ) );
NAND3_X1 _23756_ ( .A1(_02812_ ), .A2(_01927_ ), .A3(_02813_ ), .ZN(_03061_ ) );
AND3_X1 _23757_ ( .A1(_02562_ ), .A2(_02563_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03062_ ) );
AOI21_X1 _23758_ ( .A(_01249_ ), .B1(_02562_ ), .B2(_02563_ ), .ZN(_03063_ ) );
NOR2_X1 _23759_ ( .A1(_03062_ ), .A2(_03063_ ), .ZN(_03064_ ) );
NAND2_X1 _23760_ ( .A1(_03064_ ), .A2(_01778_ ), .ZN(_03065_ ) );
OAI211_X1 _23761_ ( .A(_01781_ ), .B(_02936_ ), .C1(_01767_ ), .C2(_02921_ ), .ZN(_03066_ ) );
AND2_X1 _23762_ ( .A1(_03065_ ), .A2(_03066_ ), .ZN(_03067_ ) );
OAI211_X1 _23763_ ( .A(_01207_ ), .B(_03061_ ), .C1(_03067_ ), .C2(_01927_ ), .ZN(_03068_ ) );
NAND3_X1 _23764_ ( .A1(_03060_ ), .A2(_01212_ ), .A3(_03068_ ), .ZN(_03069_ ) );
AOI21_X1 _23765_ ( .A(_01455_ ), .B1(_03059_ ), .B2(_03069_ ), .ZN(_03070_ ) );
AOI211_X1 _23766_ ( .A(_08835_ ), .B(_01597_ ), .C1(_08829_ ), .C2(_08736_ ), .ZN(_03071_ ) );
AND2_X1 _23767_ ( .A1(_08829_ ), .A2(_01353_ ), .ZN(_03072_ ) );
OAI21_X1 _23768_ ( .A(_08735_ ), .B1(_08834_ ), .B2(\exu._GEN_0 [4] ), .ZN(_03073_ ) );
OAI21_X1 _23769_ ( .A(_03071_ ), .B1(_03072_ ), .B2(_03073_ ), .ZN(_03074_ ) );
AND4_X1 _23770_ ( .A1(\exu.addi.io_imm [5] ), .A2(_01601_ ), .A3(_01602_ ), .A4(_01604_ ), .ZN(_03075_ ) );
AOI21_X1 _23771_ ( .A(_03075_ ), .B1(_10439_ ), .B2(_01607_ ), .ZN(_03076_ ) );
OAI21_X1 _23772_ ( .A(_03074_ ), .B1(_03076_ ), .B2(\exu.io_in_bits_sub ), .ZN(_03077_ ) );
AOI21_X1 _23773_ ( .A(_03070_ ), .B1(_03077_ ), .B2(_01610_ ), .ZN(_03078_ ) );
OAI221_X1 _23774_ ( .A(_01613_ ), .B1(_08734_ ), .B2(_01832_ ), .C1(_03078_ ), .C2(\exu.io_in_bits_or ), .ZN(_03079_ ) );
OAI21_X1 _23775_ ( .A(_03055_ ), .B1(_01749_ ), .B2(_02021_ ), .ZN(_03080_ ) );
NOR2_X1 _23776_ ( .A1(_03080_ ), .A2(_01579_ ), .ZN(_03081_ ) );
OAI211_X1 _23777_ ( .A(_03079_ ), .B(_01486_ ), .C1(_01614_ ), .C2(_03081_ ), .ZN(_03082_ ) );
NAND3_X1 _23778_ ( .A1(_08733_ ), .A2(_01575_ ), .A3(\exu.and_.io_is ), .ZN(_03083_ ) );
AOI21_X1 _23779_ ( .A(\exu.io_in_bits_xor ), .B1(_03082_ ), .B2(_03083_ ), .ZN(_03084_ ) );
AOI211_X1 _23780_ ( .A(\exu.io_in_bits_sll ), .B(_03084_ ), .C1(_08735_ ), .C2(_01493_ ), .ZN(_03085_ ) );
NAND2_X1 _23781_ ( .A1(_03057_ ), .A2(_01689_ ), .ZN(_03086_ ) );
AOI211_X1 _23782_ ( .A(_01574_ ), .B(_03085_ ), .C1(\exu.io_in_bits_sll ), .C2(_03086_ ), .ZN(_03087_ ) );
XNOR2_X1 _23783_ ( .A(_01366_ ), .B(_08735_ ), .ZN(_03088_ ) );
AOI21_X1 _23784_ ( .A(_03087_ ), .B1(_01828_ ), .B2(_03088_ ), .ZN(_03089_ ) );
OAI221_X1 _23785_ ( .A(_01341_ ), .B1(_01823_ ), .B2(_10441_ ), .C1(_03089_ ), .C2(\exu.io_in_bits_jal ), .ZN(_03090_ ) );
NOR2_X1 _23786_ ( .A1(_10441_ ), .A2(_01855_ ), .ZN(_03091_ ) );
OAI211_X1 _23787_ ( .A(_03090_ ), .B(_01989_ ), .C1(_01854_ ), .C2(_03091_ ), .ZN(_03092_ ) );
MUX2_X1 _23788_ ( .A(_03058_ ), .B(_03092_ ), .S(_01992_ ), .Z(_03093_ ) );
NAND2_X1 _23789_ ( .A1(_03093_ ), .A2(_01994_ ), .ZN(_03094_ ) );
AOI21_X1 _23790_ ( .A(_01797_ ), .B1(_03059_ ), .B2(_03069_ ), .ZN(_03095_ ) );
OAI211_X1 _23791_ ( .A(_03094_ ), .B(_01510_ ), .C1(_01994_ ), .C2(_03095_ ), .ZN(_03096_ ) );
OAI21_X1 _23792_ ( .A(_01186_ ), .B1(\exu.add.io_rs1_data [5] ), .B2(\exu.addi.io_imm [5] ), .ZN(_03097_ ) );
AND2_X1 _23793_ ( .A1(_03097_ ), .A2(_01181_ ), .ZN(_03098_ ) );
AOI221_X4 _23794_ ( .A(fanout_net_5 ), .B1(\exu.io_in_bits_srai ), .B2(_03056_ ), .C1(_03096_ ), .C2(_03098_ ), .ZN(_03099_ ) );
AND3_X1 _23795_ ( .A1(_09067_ ), .A2(_01864_ ), .A3(fanout_net_5 ), .ZN(_03100_ ) );
OAI21_X1 _23796_ ( .A(_01723_ ), .B1(_03099_ ), .B2(_03100_ ), .ZN(_03101_ ) );
NAND2_X1 _23797_ ( .A1(_09069_ ), .A2(_01867_ ), .ZN(_03102_ ) );
AOI21_X1 _23798_ ( .A(_01722_ ), .B1(_03101_ ), .B2(_03102_ ), .ZN(_03103_ ) );
AND2_X1 _23799_ ( .A1(\exu.addi._io_rd_T_4 [5] ), .A2(_01870_ ), .ZN(_03104_ ) );
OAI21_X1 _23800_ ( .A(_01721_ ), .B1(_03103_ ), .B2(_03104_ ), .ZN(_03105_ ) );
OAI211_X1 _23801_ ( .A(_10845_ ), .B(\exu.csrrs.io_csr_rdata [5] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_03106_ ) );
NAND2_X1 _23802_ ( .A1(_03105_ ), .A2(_03106_ ), .ZN(\exu.io_out_bits_rd_wdata [5] ) );
OAI211_X1 _23803_ ( .A(_01568_ ), .B(_01907_ ), .C1(_01912_ ), .C2(_01881_ ), .ZN(_03107_ ) );
NAND2_X1 _23804_ ( .A1(_01885_ ), .A2(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03108_ ) );
NAND3_X1 _23805_ ( .A1(_01901_ ), .A2(_01903_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03109_ ) );
NAND3_X1 _23806_ ( .A1(_03108_ ), .A2(_01888_ ), .A3(_03109_ ), .ZN(_03110_ ) );
OAI211_X1 _23807_ ( .A(_01884_ ), .B(_02989_ ), .C1(_01891_ ), .C2(_01255_ ), .ZN(_03111_ ) );
AND3_X1 _23808_ ( .A1(_03110_ ), .A2(_01734_ ), .A3(_03111_ ), .ZN(_03112_ ) );
AOI21_X1 _23809_ ( .A(_01734_ ), .B1(_02858_ ), .B2(_02860_ ), .ZN(_03113_ ) );
OR3_X1 _23810_ ( .A1(_03112_ ), .A2(_01748_ ), .A3(_03113_ ), .ZN(_03114_ ) );
OAI211_X1 _23811_ ( .A(_03114_ ), .B(_02021_ ), .C1(_01881_ ), .C2(_02552_ ), .ZN(_03115_ ) );
AND3_X1 _23812_ ( .A1(_03107_ ), .A2(_01914_ ), .A3(_03115_ ), .ZN(_03116_ ) );
OAI21_X1 _23813_ ( .A(_01878_ ), .B1(_03116_ ), .B2(_01512_ ), .ZN(_03117_ ) );
OAI21_X1 _23814_ ( .A(_01755_ ), .B1(\exu.add.io_rs1_data [4] ), .B2(\exu.addi.io_imm [4] ), .ZN(_03118_ ) );
NAND3_X1 _23815_ ( .A1(_02872_ ), .A2(_02873_ ), .A3(_01927_ ), .ZN(_03119_ ) );
NAND2_X1 _23816_ ( .A1(_01783_ ), .A2(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03120_ ) );
NAND3_X1 _23817_ ( .A1(_02562_ ), .A2(_02563_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03121_ ) );
NAND3_X1 _23818_ ( .A1(_03120_ ), .A2(_01778_ ), .A3(_03121_ ), .ZN(_03122_ ) );
OAI211_X1 _23819_ ( .A(_01781_ ), .B(_02999_ ), .C1(_01767_ ), .C2(_01255_ ), .ZN(_03123_ ) );
AND2_X1 _23820_ ( .A1(_03122_ ), .A2(_03123_ ), .ZN(_03124_ ) );
INV_X1 _23821_ ( .A(_03124_ ), .ZN(_03125_ ) );
OAI211_X1 _23822_ ( .A(_01206_ ), .B(_03119_ ), .C1(_03125_ ), .C2(_01927_ ), .ZN(_03126_ ) );
OAI21_X1 _23823_ ( .A(_01935_ ), .B1(_02559_ ), .B2(_02566_ ), .ZN(_03127_ ) );
AND3_X1 _23824_ ( .A1(_03126_ ), .A2(_01450_ ), .A3(_03127_ ), .ZN(_03128_ ) );
AOI21_X1 _23825_ ( .A(_03128_ ), .B1(_01942_ ), .B2(_01795_ ), .ZN(_03129_ ) );
NAND2_X1 _23826_ ( .A1(_03129_ ), .A2(_02283_ ), .ZN(_03130_ ) );
NOR3_X1 _23827_ ( .A1(_01949_ ), .A2(_01804_ ), .A3(_01308_ ), .ZN(_03131_ ) );
NAND2_X1 _23828_ ( .A1(_03131_ ), .A2(_01338_ ), .ZN(_03132_ ) );
NOR3_X1 _23829_ ( .A1(_01360_ ), .A2(_08732_ ), .A3(_01362_ ), .ZN(_03133_ ) );
NOR3_X1 _23830_ ( .A1(_01364_ ), .A2(_01694_ ), .A3(_03133_ ), .ZN(_03134_ ) );
NAND2_X1 _23831_ ( .A1(_03131_ ), .A2(_01689_ ), .ZN(_03135_ ) );
NAND2_X1 _23832_ ( .A1(_09203_ ), .A2(_01607_ ), .ZN(_03136_ ) );
NAND4_X1 _23833_ ( .A1(_01601_ ), .A2(\exu.addi.io_imm [4] ), .A3(_01602_ ), .A4(_01604_ ), .ZN(_03137_ ) );
AOI21_X1 _23834_ ( .A(\exu.io_in_bits_sub ), .B1(_03136_ ), .B2(_03137_ ), .ZN(_03138_ ) );
XNOR2_X1 _23835_ ( .A(_08829_ ), .B(_08732_ ), .ZN(_03139_ ) );
AOI21_X1 _23836_ ( .A(_03138_ ), .B1(_01478_ ), .B2(_03139_ ), .ZN(_03140_ ) );
NOR2_X1 _23837_ ( .A1(_03140_ ), .A2(\exu.io_in_bits_srl ), .ZN(_03141_ ) );
AND2_X1 _23838_ ( .A1(_03129_ ), .A2(_01594_ ), .ZN(_03142_ ) );
OAI21_X1 _23839_ ( .A(_02512_ ), .B1(_03141_ ), .B2(_03142_ ), .ZN(_03143_ ) );
OAI21_X1 _23840_ ( .A(_01581_ ), .B1(\exu.add.io_rs1_data [4] ), .B2(\exu._GEN_0 [4] ), .ZN(_03144_ ) );
AOI21_X1 _23841_ ( .A(\exu.io_in_bits_sra ), .B1(_03143_ ), .B2(_03144_ ), .ZN(_03145_ ) );
AND3_X1 _23842_ ( .A1(_03107_ ), .A2(_01445_ ), .A3(_03115_ ), .ZN(_03146_ ) );
OAI21_X1 _23843_ ( .A(_01486_ ), .B1(_03145_ ), .B2(_03146_ ), .ZN(_03147_ ) );
NAND3_X1 _23844_ ( .A1(_01365_ ), .A2(_10699_ ), .A3(\exu.and_.io_is ), .ZN(_03148_ ) );
AOI21_X1 _23845_ ( .A(\exu.io_in_bits_xor ), .B1(_03147_ ), .B2(_03148_ ), .ZN(_03149_ ) );
AOI21_X1 _23846_ ( .A(_03149_ ), .B1(_08732_ ), .B2(_01493_ ), .ZN(_03150_ ) );
OAI21_X1 _23847_ ( .A(_03135_ ), .B1(_03150_ ), .B2(\exu.io_in_bits_sll ), .ZN(_03151_ ) );
AOI21_X1 _23848_ ( .A(_03134_ ), .B1(_03151_ ), .B2(_01498_ ), .ZN(_03152_ ) );
OAI221_X1 _23849_ ( .A(_01341_ ), .B1(_01823_ ), .B2(_09200_ ), .C1(_03152_ ), .C2(\exu.io_in_bits_jal ), .ZN(_03153_ ) );
AND3_X1 _23850_ ( .A1(_09195_ ), .A2(_09198_ ), .A3(_09460_ ), .ZN(_03154_ ) );
OAI211_X1 _23851_ ( .A(_03153_ ), .B(_01989_ ), .C1(_01854_ ), .C2(_03154_ ), .ZN(_03155_ ) );
MUX2_X1 _23852_ ( .A(_03132_ ), .B(_03155_ ), .S(_01992_ ), .Z(_03156_ ) );
MUX2_X1 _23853_ ( .A(_03130_ ), .B(_03156_ ), .S(_01705_ ), .Z(_03157_ ) );
MUX2_X1 _23854_ ( .A(_03118_ ), .B(_03157_ ), .S(_01860_ ), .Z(_03158_ ) );
AOI21_X1 _23855_ ( .A(_03117_ ), .B1(_03158_ ), .B2(_01862_ ), .ZN(_03159_ ) );
AND3_X1 _23856_ ( .A1(_09071_ ), .A2(_01864_ ), .A3(fanout_net_5 ), .ZN(_03160_ ) );
OAI21_X1 _23857_ ( .A(_01723_ ), .B1(_03159_ ), .B2(_03160_ ), .ZN(_03161_ ) );
NAND2_X1 _23858_ ( .A1(_09050_ ), .A2(_01867_ ), .ZN(_03162_ ) );
AOI21_X1 _23859_ ( .A(_01722_ ), .B1(_03161_ ), .B2(_03162_ ), .ZN(_03163_ ) );
AND2_X1 _23860_ ( .A1(\exu.addi._io_rd_T_4 [4] ), .A2(_01870_ ), .ZN(_03164_ ) );
OAI21_X1 _23861_ ( .A(_01721_ ), .B1(_03163_ ), .B2(_03164_ ), .ZN(_03165_ ) );
OAI211_X1 _23862_ ( .A(_10845_ ), .B(\exu.csrrs.io_csr_rdata [4] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_03166_ ) );
NAND2_X1 _23863_ ( .A1(_03165_ ), .A2(_03166_ ), .ZN(\exu.io_out_bits_rd_wdata [4] ) );
NAND2_X1 _23864_ ( .A1(_02020_ ), .A2(_01568_ ), .ZN(_03167_ ) );
OAI211_X1 _23865_ ( .A(_01882_ ), .B(_02920_ ), .C1(_02924_ ), .C2(_01884_ ), .ZN(_03168_ ) );
NAND2_X1 _23866_ ( .A1(_03050_ ), .A2(_01884_ ), .ZN(_03169_ ) );
AND3_X1 _23867_ ( .A1(_01900_ ), .A2(_01902_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03170_ ) );
AOI21_X1 _23868_ ( .A(_01225_ ), .B1(_01900_ ), .B2(_01902_ ), .ZN(_03171_ ) );
OR2_X1 _23869_ ( .A1(_03170_ ), .A2(_03171_ ), .ZN(_03172_ ) );
OAI211_X1 _23870_ ( .A(_03169_ ), .B(_01734_ ), .C1(_01884_ ), .C2(_03172_ ), .ZN(_03173_ ) );
AOI21_X1 _23871_ ( .A(_01748_ ), .B1(_03168_ ), .B2(_03173_ ), .ZN(_03174_ ) );
AOI21_X1 _23872_ ( .A(_01881_ ), .B1(_02661_ ), .B2(_02665_ ), .ZN(_03175_ ) );
OAI21_X1 _23873_ ( .A(_02021_ ), .B1(_03174_ ), .B2(_03175_ ), .ZN(_03176_ ) );
NAND3_X1 _23874_ ( .A1(_03167_ ), .A2(_01914_ ), .A3(_03176_ ), .ZN(_03177_ ) );
NAND3_X1 _23875_ ( .A1(_02043_ ), .A2(_02355_ ), .A3(_01338_ ), .ZN(_03178_ ) );
INV_X1 _23876_ ( .A(_01492_ ), .ZN(_03179_ ) );
AND3_X1 _23877_ ( .A1(_01362_ ), .A2(_01575_ ), .A3(\exu.and_.io_is ), .ZN(_03180_ ) );
NAND3_X1 _23878_ ( .A1(_03167_ ), .A2(_01445_ ), .A3(_03176_ ), .ZN(_03181_ ) );
INV_X1 _23879_ ( .A(\exu.add.io_rs1_data [3] ), .ZN(_03182_ ) );
AOI21_X1 _23880_ ( .A(_01832_ ), .B1(_03182_ ), .B2(_08826_ ), .ZN(_03183_ ) );
NAND2_X1 _23881_ ( .A1(_03064_ ), .A2(_01587_ ), .ZN(_03184_ ) );
AND3_X1 _23882_ ( .A1(_01922_ ), .A2(_01923_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03185_ ) );
AOI21_X1 _23883_ ( .A(_01225_ ), .B1(_02562_ ), .B2(_02563_ ), .ZN(_03186_ ) );
OR2_X1 _23884_ ( .A1(_03185_ ), .A2(_03186_ ), .ZN(_03187_ ) );
OAI211_X1 _23885_ ( .A(_03184_ ), .B(_01788_ ), .C1(_01587_ ), .C2(_03187_ ), .ZN(_03188_ ) );
OAI211_X1 _23886_ ( .A(_01207_ ), .B(_03188_ ), .C1(_02939_ ), .C2(_01788_ ), .ZN(_03189_ ) );
NAND3_X1 _23887_ ( .A1(_02672_ ), .A2(_01935_ ), .A3(_02677_ ), .ZN(_03190_ ) );
AND3_X1 _23888_ ( .A1(_03189_ ), .A2(_03190_ ), .A3(_01212_ ), .ZN(_03191_ ) );
AOI21_X1 _23889_ ( .A(_03191_ ), .B1(_01795_ ), .B2(_02041_ ), .ZN(_03192_ ) );
NAND2_X1 _23890_ ( .A1(_03192_ ), .A2(_01594_ ), .ZN(_03193_ ) );
OR3_X1 _23891_ ( .A1(_08825_ ), .A2(_08820_ ), .A3(_08739_ ), .ZN(_03194_ ) );
OAI21_X1 _23892_ ( .A(_08739_ ), .B1(_08825_ ), .B2(_08820_ ), .ZN(_03195_ ) );
AND3_X1 _23893_ ( .A1(_03194_ ), .A2(_01478_ ), .A3(_03195_ ), .ZN(_03196_ ) );
NAND4_X1 _23894_ ( .A1(_01601_ ), .A2(\exu.addi.io_imm [3] ), .A3(_01602_ ), .A4(_01604_ ), .ZN(_03197_ ) );
OAI21_X1 _23895_ ( .A(_03197_ ), .B1(_11459_ ), .B2(_01460_ ), .ZN(_03198_ ) );
AOI21_X1 _23896_ ( .A(_03196_ ), .B1(_03198_ ), .B2(_01457_ ), .ZN(_03199_ ) );
OAI21_X1 _23897_ ( .A(_03193_ ), .B1(_03199_ ), .B2(\exu.io_in_bits_srl ), .ZN(_03200_ ) );
AOI21_X1 _23898_ ( .A(_03183_ ), .B1(_03200_ ), .B2(_02512_ ), .ZN(_03201_ ) );
OAI21_X1 _23899_ ( .A(_03181_ ), .B1(_03201_ ), .B2(\exu.io_in_bits_sra ), .ZN(_03202_ ) );
AOI21_X1 _23900_ ( .A(_03180_ ), .B1(_03202_ ), .B2(_01486_ ), .ZN(_03203_ ) );
OAI221_X1 _23901_ ( .A(_01438_ ), .B1(_08739_ ), .B2(_03179_ ), .C1(_03203_ ), .C2(\exu.io_in_bits_xor ), .ZN(_03204_ ) );
AND3_X1 _23902_ ( .A1(_02043_ ), .A2(_02354_ ), .A3(_01441_ ), .ZN(_03205_ ) );
OAI211_X1 _23903_ ( .A(_03204_ ), .B(_01498_ ), .C1(_01438_ ), .C2(_03205_ ), .ZN(_03206_ ) );
NAND3_X1 _23904_ ( .A1(_01357_ ), .A2(_01359_ ), .A3(_08739_ ), .ZN(_03207_ ) );
NAND3_X1 _23905_ ( .A1(_01361_ ), .A2(_01828_ ), .A3(_03207_ ), .ZN(_03208_ ) );
AOI21_X1 _23906_ ( .A(\exu.io_in_bits_jal ), .B1(_03206_ ), .B2(_03208_ ), .ZN(_03209_ ) );
AOI21_X1 _23907_ ( .A(_03209_ ), .B1(_09452_ ), .B2(_11443_ ), .ZN(_03210_ ) );
NOR2_X1 _23908_ ( .A1(_03210_ ), .A2(\exu.io_in_bits_jalr ), .ZN(_03211_ ) );
AND2_X1 _23909_ ( .A1(_11443_ ), .A2(_01699_ ), .ZN(_03212_ ) );
OAI21_X1 _23910_ ( .A(_01989_ ), .B1(_03211_ ), .B2(_03212_ ), .ZN(_03213_ ) );
MUX2_X1 _23911_ ( .A(_03178_ ), .B(_03213_ ), .S(_01992_ ), .Z(_03214_ ) );
NAND2_X1 _23912_ ( .A1(_03214_ ), .A2(_01994_ ), .ZN(_03215_ ) );
AOI211_X1 _23913_ ( .A(_01797_ ), .B(_03191_ ), .C1(_01795_ ), .C2(_02041_ ), .ZN(_03216_ ) );
OAI211_X1 _23914_ ( .A(_03215_ ), .B(_01510_ ), .C1(_01994_ ), .C2(_03216_ ), .ZN(_03217_ ) );
AOI21_X1 _23915_ ( .A(\exu.io_in_bits_srai ), .B1(_09066_ ), .B2(_01755_ ), .ZN(_03218_ ) );
AOI221_X4 _23916_ ( .A(fanout_net_5 ), .B1(\exu.io_in_bits_srai ), .B2(_03177_ ), .C1(_03217_ ), .C2(_03218_ ), .ZN(_03219_ ) );
AND3_X1 _23917_ ( .A1(_09061_ ), .A2(_01864_ ), .A3(fanout_net_5 ), .ZN(_03220_ ) );
OAI21_X1 _23918_ ( .A(_01723_ ), .B1(_03219_ ), .B2(_03220_ ), .ZN(_03221_ ) );
NAND3_X1 _23919_ ( .A1(_09062_ ), .A2(_09066_ ), .A3(_01867_ ), .ZN(_03222_ ) );
AOI21_X1 _23920_ ( .A(_01722_ ), .B1(_03221_ ), .B2(_03222_ ), .ZN(_03223_ ) );
NOR2_X1 _23921_ ( .A1(_11473_ ), .A2(_02249_ ), .ZN(_03224_ ) );
OAI21_X1 _23922_ ( .A(_01721_ ), .B1(_03223_ ), .B2(_03224_ ), .ZN(_03225_ ) );
OAI211_X1 _23923_ ( .A(_10845_ ), .B(\exu.csrrs.io_csr_rdata [3] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_03226_ ) );
NAND2_X1 _23924_ ( .A1(_03225_ ), .A2(_03226_ ), .ZN(\exu.io_out_bits_rd_wdata [3] ) );
NAND3_X1 _23925_ ( .A1(_09057_ ), .A2(_10842_ ), .A3(fanout_net_5 ), .ZN(_03227_ ) );
NAND3_X1 _23926_ ( .A1(_03108_ ), .A2(_01884_ ), .A3(_03109_ ), .ZN(_03228_ ) );
AND3_X1 _23927_ ( .A1(_01901_ ), .A2(_01903_ ), .A3(_01225_ ), .ZN(_03229_ ) );
AOI21_X1 _23928_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B1(_01901_ ), .B2(_01903_ ), .ZN(_03230_ ) );
NOR2_X1 _23929_ ( .A1(_03229_ ), .A2(_03230_ ), .ZN(_03231_ ) );
OAI211_X1 _23930_ ( .A(_03228_ ), .B(_01547_ ), .C1(_01884_ ), .C2(_03231_ ), .ZN(_03232_ ) );
NAND3_X1 _23931_ ( .A1(_02988_ ), .A2(_02990_ ), .A3(_01562_ ), .ZN(_03233_ ) );
NAND3_X1 _23932_ ( .A1(_03232_ ), .A2(_03233_ ), .A3(_01541_ ), .ZN(_03234_ ) );
NAND3_X1 _23933_ ( .A1(_02734_ ), .A2(_01747_ ), .A3(_02739_ ), .ZN(_03235_ ) );
AND3_X1 _23934_ ( .A1(_03234_ ), .A2(_01879_ ), .A3(_03235_ ), .ZN(_03236_ ) );
AOI21_X1 _23935_ ( .A(_03236_ ), .B1(_02116_ ), .B2(_01567_ ), .ZN(_03237_ ) );
NAND2_X1 _23936_ ( .A1(_03237_ ), .A2(_01530_ ), .ZN(_03238_ ) );
INV_X1 _23937_ ( .A(_09058_ ), .ZN(_03239_ ) );
NAND2_X1 _23938_ ( .A1(_03239_ ), .A2(_01185_ ), .ZN(_03240_ ) );
NAND3_X1 _23939_ ( .A1(_03120_ ), .A2(_01587_ ), .A3(_03121_ ), .ZN(_03241_ ) );
NAND2_X1 _23940_ ( .A1(_01783_ ), .A2(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03242_ ) );
NAND3_X1 _23941_ ( .A1(_02562_ ), .A2(_02563_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03243_ ) );
NAND2_X1 _23942_ ( .A1(_03242_ ), .A2(_03243_ ), .ZN(_03244_ ) );
OAI211_X1 _23943_ ( .A(_03241_ ), .B(_01590_ ), .C1(_03244_ ), .C2(_01587_ ), .ZN(_03245_ ) );
OAI211_X1 _23944_ ( .A(_03245_ ), .B(_01591_ ), .C1(_01788_ ), .C2(_03001_ ), .ZN(_03246_ ) );
NAND3_X1 _23945_ ( .A1(_02744_ ), .A2(_01790_ ), .A3(_02749_ ), .ZN(_03247_ ) );
AND3_X1 _23946_ ( .A1(_03246_ ), .A2(_01211_ ), .A3(_03247_ ), .ZN(_03248_ ) );
AOI21_X1 _23947_ ( .A(_03248_ ), .B1(_02133_ ), .B2(_01794_ ), .ZN(_03249_ ) );
NAND2_X1 _23948_ ( .A1(_03249_ ), .A2(_01217_ ), .ZN(_03250_ ) );
NAND3_X1 _23949_ ( .A1(_02135_ ), .A2(_02354_ ), .A3(_01336_ ), .ZN(_03251_ ) );
AND2_X1 _23950_ ( .A1(_03249_ ), .A2(_01593_ ), .ZN(_03252_ ) );
OAI21_X1 _23951_ ( .A(_01477_ ), .B1(_08824_ ), .B2(_08779_ ), .ZN(_03253_ ) );
AOI21_X1 _23952_ ( .A(_03253_ ), .B1(_08824_ ), .B2(_08779_ ), .ZN(_03254_ ) );
NAND4_X1 _23953_ ( .A1(_01465_ ), .A2(\exu.addi.io_imm [2] ), .A3(_01462_ ), .A4(_01467_ ), .ZN(_03255_ ) );
OAI21_X1 _23954_ ( .A(_03255_ ), .B1(_11412_ ), .B2(_01460_ ), .ZN(_03256_ ) );
AOI21_X1 _23955_ ( .A(_03254_ ), .B1(_03256_ ), .B2(_01457_ ), .ZN(_03257_ ) );
NOR2_X1 _23956_ ( .A1(_03257_ ), .A2(\exu.io_in_bits_srl ), .ZN(_03258_ ) );
OAI21_X1 _23957_ ( .A(_02512_ ), .B1(_03252_ ), .B2(_03258_ ), .ZN(_03259_ ) );
OAI21_X1 _23958_ ( .A(_01448_ ), .B1(\exu.add.io_rs1_data [2] ), .B2(\exu._GEN_0 [2] ), .ZN(_03260_ ) );
AOI21_X1 _23959_ ( .A(\exu.io_in_bits_sra ), .B1(_03259_ ), .B2(_03260_ ), .ZN(_03261_ ) );
AND2_X1 _23960_ ( .A1(_03237_ ), .A2(_01445_ ), .ZN(_03262_ ) );
OAI21_X1 _23961_ ( .A(_01485_ ), .B1(_03261_ ), .B2(_03262_ ), .ZN(_03263_ ) );
NAND3_X1 _23962_ ( .A1(_01358_ ), .A2(_10698_ ), .A3(\exu.and_.io_is ), .ZN(_03264_ ) );
AOI21_X1 _23963_ ( .A(\exu.io_in_bits_xor ), .B1(_03263_ ), .B2(_03264_ ), .ZN(_03265_ ) );
AND2_X1 _23964_ ( .A1(_08779_ ), .A2(_01492_ ), .ZN(_03266_ ) );
OAI21_X1 _23965_ ( .A(_01438_ ), .B1(_03265_ ), .B2(_03266_ ), .ZN(_03267_ ) );
NAND3_X1 _23966_ ( .A1(_02135_ ), .A2(_01332_ ), .A3(_01440_ ), .ZN(_03268_ ) );
AOI21_X1 _23967_ ( .A(_01572_ ), .B1(_03267_ ), .B2(_03268_ ), .ZN(_03269_ ) );
OR3_X1 _23968_ ( .A1(_01355_ ), .A2(_01356_ ), .A3(_08779_ ), .ZN(_03270_ ) );
AND3_X1 _23969_ ( .A1(_03270_ ), .A2(_01357_ ), .A3(_01435_ ), .ZN(_03271_ ) );
OAI21_X1 _23970_ ( .A(_09410_ ), .B1(_03269_ ), .B2(_03271_ ), .ZN(_03272_ ) );
OAI211_X1 _23971_ ( .A(_03272_ ), .B(_09657_ ), .C1(\exu.auipc.io_rs1_data [2] ), .C2(_09999_ ), .ZN(_03273_ ) );
NOR3_X1 _23972_ ( .A1(_09657_ ), .A2(fanout_net_27 ), .A3(\exu.auipc.io_rs1_data [2] ), .ZN(_03274_ ) );
OAI211_X1 _23973_ ( .A(_03273_ ), .B(_01501_ ), .C1(_09657_ ), .C2(_03274_ ), .ZN(_03275_ ) );
MUX2_X1 _23974_ ( .A(_03251_ ), .B(_03275_ ), .S(_01504_ ), .Z(_03276_ ) );
MUX2_X1 _23975_ ( .A(_03250_ ), .B(_03276_ ), .S(_01214_ ), .Z(_03277_ ) );
MUX2_X1 _23976_ ( .A(_03240_ ), .B(_03277_ ), .S(_02023_ ), .Z(_03278_ ) );
MUX2_X1 _23977_ ( .A(_03238_ ), .B(_03278_ ), .S(_01181_ ), .Z(_03279_ ) );
MUX2_X1 _23978_ ( .A(_03227_ ), .B(_03279_ ), .S(_01176_ ), .Z(_03280_ ) );
OR2_X1 _23979_ ( .A1(_03280_ ), .A2(\exu.io_in_bits_xori ), .ZN(_03281_ ) );
NAND3_X1 _23980_ ( .A1(_09063_ ), .A2(_03239_ ), .A3(_01519_ ), .ZN(_03282_ ) );
AOI21_X1 _23981_ ( .A(_01173_ ), .B1(_03281_ ), .B2(_03282_ ), .ZN(_03283_ ) );
AOI211_X1 _23982_ ( .A(_01718_ ), .B(_03283_ ), .C1(\exu.addi._io_rd_T_4 [2] ), .C2(_02003_ ), .ZN(_03284_ ) );
AOI21_X1 _23983_ ( .A(_01109_ ), .B1(_10845_ ), .B2(\exu.csrrs.io_csr_rdata [2] ), .ZN(_03285_ ) );
NOR2_X1 _23984_ ( .A1(_03284_ ), .A2(_03285_ ), .ZN(\exu.io_out_bits_rd_wdata [2] ) );
OAI21_X1 _23985_ ( .A(_01536_ ), .B1(_02554_ ), .B2(_01568_ ), .ZN(_03286_ ) );
NOR2_X1 _23986_ ( .A1(_03286_ ), .A2(_01752_ ), .ZN(_03287_ ) );
OAI21_X1 _23987_ ( .A(_01515_ ), .B1(_03287_ ), .B2(_01182_ ), .ZN(_03288_ ) );
OAI21_X1 _23988_ ( .A(_01186_ ), .B1(\exu.add.io_rs1_data [28] ), .B2(\exu.addi.io_imm [28] ), .ZN(_03289_ ) );
NAND4_X1 _23989_ ( .A1(_01941_ ), .A2(_01207_ ), .A3(_01213_ ), .A4(_02283_ ), .ZN(_03290_ ) );
OR3_X1 _23990_ ( .A1(_01960_ ), .A2(_01271_ ), .A3(_01963_ ), .ZN(_03291_ ) );
OAI211_X1 _23991_ ( .A(_01253_ ), .B(_01665_ ), .C1(_01297_ ), .C2(_01666_ ), .ZN(_03292_ ) );
OAI211_X1 _23992_ ( .A(_01299_ ), .B(_01673_ ), .C1(_01297_ ), .C2(_01283_ ), .ZN(_03293_ ) );
NAND2_X1 _23993_ ( .A1(_03292_ ), .A2(_03293_ ), .ZN(_03294_ ) );
NAND2_X1 _23994_ ( .A1(_03294_ ), .A2(_01325_ ), .ZN(_03295_ ) );
NOR2_X1 _23995_ ( .A1(_01676_ ), .A2(_01677_ ), .ZN(_03296_ ) );
MUX2_X1 _23996_ ( .A(_03296_ ), .B(_01682_ ), .S(_01299_ ), .Z(_03297_ ) );
OAI211_X1 _23997_ ( .A(_01271_ ), .B(_03295_ ), .C1(_03297_ ), .C2(_01325_ ), .ZN(_03298_ ) );
NAND3_X1 _23998_ ( .A1(_03291_ ), .A2(_02354_ ), .A3(_03298_ ), .ZN(_03299_ ) );
OAI21_X1 _23999_ ( .A(_03299_ ), .B1(_02571_ ), .B2(_02354_ ), .ZN(_03300_ ) );
NAND2_X1 _24000_ ( .A1(_03300_ ), .A2(_01338_ ), .ZN(_03301_ ) );
NAND3_X1 _24001_ ( .A1(_01427_ ), .A2(_10698_ ), .A3(\exu.and_.io_is ), .ZN(_03302_ ) );
NOR2_X1 _24002_ ( .A1(_03286_ ), .A2(_01579_ ), .ZN(_03303_ ) );
OAI21_X1 _24003_ ( .A(_01448_ ), .B1(\exu.add.io_rs1_data [28] ), .B2(\exu._GEN_0 [28] ), .ZN(_03304_ ) );
AND3_X1 _24004_ ( .A1(_02569_ ), .A2(_01450_ ), .A3(_01594_ ), .ZN(_03305_ ) );
NAND2_X1 _24005_ ( .A1(_01472_ ), .A2(_08765_ ), .ZN(_03306_ ) );
NAND3_X1 _24006_ ( .A1(_02634_ ), .A2(_01478_ ), .A3(_03306_ ), .ZN(_03307_ ) );
AND4_X1 _24007_ ( .A1(\exu.addi.io_imm [28] ), .A2(_01600_ ), .A3(_01463_ ), .A4(_01603_ ), .ZN(_03308_ ) );
AOI21_X1 _24008_ ( .A(_03308_ ), .B1(_09353_ ), .B2(_01606_ ), .ZN(_03309_ ) );
OAI21_X1 _24009_ ( .A(_03307_ ), .B1(_03309_ ), .B2(\exu.io_in_bits_sub ), .ZN(_03310_ ) );
AOI21_X1 _24010_ ( .A(_03305_ ), .B1(_03310_ ), .B2(_01481_ ), .ZN(_03311_ ) );
OAI21_X1 _24011_ ( .A(_03304_ ), .B1(_03311_ ), .B2(\exu.io_in_bits_or ), .ZN(_03312_ ) );
AOI21_X1 _24012_ ( .A(_03303_ ), .B1(_03312_ ), .B2(_01613_ ), .ZN(_03313_ ) );
OAI21_X1 _24013_ ( .A(_03302_ ), .B1(_03313_ ), .B2(\exu.and_.io_is ), .ZN(_03314_ ) );
AOI221_X4 _24014_ ( .A(\exu.io_in_bits_sll ), .B1(_08765_ ), .B2(_01968_ ), .C1(_03314_ ), .C2(_01617_ ), .ZN(_03315_ ) );
NAND2_X1 _24015_ ( .A1(_03300_ ), .A2(_01441_ ), .ZN(_03316_ ) );
AOI211_X1 _24016_ ( .A(_01573_ ), .B(_03315_ ), .C1(\exu.io_in_bits_sll ), .C2(_03316_ ), .ZN(_03317_ ) );
AND3_X1 _24017_ ( .A1(_01422_ ), .A2(_01344_ ), .A3(_01425_ ), .ZN(_03318_ ) );
NOR3_X1 _24018_ ( .A1(_03318_ ), .A2(_01426_ ), .A3(_01694_ ), .ZN(_03319_ ) );
OAI21_X1 _24019_ ( .A(_01571_ ), .B1(_03317_ ), .B2(_03319_ ), .ZN(_03320_ ) );
NAND2_X1 _24020_ ( .A1(_09357_ ), .A2(_09452_ ), .ZN(_03321_ ) );
AOI21_X1 _24021_ ( .A(\exu.io_in_bits_jalr ), .B1(_03320_ ), .B2(_03321_ ), .ZN(_03322_ ) );
AND2_X1 _24022_ ( .A1(_09357_ ), .A2(_01699_ ), .ZN(_03323_ ) );
OAI21_X1 _24023_ ( .A(_01501_ ), .B1(_03322_ ), .B2(_03323_ ), .ZN(_03324_ ) );
MUX2_X1 _24024_ ( .A(_03301_ ), .B(_03324_ ), .S(_01505_ ), .Z(_03325_ ) );
MUX2_X1 _24025_ ( .A(_03290_ ), .B(_03325_ ), .S(_01705_ ), .Z(_03326_ ) );
MUX2_X1 _24026_ ( .A(_03289_ ), .B(_03326_ ), .S(_01510_ ), .Z(_03327_ ) );
AOI21_X1 _24027_ ( .A(_03288_ ), .B1(_03327_ ), .B2(_01862_ ), .ZN(_03328_ ) );
AND3_X1 _24028_ ( .A1(_09389_ ), .A2(_10843_ ), .A3(fanout_net_5 ), .ZN(_03329_ ) );
OAI21_X1 _24029_ ( .A(_01175_ ), .B1(_03328_ ), .B2(_03329_ ), .ZN(_03330_ ) );
NAND2_X1 _24030_ ( .A1(_09391_ ), .A2(_01519_ ), .ZN(_03331_ ) );
AOI21_X1 _24031_ ( .A(_01173_ ), .B1(_03330_ ), .B2(_03331_ ), .ZN(_03332_ ) );
NOR3_X1 _24032_ ( .A1(_09393_ ), .A2(_09394_ ), .A3(_02249_ ), .ZN(_03333_ ) );
OAI21_X1 _24033_ ( .A(_01721_ ), .B1(_03332_ ), .B2(_03333_ ), .ZN(_03334_ ) );
OAI211_X1 _24034_ ( .A(_01873_ ), .B(\exu.csrrs.io_csr_rdata [28] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_03335_ ) );
NAND2_X1 _24035_ ( .A1(_03334_ ), .A2(_03335_ ), .ZN(\exu.io_out_bits_rd_wdata [28] ) );
NAND3_X1 _24036_ ( .A1(_09051_ ), .A2(_10842_ ), .A3(\exu.andi.io_is ), .ZN(_03336_ ) );
NAND2_X1 _24037_ ( .A1(_02191_ ), .A2(_01566_ ), .ZN(_03337_ ) );
NAND3_X1 _24038_ ( .A1(_02257_ ), .A2(_02258_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03338_ ) );
OAI211_X1 _24039_ ( .A(_01887_ ), .B(_03338_ ), .C1(_01890_ ), .C2(_01629_ ), .ZN(_03339_ ) );
OAI211_X1 _24040_ ( .A(_01546_ ), .B(_03339_ ), .C1(_03172_ ), .C2(_01888_ ), .ZN(_03340_ ) );
OAI211_X1 _24041_ ( .A(_03340_ ), .B(_01541_ ), .C1(_03053_ ), .C2(_01547_ ), .ZN(_03341_ ) );
OAI211_X1 _24042_ ( .A(_03341_ ), .B(_01533_ ), .C1(_02800_ ), .C2(_01541_ ), .ZN(_03342_ ) );
NAND3_X1 _24043_ ( .A1(_03337_ ), .A2(_01914_ ), .A3(_03342_ ), .ZN(_03343_ ) );
NAND2_X1 _24044_ ( .A1(_11355_ ), .A2(_01185_ ), .ZN(_03344_ ) );
NAND3_X1 _24045_ ( .A1(_02562_ ), .A2(_02563_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03345_ ) );
OAI211_X1 _24046_ ( .A(_01763_ ), .B(_03345_ ), .C1(_01767_ ), .C2(_01629_ ), .ZN(_03346_ ) );
OAI211_X1 _24047_ ( .A(_01590_ ), .B(_03346_ ), .C1(_03187_ ), .C2(_01778_ ), .ZN(_03347_ ) );
NAND3_X1 _24048_ ( .A1(_03065_ ), .A2(_01771_ ), .A3(_03066_ ), .ZN(_03348_ ) );
NAND3_X1 _24049_ ( .A1(_03347_ ), .A2(_03348_ ), .A3(_01591_ ), .ZN(_03349_ ) );
OAI211_X1 _24050_ ( .A(_01211_ ), .B(_03349_ ), .C1(_02816_ ), .C2(_01591_ ), .ZN(_03350_ ) );
NAND3_X1 _24051_ ( .A1(_02199_ ), .A2(_01793_ ), .A3(_02206_ ), .ZN(_03351_ ) );
NAND3_X1 _24052_ ( .A1(_03350_ ), .A2(_01217_ ), .A3(_03351_ ), .ZN(_03352_ ) );
AND2_X1 _24053_ ( .A1(_02220_ ), .A2(_01271_ ), .ZN(_03353_ ) );
NAND3_X1 _24054_ ( .A1(_03353_ ), .A2(_02355_ ), .A3(_01337_ ), .ZN(_03354_ ) );
NAND3_X1 _24055_ ( .A1(_01356_ ), .A2(_09463_ ), .A3(\exu.and_.io_is ), .ZN(_03355_ ) );
AND3_X1 _24056_ ( .A1(_03337_ ), .A2(_01444_ ), .A3(_03342_ ), .ZN(_03356_ ) );
OAI21_X1 _24057_ ( .A(_01447_ ), .B1(\exu.add.io_rs1_data [1] ), .B2(\exu._GEN_0 [1] ), .ZN(_03357_ ) );
AND3_X1 _24058_ ( .A1(_03350_ ), .A2(_01593_ ), .A3(_03351_ ), .ZN(_03358_ ) );
AND3_X1 _24059_ ( .A1(_08778_ ), .A2(_08821_ ), .A3(\exu._GEN_0 [0] ), .ZN(_03359_ ) );
OR3_X1 _24060_ ( .A1(_03359_ ), .A2(_08822_ ), .A3(_01596_ ), .ZN(_03360_ ) );
AND4_X1 _24061_ ( .A1(\exu.addi.io_imm [1] ), .A2(_01465_ ), .A3(_01462_ ), .A4(_01467_ ), .ZN(_03361_ ) );
AOI21_X1 _24062_ ( .A(_03361_ ), .B1(_11330_ ), .B2(_01606_ ), .ZN(_03362_ ) );
OAI21_X1 _24063_ ( .A(_03360_ ), .B1(_03362_ ), .B2(\exu.io_in_bits_sub ), .ZN(_03363_ ) );
AOI21_X1 _24064_ ( .A(_03358_ ), .B1(_01452_ ), .B2(_03363_ ), .ZN(_03364_ ) );
OAI21_X1 _24065_ ( .A(_03357_ ), .B1(_03364_ ), .B2(\exu.io_in_bits_or ), .ZN(_03365_ ) );
AOI21_X1 _24066_ ( .A(_03356_ ), .B1(_03365_ ), .B2(_01443_ ), .ZN(_03366_ ) );
OAI21_X1 _24067_ ( .A(_03355_ ), .B1(_03366_ ), .B2(\exu.and_.io_is ), .ZN(_03367_ ) );
AOI221_X4 _24068_ ( .A(\exu.io_in_bits_sll ), .B1(_08778_ ), .B2(_01491_ ), .C1(_03367_ ), .C2(_01617_ ), .ZN(_03368_ ) );
NAND3_X1 _24069_ ( .A1(_03353_ ), .A2(_01332_ ), .A3(_01440_ ), .ZN(_03369_ ) );
AOI211_X1 _24070_ ( .A(_01572_ ), .B(_03368_ ), .C1(\exu.io_in_bits_sll ), .C2(_03369_ ), .ZN(_03370_ ) );
NOR2_X1 _24071_ ( .A1(_08778_ ), .A2(_01354_ ), .ZN(_03371_ ) );
NOR3_X1 _24072_ ( .A1(_01355_ ), .A2(_03371_ ), .A3(_01693_ ), .ZN(_03372_ ) );
NOR2_X1 _24073_ ( .A1(_03370_ ), .A2(_03372_ ), .ZN(_03373_ ) );
OAI221_X1 _24074_ ( .A(_09657_ ), .B1(\exu.addi._io_rd_T_4_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_B ), .B2(_09999_ ), .C1(_03373_ ), .C2(\exu.io_in_bits_jal ), .ZN(_03374_ ) );
NOR3_X1 _24075_ ( .A1(_09657_ ), .A2(fanout_net_27 ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_B ), .ZN(_03375_ ) );
OAI211_X1 _24076_ ( .A(_03374_ ), .B(_01501_ ), .C1(_01340_ ), .C2(_03375_ ), .ZN(_03376_ ) );
MUX2_X1 _24077_ ( .A(_03354_ ), .B(_03376_ ), .S(_01504_ ), .Z(_03377_ ) );
MUX2_X1 _24078_ ( .A(_03352_ ), .B(_03377_ ), .S(_01214_ ), .Z(_03378_ ) );
MUX2_X1 _24079_ ( .A(_03344_ ), .B(_03378_ ), .S(_02023_ ), .Z(_03379_ ) );
MUX2_X1 _24080_ ( .A(_03343_ ), .B(_03379_ ), .S(_01181_ ), .Z(_03380_ ) );
MUX2_X1 _24081_ ( .A(_03336_ ), .B(_03380_ ), .S(_01176_ ), .Z(_03381_ ) );
OR2_X1 _24082_ ( .A1(_03381_ ), .A2(\exu.io_in_bits_xori ), .ZN(_03382_ ) );
NAND3_X1 _24083_ ( .A1(_09052_ ), .A2(_11355_ ), .A3(_01867_ ), .ZN(_03383_ ) );
AOI21_X1 _24084_ ( .A(_01722_ ), .B1(_03382_ ), .B2(_03383_ ), .ZN(_03384_ ) );
AOI211_X1 _24085_ ( .A(_01718_ ), .B(_03384_ ), .C1(_11358_ ), .C2(_02003_ ), .ZN(_03385_ ) );
AOI21_X1 _24086_ ( .A(_01721_ ), .B1(_01058_ ), .B2(\exu.csrrs.io_csr_rdata [1] ), .ZN(_03386_ ) );
NOR2_X1 _24087_ ( .A1(_03385_ ), .A2(_03386_ ), .ZN(\exu.io_out_bits_rd_wdata [1] ) );
OAI21_X1 _24088_ ( .A(_01747_ ), .B1(_02861_ ), .B2(_02862_ ), .ZN(_03387_ ) );
NAND3_X1 _24089_ ( .A1(_03110_ ), .A2(_01882_ ), .A3(_03111_ ), .ZN(_03388_ ) );
NAND3_X1 _24090_ ( .A1(_01901_ ), .A2(_01903_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03389_ ) );
INV_X1 _24091_ ( .A(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03390_ ) );
OAI211_X1 _24092_ ( .A(_01888_ ), .B(_03389_ ), .C1(_01891_ ), .C2(_03390_ ), .ZN(_03391_ ) );
OAI211_X1 _24093_ ( .A(_03391_ ), .B(_01547_ ), .C1(_03231_ ), .C2(_01888_ ), .ZN(_03392_ ) );
NAND3_X1 _24094_ ( .A1(_03388_ ), .A2(_01541_ ), .A3(_03392_ ), .ZN(_03393_ ) );
AOI21_X1 _24095_ ( .A(_01567_ ), .B1(_03387_ ), .B2(_03393_ ), .ZN(_03394_ ) );
AOI21_X1 _24096_ ( .A(_03394_ ), .B1(_02267_ ), .B2(_01567_ ), .ZN(_03395_ ) );
OR2_X1 _24097_ ( .A1(_03395_ ), .A2(_01578_ ), .ZN(_03396_ ) );
AOI21_X1 _24098_ ( .A(_01832_ ), .B1(_08821_ ), .B2(_01089_ ), .ZN(_03397_ ) );
NAND3_X1 _24099_ ( .A1(_02562_ ), .A2(_02563_ ), .A3(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03398_ ) );
OAI211_X1 _24100_ ( .A(_01778_ ), .B(_03398_ ), .C1(_01767_ ), .C2(_03390_ ), .ZN(_03399_ ) );
OAI211_X1 _24101_ ( .A(_01590_ ), .B(_03399_ ), .C1(_03244_ ), .C2(_01778_ ), .ZN(_03400_ ) );
OAI211_X1 _24102_ ( .A(_01591_ ), .B(_03400_ ), .C1(_03125_ ), .C2(_01788_ ), .ZN(_03401_ ) );
OAI21_X1 _24103_ ( .A(_03401_ ), .B1(_02875_ ), .B2(_01205_ ), .ZN(_03402_ ) );
MUX2_X1 _24104_ ( .A(_03402_ ), .B(_02282_ ), .S(_01794_ ), .Z(_03403_ ) );
NAND2_X1 _24105_ ( .A1(_03403_ ), .A2(_01593_ ), .ZN(_03404_ ) );
NAND2_X1 _24106_ ( .A1(_11366_ ), .A2(_01606_ ), .ZN(_03405_ ) );
NAND4_X1 _24107_ ( .A1(_01465_ ), .A2(\exu.addi.io_imm [0] ), .A3(_01462_ ), .A4(_01467_ ), .ZN(_03406_ ) );
AOI21_X1 _24108_ ( .A(\exu.io_in_bits_sub ), .B1(_03405_ ), .B2(_03406_ ), .ZN(_03407_ ) );
AOI21_X1 _24109_ ( .A(_03407_ ), .B1(_08740_ ), .B2(_01478_ ), .ZN(_03408_ ) );
OAI21_X1 _24110_ ( .A(_03404_ ), .B1(\exu.io_in_bits_srl ), .B2(_03408_ ), .ZN(_03409_ ) );
AOI21_X1 _24111_ ( .A(_03397_ ), .B1(_03409_ ), .B2(_02512_ ), .ZN(_03410_ ) );
OAI211_X1 _24112_ ( .A(_01485_ ), .B(_03396_ ), .C1(_03410_ ), .C2(\exu.io_in_bits_sra ), .ZN(_03411_ ) );
AND3_X1 _24113_ ( .A1(_01354_ ), .A2(_09463_ ), .A3(\exu.and_.io_is ), .ZN(_03412_ ) );
OAI211_X1 _24114_ ( .A(_03411_ ), .B(_01617_ ), .C1(_01486_ ), .C2(_03412_ ), .ZN(_03413_ ) );
OAI211_X1 _24115_ ( .A(_03413_ ), .B(_01438_ ), .C1(_08741_ ), .C2(_03179_ ), .ZN(_03414_ ) );
AND3_X1 _24116_ ( .A1(_01944_ ), .A2(_01270_ ), .A3(_01279_ ), .ZN(_03415_ ) );
AND3_X1 _24117_ ( .A1(_03415_ ), .A2(_01332_ ), .A3(_01439_ ), .ZN(_03416_ ) );
OAI21_X1 _24118_ ( .A(_03414_ ), .B1(_01438_ ), .B2(_03416_ ), .ZN(_03417_ ) );
MUX2_X1 _24119_ ( .A(_09798_ ), .B(_03417_ ), .S(_01497_ ), .Z(_03418_ ) );
MUX2_X1 _24120_ ( .A(_03418_ ), .B(_09535_ ), .S(\exu.io_in_bits_sltu ), .Z(_03419_ ) );
NAND2_X1 _24121_ ( .A1(_08740_ ), .A2(_01828_ ), .ZN(_03420_ ) );
MUX2_X1 _24122_ ( .A(_03419_ ), .B(_03420_ ), .S(\exu.add.io_is ), .Z(_03421_ ) );
OAI221_X1 _24123_ ( .A(_01854_ ), .B1(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .B2(_01823_ ), .C1(_03421_ ), .C2(\exu.io_in_bits_jal ), .ZN(_03422_ ) );
NOR3_X1 _24124_ ( .A1(_01854_ ), .A2(fanout_net_27 ), .A3(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03423_ ) );
OAI211_X1 _24125_ ( .A(_03422_ ), .B(_01570_ ), .C1(_01854_ ), .C2(_03423_ ), .ZN(_03424_ ) );
NAND3_X1 _24126_ ( .A1(_03415_ ), .A2(_02355_ ), .A3(_01702_ ), .ZN(_03425_ ) );
AOI21_X1 _24127_ ( .A(\exu.io_in_bits_srli ), .B1(_03424_ ), .B2(_03425_ ), .ZN(_03426_ ) );
AND2_X1 _24128_ ( .A1(_03403_ ), .A2(_02283_ ), .ZN(_03427_ ) );
OAI21_X1 _24129_ ( .A(_01510_ ), .B1(_03426_ ), .B2(_03427_ ), .ZN(_03428_ ) );
OAI211_X1 _24130_ ( .A(_10699_ ), .B(\exu.io_in_bits_ori ), .C1(\exu.addi.io_imm [0] ), .C2(\exu.add.io_rs1_data [0] ), .ZN(_03429_ ) );
AOI21_X1 _24131_ ( .A(\exu.io_in_bits_srai ), .B1(_03428_ ), .B2(_03429_ ), .ZN(_03430_ ) );
NOR2_X1 _24132_ ( .A1(_03395_ ), .A2(_01751_ ), .ZN(_03431_ ) );
OAI21_X1 _24133_ ( .A(_01176_ ), .B1(_03430_ ), .B2(_03431_ ), .ZN(_03432_ ) );
NAND4_X1 _24134_ ( .A1(_10842_ ), .A2(\exu.addi.io_imm [0] ), .A3(\exu.add.io_rs1_data [0] ), .A4(\exu.andi.io_is ), .ZN(_03433_ ) );
AOI21_X1 _24135_ ( .A(\exu.io_in_bits_xori ), .B1(_03432_ ), .B2(_03433_ ), .ZN(_03434_ ) );
AND3_X1 _24136_ ( .A1(_09054_ ), .A2(_12829_ ), .A3(_01518_ ), .ZN(_03435_ ) );
OAI21_X1 _24137_ ( .A(_01169_ ), .B1(_03434_ ), .B2(_03435_ ), .ZN(_03436_ ) );
NOR2_X1 _24138_ ( .A1(_09766_ ), .A2(_09709_ ), .ZN(_03437_ ) );
AND3_X1 _24139_ ( .A1(_03437_ ), .A2(_09392_ ), .A3(_09702_ ), .ZN(_03438_ ) );
NOR4_X1 _24140_ ( .A1(_09387_ ), .A2(_09172_ ), .A3(_09163_ ), .A4(_09166_ ), .ZN(_03439_ ) );
AND2_X1 _24141_ ( .A1(_03438_ ), .A2(_03439_ ), .ZN(_03440_ ) );
INV_X1 _24142_ ( .A(_03440_ ), .ZN(_03441_ ) );
OAI211_X1 _24143_ ( .A(_09154_ ), .B(_09155_ ), .C1(_09148_ ), .C2(_09149_ ), .ZN(_03442_ ) );
NOR2_X1 _24144_ ( .A1(_03442_ ), .A2(_09147_ ), .ZN(_03443_ ) );
NOR2_X1 _24145_ ( .A1(_09045_ ), .A2(_09048_ ), .ZN(_03444_ ) );
NAND2_X1 _24146_ ( .A1(_03443_ ), .A2(_03444_ ), .ZN(_03445_ ) );
NOR3_X1 _24147_ ( .A1(_03445_ ), .A2(_09126_ ), .A3(_09129_ ), .ZN(_03446_ ) );
INV_X1 _24148_ ( .A(_03446_ ), .ZN(_03447_ ) );
NOR2_X1 _24149_ ( .A1(_09105_ ), .A2(_09108_ ), .ZN(_03448_ ) );
INV_X1 _24150_ ( .A(_03448_ ), .ZN(_03449_ ) );
NOR3_X1 _24151_ ( .A1(_03449_ ), .A2(_09111_ ), .A3(_09114_ ), .ZN(_03450_ ) );
NOR2_X1 _24152_ ( .A1(_09089_ ), .A2(_09092_ ), .ZN(_03451_ ) );
INV_X1 _24153_ ( .A(_03451_ ), .ZN(_03452_ ) );
OR3_X1 _24154_ ( .A1(_03452_ ), .A2(_09082_ ), .A3(_09085_ ), .ZN(_03453_ ) );
NOR3_X1 _24155_ ( .A1(_10514_ ), .A2(_08831_ ), .A3(\exu.addi.io_imm [6] ), .ZN(_03454_ ) );
OR3_X1 _24156_ ( .A1(_09069_ ), .A2(_08834_ ), .A3(\exu.addi.io_imm [4] ), .ZN(_03455_ ) );
NAND2_X1 _24157_ ( .A1(_08607_ ), .A2(\exu.add.io_rs1_data [5] ), .ZN(_03456_ ) );
AOI211_X1 _24158_ ( .A(_10425_ ), .B(_10514_ ), .C1(_03455_ ), .C2(_03456_ ), .ZN(_03457_ ) );
INV_X1 _24159_ ( .A(\exu.addi.io_imm [7] ), .ZN(_03458_ ) );
AOI211_X1 _24160_ ( .A(_03454_ ), .B(_03457_ ), .C1(\exu.add.io_rs1_data [7] ), .C2(_03458_ ), .ZN(_03459_ ) );
NOR4_X1 _24161_ ( .A1(_10425_ ), .A2(_09050_ ), .A3(_09069_ ), .A4(_10514_ ), .ZN(_03460_ ) );
OR3_X1 _24162_ ( .A1(_11471_ ), .A2(_08819_ ), .A3(\exu.addi.io_imm [2] ), .ZN(_03461_ ) );
OAI21_X1 _24163_ ( .A(_03461_ ), .B1(_03182_ ), .B2(\exu.addi.io_imm [3] ), .ZN(_03462_ ) );
NAND2_X1 _24164_ ( .A1(_08590_ ), .A2(\exu.add.io_rs1_data [1] ), .ZN(_03463_ ) );
NAND2_X1 _24165_ ( .A1(_08821_ ), .A2(\exu.addi.io_imm [0] ), .ZN(_03464_ ) );
OAI21_X1 _24166_ ( .A(_03464_ ), .B1(_09051_ ), .B2(_09055_ ), .ZN(_03465_ ) );
AOI211_X1 _24167_ ( .A(_09059_ ), .B(_11471_ ), .C1(_03463_ ), .C2(_03465_ ), .ZN(_03466_ ) );
OAI21_X1 _24168_ ( .A(_03460_ ), .B1(_03462_ ), .B2(_03466_ ), .ZN(_03467_ ) );
AOI21_X1 _24169_ ( .A(_03453_ ), .B1(_03459_ ), .B2(_03467_ ), .ZN(_03468_ ) );
NOR3_X1 _24170_ ( .A1(_09085_ ), .A2(_08841_ ), .A3(\exu.addi.io_imm [8] ), .ZN(_03469_ ) );
INV_X1 _24171_ ( .A(\exu.add.io_rs1_data [9] ), .ZN(_03470_ ) );
NOR2_X1 _24172_ ( .A1(_03470_ ), .A2(\exu.addi.io_imm [9] ), .ZN(_03471_ ) );
OAI21_X1 _24173_ ( .A(_03451_ ), .B1(_03469_ ), .B2(_03471_ ), .ZN(_03472_ ) );
OR2_X1 _24174_ ( .A1(_08848_ ), .A2(\exu.addi.io_imm [11] ), .ZN(_03473_ ) );
OR3_X1 _24175_ ( .A1(_09092_ ), .A2(_08850_ ), .A3(\exu.addi.io_imm [10] ), .ZN(_03474_ ) );
NAND3_X1 _24176_ ( .A1(_03472_ ), .A2(_03473_ ), .A3(_03474_ ), .ZN(_03475_ ) );
OAI21_X1 _24177_ ( .A(_03450_ ), .B1(_03468_ ), .B2(_03475_ ), .ZN(_03476_ ) );
NOR2_X1 _24178_ ( .A1(_08855_ ), .A2(\exu.addi.io_imm [12] ), .ZN(_03477_ ) );
OAI21_X1 _24179_ ( .A(_03477_ ), .B1(_09109_ ), .B2(_09110_ ), .ZN(_03478_ ) );
NAND2_X1 _24180_ ( .A1(_08649_ ), .A2(\exu.add.io_rs1_data [13] ), .ZN(_03479_ ) );
AOI21_X1 _24181_ ( .A(_03449_ ), .B1(_03478_ ), .B2(_03479_ ), .ZN(_03480_ ) );
NOR2_X1 _24182_ ( .A1(_08862_ ), .A2(\exu.addi.io_imm [15] ), .ZN(_03481_ ) );
NOR3_X1 _24183_ ( .A1(_09105_ ), .A2(_08860_ ), .A3(\exu.addi.io_imm [14] ), .ZN(_03482_ ) );
NOR3_X1 _24184_ ( .A1(_03480_ ), .A2(_03481_ ), .A3(_03482_ ), .ZN(_03483_ ) );
AOI21_X1 _24185_ ( .A(_03447_ ), .B1(_03476_ ), .B2(_03483_ ), .ZN(_03484_ ) );
INV_X1 _24186_ ( .A(_03484_ ), .ZN(_03485_ ) );
NAND3_X1 _24187_ ( .A1(_09154_ ), .A2(\exu.add.io_rs1_data [22] ), .A3(_09157_ ), .ZN(_03486_ ) );
NOR3_X1 _24188_ ( .A1(_09147_ ), .A2(_08891_ ), .A3(\exu.addi.io_imm [20] ), .ZN(_03487_ ) );
INV_X1 _24189_ ( .A(\exu.addi.io_imm [21] ), .ZN(_03488_ ) );
AOI21_X1 _24190_ ( .A(_03487_ ), .B1(\exu.add.io_rs1_data [21] ), .B2(_03488_ ), .ZN(_03489_ ) );
NOR3_X1 _24191_ ( .A1(_03489_ ), .A2(_09141_ ), .A3(_09144_ ), .ZN(_03490_ ) );
AOI21_X1 _24192_ ( .A(_03490_ ), .B1(\exu.add.io_rs1_data [23] ), .B2(_08667_ ), .ZN(_03491_ ) );
AND3_X1 _24193_ ( .A1(_03485_ ), .A2(_03486_ ), .A3(_03491_ ), .ZN(_03492_ ) );
NOR3_X1 _24194_ ( .A1(_09129_ ), .A2(_08877_ ), .A3(\exu.addi.io_imm [16] ), .ZN(_03493_ ) );
INV_X1 _24195_ ( .A(\exu.add.io_rs1_data [17] ), .ZN(_03494_ ) );
NOR2_X1 _24196_ ( .A1(_03494_ ), .A2(\exu.addi.io_imm [17] ), .ZN(_03495_ ) );
OAI21_X1 _24197_ ( .A(_03444_ ), .B1(_03493_ ), .B2(_03495_ ), .ZN(_03496_ ) );
OR3_X1 _24198_ ( .A1(_09045_ ), .A2(_08884_ ), .A3(\exu.addi.io_imm [18] ), .ZN(_03497_ ) );
NAND2_X1 _24199_ ( .A1(_03496_ ), .A2(_03497_ ), .ZN(_03498_ ) );
NOR2_X1 _24200_ ( .A1(_08882_ ), .A2(\exu.addi.io_imm [19] ), .ZN(_03499_ ) );
OAI21_X1 _24201_ ( .A(_03443_ ), .B1(_03498_ ), .B2(_03499_ ), .ZN(_03500_ ) );
AOI21_X1 _24202_ ( .A(_03441_ ), .B1(_03492_ ), .B2(_03500_ ), .ZN(_03501_ ) );
INV_X1 _24203_ ( .A(_03501_ ), .ZN(_03502_ ) );
OAI211_X1 _24204_ ( .A(\exu.add.io_rs1_data [28] ), .B(_09704_ ), .C1(_09699_ ), .C2(_09700_ ), .ZN(_03503_ ) );
OAI21_X1 _24205_ ( .A(_03503_ ), .B1(_08869_ ), .B2(\exu.addi.io_imm [29] ), .ZN(_03504_ ) );
AND2_X1 _24206_ ( .A1(_03504_ ), .A2(_03437_ ), .ZN(_03505_ ) );
INV_X1 _24207_ ( .A(\exu.add.io_rs1_data [30] ), .ZN(_03506_ ) );
NOR3_X1 _24208_ ( .A1(_09766_ ), .A2(_03506_ ), .A3(\exu.addi.io_imm [30] ), .ZN(_03507_ ) );
NOR2_X1 _24209_ ( .A1(_08875_ ), .A2(\exu.addi.io_imm [31] ), .ZN(_03508_ ) );
OR3_X1 _24210_ ( .A1(_03505_ ), .A2(_03507_ ), .A3(_03508_ ), .ZN(_03509_ ) );
NOR3_X1 _24211_ ( .A1(_09387_ ), .A2(_08911_ ), .A3(\exu.addi.io_imm [26] ), .ZN(_03510_ ) );
OR3_X1 _24212_ ( .A1(_09166_ ), .A2(_08903_ ), .A3(\exu.addi.io_imm [24] ), .ZN(_03511_ ) );
OAI21_X1 _24213_ ( .A(_03511_ ), .B1(_08908_ ), .B2(\exu.addi.io_imm [25] ), .ZN(_03512_ ) );
NOR2_X1 _24214_ ( .A1(_09387_ ), .A2(_09172_ ), .ZN(_03513_ ) );
AOI21_X1 _24215_ ( .A(_03510_ ), .B1(_03512_ ), .B2(_03513_ ), .ZN(_03514_ ) );
OAI21_X1 _24216_ ( .A(_03514_ ), .B1(_08913_ ), .B2(\exu.addi.io_imm [27] ), .ZN(_03515_ ) );
AOI21_X1 _24217_ ( .A(_03509_ ), .B1(_03515_ ), .B2(_03438_ ), .ZN(_03516_ ) );
AND2_X1 _24218_ ( .A1(_03502_ ), .A2(_03516_ ), .ZN(_03517_ ) );
NAND3_X1 _24219_ ( .A1(_03517_ ), .A2(_10844_ ), .A3(\exu.io_in_bits_sltiu ), .ZN(_03518_ ) );
AOI21_X1 _24220_ ( .A(\exu.io_in_bits_slti ), .B1(_03436_ ), .B2(_03518_ ), .ZN(_03519_ ) );
OAI21_X1 _24221_ ( .A(\exu.io_in_bits_slti ), .B1(_03517_ ), .B2(_09766_ ), .ZN(_03520_ ) );
AOI211_X1 _24222_ ( .A(fanout_net_27 ), .B(_03520_ ), .C1(_09766_ ), .C2(_03517_ ), .ZN(_03521_ ) );
OAI21_X1 _24223_ ( .A(_01522_ ), .B1(_03519_ ), .B2(_03521_ ), .ZN(_03522_ ) );
OAI21_X1 _24224_ ( .A(_03522_ ), .B1(_12827_ ), .B2(_02249_ ), .ZN(_03523_ ) );
NAND2_X1 _24225_ ( .A1(_03523_ ), .A2(_01875_ ), .ZN(_03524_ ) );
OAI211_X1 _24226_ ( .A(_10845_ ), .B(\exu.csrrs.io_csr_rdata [0] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_03525_ ) );
NAND2_X1 _24227_ ( .A1(_03524_ ), .A2(_03525_ ), .ZN(\exu.io_out_bits_rd_wdata [0] ) );
OAI21_X1 _24228_ ( .A(_01536_ ), .B1(_02668_ ), .B2(_01567_ ), .ZN(_03526_ ) );
NOR2_X1 _24229_ ( .A1(_03526_ ), .A2(_01752_ ), .ZN(_03527_ ) );
OAI21_X1 _24230_ ( .A(_01515_ ), .B1(_03527_ ), .B2(_01182_ ), .ZN(_03528_ ) );
OAI21_X1 _24231_ ( .A(_01186_ ), .B1(\exu.add.io_rs1_data [27] ), .B2(\exu.addi.io_imm [27] ), .ZN(_03529_ ) );
NAND4_X1 _24232_ ( .A1(_02040_ ), .A2(_01207_ ), .A3(_01213_ ), .A4(_02283_ ), .ZN(_03530_ ) );
NAND2_X1 _24233_ ( .A1(_02684_ ), .A2(_01804_ ), .ZN(_03531_ ) );
OR3_X1 _24234_ ( .A1(_01314_ ), .A2(_01316_ ), .A3(_01254_ ), .ZN(_03532_ ) );
AND3_X1 _24235_ ( .A1(_03532_ ), .A2(_01325_ ), .A3(_01313_ ), .ZN(_03533_ ) );
AOI21_X1 _24236_ ( .A(_01325_ ), .B1(_01289_ ), .B2(_01295_ ), .ZN(_03534_ ) );
OAI21_X1 _24237_ ( .A(_01686_ ), .B1(_03533_ ), .B2(_03534_ ), .ZN(_03535_ ) );
OAI211_X1 _24238_ ( .A(_03535_ ), .B(_02354_ ), .C1(_02046_ ), .C2(_01686_ ), .ZN(_03536_ ) );
NAND2_X1 _24239_ ( .A1(_03531_ ), .A2(_03536_ ), .ZN(_03537_ ) );
NAND2_X1 _24240_ ( .A1(_03537_ ), .A2(_01338_ ), .ZN(_03538_ ) );
NAND3_X1 _24241_ ( .A1(_01423_ ), .A2(_10698_ ), .A3(\exu.and_.io_is ), .ZN(_03539_ ) );
NOR2_X1 _24242_ ( .A1(_03526_ ), .A2(_01579_ ), .ZN(_03540_ ) );
OAI21_X1 _24243_ ( .A(_01448_ ), .B1(\exu.add.io_rs1_data [27] ), .B2(\exu._GEN_0 [27] ), .ZN(_03541_ ) );
NAND3_X1 _24244_ ( .A1(_02040_ ), .A2(_01207_ ), .A3(_01450_ ), .ZN(_03542_ ) );
NOR2_X1 _24245_ ( .A1(_03542_ ), .A2(_01455_ ), .ZN(_03543_ ) );
AOI21_X1 _24246_ ( .A(_01460_ ), .B1(_09424_ ), .B2(_09425_ ), .ZN(_03544_ ) );
AND4_X1 _24247_ ( .A1(\exu.addi.io_imm [27] ), .A2(_01600_ ), .A3(_01463_ ), .A4(_01603_ ), .ZN(_03545_ ) );
OAI21_X1 _24248_ ( .A(_01457_ ), .B1(_03544_ ), .B2(_03545_ ), .ZN(_03546_ ) );
AOI21_X1 _24249_ ( .A(_08909_ ), .B1(_01471_ ), .B2(_08770_ ), .ZN(_03547_ ) );
NOR2_X1 _24250_ ( .A1(_03547_ ), .A2(_08772_ ), .ZN(_03548_ ) );
INV_X1 _24251_ ( .A(_03548_ ), .ZN(_03549_ ) );
OAI21_X1 _24252_ ( .A(_03549_ ), .B1(_08911_ ), .B2(\exu._GEN_0 [26] ), .ZN(_03550_ ) );
INV_X1 _24253_ ( .A(_08771_ ), .ZN(_03551_ ) );
XNOR2_X1 _24254_ ( .A(_03550_ ), .B(_03551_ ), .ZN(_03552_ ) );
OAI21_X1 _24255_ ( .A(_03546_ ), .B1(_01597_ ), .B2(_03552_ ), .ZN(_03553_ ) );
AOI21_X1 _24256_ ( .A(_03543_ ), .B1(_03553_ ), .B2(_01481_ ), .ZN(_03554_ ) );
OAI21_X1 _24257_ ( .A(_03541_ ), .B1(_03554_ ), .B2(\exu.io_in_bits_or ), .ZN(_03555_ ) );
AOI21_X1 _24258_ ( .A(_03540_ ), .B1(_03555_ ), .B2(_01613_ ), .ZN(_03556_ ) );
OAI21_X1 _24259_ ( .A(_03539_ ), .B1(_03556_ ), .B2(\exu.and_.io_is ), .ZN(_03557_ ) );
AOI221_X4 _24260_ ( .A(\exu.io_in_bits_sll ), .B1(_08771_ ), .B2(_01968_ ), .C1(_03557_ ), .C2(_01617_ ), .ZN(_03558_ ) );
NAND2_X1 _24261_ ( .A1(_03537_ ), .A2(_01441_ ), .ZN(_03559_ ) );
AOI211_X1 _24262_ ( .A(_01573_ ), .B(_03558_ ), .C1(\exu.io_in_bits_sll ), .C2(_03559_ ), .ZN(_03560_ ) );
OAI21_X1 _24263_ ( .A(_08772_ ), .B1(_01417_ ), .B2(_01421_ ), .ZN(_03561_ ) );
INV_X1 _24264_ ( .A(_01424_ ), .ZN(_03562_ ) );
AND3_X1 _24265_ ( .A1(_03561_ ), .A2(_03551_ ), .A3(_03562_ ), .ZN(_03563_ ) );
AOI21_X1 _24266_ ( .A(_03551_ ), .B1(_03561_ ), .B2(_03562_ ), .ZN(_03564_ ) );
NOR3_X1 _24267_ ( .A1(_03563_ ), .A2(_03564_ ), .A3(_01694_ ), .ZN(_03565_ ) );
OAI21_X1 _24268_ ( .A(_01571_ ), .B1(_03560_ ), .B2(_03565_ ), .ZN(_03566_ ) );
OR2_X1 _24269_ ( .A1(_09420_ ), .A2(_01342_ ), .ZN(_03567_ ) );
AOI21_X1 _24270_ ( .A(\exu.io_in_bits_jalr ), .B1(_03566_ ), .B2(_03567_ ), .ZN(_03568_ ) );
NOR2_X1 _24271_ ( .A1(_09420_ ), .A2(_01855_ ), .ZN(_03569_ ) );
OAI21_X1 _24272_ ( .A(_01501_ ), .B1(_03568_ ), .B2(_03569_ ), .ZN(_03570_ ) );
MUX2_X1 _24273_ ( .A(_03538_ ), .B(_03570_ ), .S(_01505_ ), .Z(_03571_ ) );
MUX2_X1 _24274_ ( .A(_03530_ ), .B(_03571_ ), .S(_01507_ ), .Z(_03572_ ) );
MUX2_X1 _24275_ ( .A(_03529_ ), .B(_03572_ ), .S(_01510_ ), .Z(_03573_ ) );
AOI21_X1 _24276_ ( .A(_03528_ ), .B1(_03573_ ), .B2(_01512_ ), .ZN(_03574_ ) );
AND3_X1 _24277_ ( .A1(_09383_ ), .A2(_10843_ ), .A3(\exu.andi.io_is ), .ZN(_03575_ ) );
OAI21_X1 _24278_ ( .A(_01175_ ), .B1(_03574_ ), .B2(_03575_ ), .ZN(_03576_ ) );
NAND2_X1 _24279_ ( .A1(_09387_ ), .A2(_01519_ ), .ZN(_03577_ ) );
AOI21_X1 _24280_ ( .A(_01173_ ), .B1(_03576_ ), .B2(_03577_ ), .ZN(_03578_ ) );
AND2_X1 _24281_ ( .A1(\exu.addi._io_rd_T_4 [27] ), .A2(_01523_ ), .ZN(_03579_ ) );
OAI21_X1 _24282_ ( .A(_01109_ ), .B1(_03578_ ), .B2(_03579_ ), .ZN(_03580_ ) );
INV_X1 _24283_ ( .A(_03580_ ), .ZN(_03581_ ) );
NOR3_X1 _24284_ ( .A1(_01721_ ), .A2(fanout_net_27 ), .A3(_09455_ ), .ZN(_03582_ ) );
NOR2_X1 _24285_ ( .A1(_03581_ ), .A2(_03582_ ), .ZN(_03583_ ) );
INV_X1 _24286_ ( .A(_03583_ ), .ZN(\exu.io_out_bits_rd_wdata [27] ) );
AOI211_X1 _24287_ ( .A(_01752_ ), .B(_01534_ ), .C1(_02732_ ), .C2(_02021_ ), .ZN(_03584_ ) );
OAI21_X1 _24288_ ( .A(_01878_ ), .B1(_03584_ ), .B2(_01512_ ), .ZN(_03585_ ) );
OAI21_X1 _24289_ ( .A(_01755_ ), .B1(\exu.add.io_rs1_data [26] ), .B2(\exu.addi.io_imm [26] ), .ZN(_03586_ ) );
NAND4_X1 _24290_ ( .A1(_02132_ ), .A2(_01207_ ), .A3(_01213_ ), .A4(_02283_ ), .ZN(_03587_ ) );
NAND2_X1 _24291_ ( .A1(_02756_ ), .A2(_01654_ ), .ZN(_03588_ ) );
AND2_X1 _24292_ ( .A1(_01667_ ), .A2(_01670_ ), .ZN(_03589_ ) );
MUX2_X1 _24293_ ( .A(_03589_ ), .B(_01679_ ), .S(_01306_ ), .Z(_03590_ ) );
MUX2_X1 _24294_ ( .A(_03590_ ), .B(_02138_ ), .S(_01308_ ), .Z(_03591_ ) );
OAI21_X1 _24295_ ( .A(_03588_ ), .B1(_03591_ ), .B2(_01654_ ), .ZN(_03592_ ) );
NAND2_X1 _24296_ ( .A1(_03592_ ), .A2(_01702_ ), .ZN(_03593_ ) );
NAND3_X1 _24297_ ( .A1(_01424_ ), .A2(_01575_ ), .A3(\exu.and_.io_is ), .ZN(_03594_ ) );
NAND2_X1 _24298_ ( .A1(_02732_ ), .A2(_01880_ ), .ZN(_03595_ ) );
AND3_X1 _24299_ ( .A1(_03595_ ), .A2(_01445_ ), .A3(_01536_ ), .ZN(_03596_ ) );
OAI21_X1 _24300_ ( .A(_01581_ ), .B1(\exu.add.io_rs1_data [26] ), .B2(\exu._GEN_0 [26] ), .ZN(_03597_ ) );
NAND3_X1 _24301_ ( .A1(_02132_ ), .A2(_01207_ ), .A3(_01212_ ), .ZN(_03598_ ) );
NOR2_X1 _24302_ ( .A1(_03598_ ), .A2(_01455_ ), .ZN(_03599_ ) );
NAND2_X1 _24303_ ( .A1(_03547_ ), .A2(_08772_ ), .ZN(_03600_ ) );
NAND3_X1 _24304_ ( .A1(_03549_ ), .A2(_03600_ ), .A3(_01478_ ), .ZN(_03601_ ) );
AND4_X1 _24305_ ( .A1(\exu.addi.io_imm [26] ), .A2(_01601_ ), .A3(_01602_ ), .A4(_01604_ ), .ZN(_03602_ ) );
AOI21_X1 _24306_ ( .A(_03602_ ), .B1(_08697_ ), .B2(_01607_ ), .ZN(_03603_ ) );
OAI21_X1 _24307_ ( .A(_03601_ ), .B1(_03603_ ), .B2(\exu.io_in_bits_sub ), .ZN(_03604_ ) );
AOI21_X1 _24308_ ( .A(_03599_ ), .B1(_03604_ ), .B2(_01610_ ), .ZN(_03605_ ) );
OAI21_X1 _24309_ ( .A(_03597_ ), .B1(_03605_ ), .B2(\exu.io_in_bits_or ), .ZN(_03606_ ) );
AOI21_X1 _24310_ ( .A(_03596_ ), .B1(_03606_ ), .B2(_01614_ ), .ZN(_03607_ ) );
OAI21_X1 _24311_ ( .A(_03594_ ), .B1(_03607_ ), .B2(\exu.and_.io_is ), .ZN(_03608_ ) );
AOI221_X4 _24312_ ( .A(\exu.io_in_bits_sll ), .B1(_08772_ ), .B2(_01493_ ), .C1(_03608_ ), .C2(_01618_ ), .ZN(_03609_ ) );
NAND2_X1 _24313_ ( .A1(_03592_ ), .A2(_01689_ ), .ZN(_03610_ ) );
AOI211_X1 _24314_ ( .A(_01574_ ), .B(_03609_ ), .C1(\exu.io_in_bits_sll ), .C2(_03610_ ), .ZN(_03611_ ) );
OR3_X1 _24315_ ( .A1(_01417_ ), .A2(_08772_ ), .A3(_01421_ ), .ZN(_03612_ ) );
AND3_X1 _24316_ ( .A1(_03612_ ), .A2(_01828_ ), .A3(_03561_ ), .ZN(_03613_ ) );
OAI21_X1 _24317_ ( .A(_01571_ ), .B1(_03611_ ), .B2(_03613_ ), .ZN(_03614_ ) );
NAND3_X1 _24318_ ( .A1(_08809_ ), .A2(_09452_ ), .A3(_08810_ ), .ZN(_03615_ ) );
AOI21_X1 _24319_ ( .A(\exu.io_in_bits_jalr ), .B1(_03614_ ), .B2(_03615_ ), .ZN(_03616_ ) );
AND3_X1 _24320_ ( .A1(_08809_ ), .A2(_01699_ ), .A3(_08810_ ), .ZN(_03617_ ) );
OAI21_X1 _24321_ ( .A(_01989_ ), .B1(_03616_ ), .B2(_03617_ ), .ZN(_03618_ ) );
MUX2_X1 _24322_ ( .A(_03593_ ), .B(_03618_ ), .S(_01992_ ), .Z(_03619_ ) );
MUX2_X1 _24323_ ( .A(_03587_ ), .B(_03619_ ), .S(_01705_ ), .Z(_03620_ ) );
MUX2_X1 _24324_ ( .A(_03586_ ), .B(_03620_ ), .S(_01860_ ), .Z(_03621_ ) );
AOI21_X1 _24325_ ( .A(_03585_ ), .B1(_03621_ ), .B2(_01862_ ), .ZN(_03622_ ) );
AND3_X1 _24326_ ( .A1(_09170_ ), .A2(_01864_ ), .A3(\exu.andi.io_is ), .ZN(_03623_ ) );
OAI21_X1 _24327_ ( .A(_01877_ ), .B1(_03622_ ), .B2(_03623_ ), .ZN(_03624_ ) );
NAND2_X1 _24328_ ( .A1(_09172_ ), .A2(_02000_ ), .ZN(_03625_ ) );
AOI21_X1 _24329_ ( .A(_01876_ ), .B1(_03624_ ), .B2(_03625_ ), .ZN(_03626_ ) );
AND2_X1 _24330_ ( .A1(\exu.addi._io_rd_T_4 [26] ), .A2(_02003_ ), .ZN(_03627_ ) );
OAI21_X1 _24331_ ( .A(_01875_ ), .B1(_03626_ ), .B2(_03627_ ), .ZN(_03628_ ) );
OAI211_X1 _24332_ ( .A(_01058_ ), .B(\exu.csrrs.io_csr_rdata [26] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_03629_ ) );
NAND2_X1 _24333_ ( .A1(_03628_ ), .A2(_03629_ ), .ZN(\exu.io_out_bits_rd_wdata [26] ) );
NAND2_X1 _24334_ ( .A1(_02802_ ), .A2(_02021_ ), .ZN(_03630_ ) );
NAND3_X1 _24335_ ( .A1(_03630_ ), .A2(_01914_ ), .A3(_01537_ ), .ZN(_03631_ ) );
NAND3_X1 _24336_ ( .A1(_01418_ ), .A2(_10699_ ), .A3(\exu.and_.io_is ), .ZN(_03632_ ) );
AND3_X1 _24337_ ( .A1(_03630_ ), .A2(_01445_ ), .A3(_01537_ ), .ZN(_03633_ ) );
OAI21_X1 _24338_ ( .A(_01581_ ), .B1(\exu.add.io_rs1_data [25] ), .B2(\exu._GEN_0 [25] ), .ZN(_03634_ ) );
AND3_X1 _24339_ ( .A1(_02818_ ), .A2(_01212_ ), .A3(_01594_ ), .ZN(_03635_ ) );
AND2_X1 _24340_ ( .A1(_01471_ ), .A2(_01346_ ), .ZN(_03636_ ) );
OR3_X1 _24341_ ( .A1(_03636_ ), .A2(_01345_ ), .A3(_08904_ ), .ZN(_03637_ ) );
AOI211_X1 _24342_ ( .A(_08906_ ), .B(_01597_ ), .C1(_01471_ ), .C2(_08770_ ), .ZN(_03638_ ) );
NAND2_X1 _24343_ ( .A1(_03637_ ), .A2(_03638_ ), .ZN(_03639_ ) );
AND4_X1 _24344_ ( .A1(\exu.addi.io_imm [25] ), .A2(_01601_ ), .A3(_01602_ ), .A4(_01604_ ), .ZN(_03640_ ) );
AOI21_X1 _24345_ ( .A(_03640_ ), .B1(_09292_ ), .B2(_01607_ ), .ZN(_03641_ ) );
OAI21_X1 _24346_ ( .A(_03639_ ), .B1(_03641_ ), .B2(\exu.io_in_bits_sub ), .ZN(_03642_ ) );
AOI21_X1 _24347_ ( .A(_03635_ ), .B1(_03642_ ), .B2(_01610_ ), .ZN(_03643_ ) );
OAI21_X1 _24348_ ( .A(_03634_ ), .B1(_03643_ ), .B2(\exu.io_in_bits_or ), .ZN(_03644_ ) );
AOI21_X1 _24349_ ( .A(_03633_ ), .B1(_03644_ ), .B2(_01614_ ), .ZN(_03645_ ) );
OAI21_X1 _24350_ ( .A(_03632_ ), .B1(_03645_ ), .B2(\exu.and_.io_is ), .ZN(_03646_ ) );
AOI221_X4 _24351_ ( .A(\exu.io_in_bits_sll ), .B1(_08768_ ), .B2(_01493_ ), .C1(_03646_ ), .C2(_01618_ ), .ZN(_03647_ ) );
OR2_X1 _24352_ ( .A1(_02806_ ), .A2(_02354_ ), .ZN(_03648_ ) );
AND2_X1 _24353_ ( .A1(_01806_ ), .A2(_01807_ ), .ZN(_03649_ ) );
MUX2_X1 _24354_ ( .A(_03649_ ), .B(_02617_ ), .S(_01306_ ), .Z(_03650_ ) );
MUX2_X1 _24355_ ( .A(_03650_ ), .B(_02227_ ), .S(_01308_ ), .Z(_03651_ ) );
OAI21_X1 _24356_ ( .A(_03648_ ), .B1(_01654_ ), .B2(_03651_ ), .ZN(_03652_ ) );
NAND2_X1 _24357_ ( .A1(_03652_ ), .A2(_01689_ ), .ZN(_03653_ ) );
AOI211_X1 _24358_ ( .A(_01574_ ), .B(_03647_ ), .C1(\exu.io_in_bits_sll ), .C2(_03653_ ), .ZN(_03654_ ) );
AOI21_X1 _24359_ ( .A(_01346_ ), .B1(_01399_ ), .B2(_01416_ ), .ZN(_03655_ ) );
OR3_X1 _24360_ ( .A1(_03655_ ), .A2(_08768_ ), .A3(_01419_ ), .ZN(_03656_ ) );
OAI21_X1 _24361_ ( .A(_08768_ ), .B1(_03655_ ), .B2(_01419_ ), .ZN(_03657_ ) );
AND3_X1 _24362_ ( .A1(_03656_ ), .A2(_01828_ ), .A3(_03657_ ), .ZN(_03658_ ) );
OAI21_X1 _24363_ ( .A(_01571_ ), .B1(_03654_ ), .B2(_03658_ ), .ZN(_03659_ ) );
OR2_X1 _24364_ ( .A1(_09268_ ), .A2(_01823_ ), .ZN(_03660_ ) );
AOI21_X1 _24365_ ( .A(\exu.io_in_bits_jalr ), .B1(_03659_ ), .B2(_03660_ ), .ZN(_03661_ ) );
NOR2_X1 _24366_ ( .A1(_09268_ ), .A2(_01855_ ), .ZN(_03662_ ) );
OAI21_X1 _24367_ ( .A(_01570_ ), .B1(_03661_ ), .B2(_03662_ ), .ZN(_03663_ ) );
NAND2_X1 _24368_ ( .A1(_03652_ ), .A2(_01702_ ), .ZN(_03664_ ) );
NAND3_X1 _24369_ ( .A1(_03663_ ), .A2(_01994_ ), .A3(_03664_ ), .ZN(_03665_ ) );
AND3_X1 _24370_ ( .A1(_02818_ ), .A2(_01213_ ), .A3(_02283_ ), .ZN(_03666_ ) );
OAI211_X1 _24371_ ( .A(_03665_ ), .B(_01860_ ), .C1(_01994_ ), .C2(_03666_ ), .ZN(_03667_ ) );
OAI21_X1 _24372_ ( .A(_01186_ ), .B1(\exu.add.io_rs1_data [25] ), .B2(\exu.addi.io_imm [25] ), .ZN(_03668_ ) );
AND2_X1 _24373_ ( .A1(_03668_ ), .A2(_01182_ ), .ZN(_03669_ ) );
AOI221_X4 _24374_ ( .A(\exu.andi.io_is ), .B1(\exu.io_in_bits_srai ), .B2(_03631_ ), .C1(_03667_ ), .C2(_03669_ ), .ZN(_03670_ ) );
AND3_X1 _24375_ ( .A1(_09164_ ), .A2(_01864_ ), .A3(\exu.andi.io_is ), .ZN(_03671_ ) );
OAI21_X1 _24376_ ( .A(_01877_ ), .B1(_03670_ ), .B2(_03671_ ), .ZN(_03672_ ) );
NAND2_X1 _24377_ ( .A1(_09166_ ), .A2(_02000_ ), .ZN(_03673_ ) );
AOI21_X1 _24378_ ( .A(_01876_ ), .B1(_03672_ ), .B2(_03673_ ), .ZN(_03674_ ) );
AND2_X1 _24379_ ( .A1(\exu.addi._io_rd_T_4 [25] ), .A2(_02003_ ), .ZN(_03675_ ) );
OAI21_X1 _24380_ ( .A(_01875_ ), .B1(_03674_ ), .B2(_03675_ ), .ZN(_03676_ ) );
OAI211_X1 _24381_ ( .A(_01058_ ), .B(\exu.csrrs.io_csr_rdata [25] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_03677_ ) );
NAND2_X1 _24382_ ( .A1(_03676_ ), .A2(_03677_ ), .ZN(\exu.io_out_bits_rd_wdata [25] ) );
OAI21_X1 _24383_ ( .A(_01536_ ), .B1(_02865_ ), .B2(_01568_ ), .ZN(_03678_ ) );
NOR2_X1 _24384_ ( .A1(_03678_ ), .A2(_01752_ ), .ZN(_03679_ ) );
OAI21_X1 _24385_ ( .A(_01878_ ), .B1(_03679_ ), .B2(_01512_ ), .ZN(_03680_ ) );
OAI21_X1 _24386_ ( .A(_01755_ ), .B1(\exu.add.io_rs1_data [24] ), .B2(\exu.addi.io_imm [24] ), .ZN(_03681_ ) );
NAND4_X1 _24387_ ( .A1(_02273_ ), .A2(_01207_ ), .A3(_01213_ ), .A4(_02283_ ), .ZN(_03682_ ) );
OAI21_X1 _24388_ ( .A(_01308_ ), .B1(_02290_ ), .B2(_02291_ ), .ZN(_03683_ ) );
AOI21_X1 _24389_ ( .A(_01306_ ), .B1(_01961_ ), .B2(_01962_ ), .ZN(_03684_ ) );
AND3_X1 _24390_ ( .A1(_03292_ ), .A2(_03293_ ), .A3(_01279_ ), .ZN(_03685_ ) );
OAI21_X1 _24391_ ( .A(_01271_ ), .B1(_03684_ ), .B2(_03685_ ), .ZN(_03686_ ) );
AND2_X1 _24392_ ( .A1(_03683_ ), .A2(_03686_ ), .ZN(_03687_ ) );
MUX2_X1 _24393_ ( .A(_02880_ ), .B(_03687_ ), .S(_01333_ ), .Z(_03688_ ) );
NAND2_X1 _24394_ ( .A1(_03688_ ), .A2(_01702_ ), .ZN(_03689_ ) );
NAND3_X1 _24395_ ( .A1(_01419_ ), .A2(_01575_ ), .A3(\exu.and_.io_is ), .ZN(_03690_ ) );
NOR2_X1 _24396_ ( .A1(_03678_ ), .A2(_01579_ ), .ZN(_03691_ ) );
OAI21_X1 _24397_ ( .A(_01581_ ), .B1(\exu.add.io_rs1_data [24] ), .B2(\exu._GEN_0 [24] ), .ZN(_03692_ ) );
AND3_X1 _24398_ ( .A1(_02273_ ), .A2(_01207_ ), .A3(_01450_ ), .ZN(_03693_ ) );
AND2_X1 _24399_ ( .A1(_03693_ ), .A2(_01594_ ), .ZN(_03694_ ) );
AOI21_X1 _24400_ ( .A(_01597_ ), .B1(_01471_ ), .B2(_01346_ ), .ZN(_03695_ ) );
OAI21_X1 _24401_ ( .A(_03695_ ), .B1(_01346_ ), .B2(_01471_ ), .ZN(_03696_ ) );
AND4_X1 _24402_ ( .A1(\exu.addi.io_imm [24] ), .A2(_01600_ ), .A3(_01463_ ), .A4(_01603_ ), .ZN(_03697_ ) );
AOI21_X1 _24403_ ( .A(_03697_ ), .B1(_09614_ ), .B2(_01606_ ), .ZN(_03698_ ) );
OAI21_X1 _24404_ ( .A(_03696_ ), .B1(_03698_ ), .B2(\exu.io_in_bits_sub ), .ZN(_03699_ ) );
AOI21_X1 _24405_ ( .A(_03694_ ), .B1(_03699_ ), .B2(_01481_ ), .ZN(_03700_ ) );
OAI21_X1 _24406_ ( .A(_03692_ ), .B1(_03700_ ), .B2(\exu.io_in_bits_or ), .ZN(_03701_ ) );
AOI21_X1 _24407_ ( .A(_03691_ ), .B1(_03701_ ), .B2(_01613_ ), .ZN(_03702_ ) );
OAI21_X1 _24408_ ( .A(_03690_ ), .B1(_03702_ ), .B2(\exu.and_.io_is ), .ZN(_03703_ ) );
AOI221_X4 _24409_ ( .A(\exu.io_in_bits_sll ), .B1(_08769_ ), .B2(_01968_ ), .C1(_03703_ ), .C2(_01618_ ), .ZN(_03704_ ) );
NAND2_X1 _24410_ ( .A1(_03688_ ), .A2(_01689_ ), .ZN(_03705_ ) );
AOI211_X1 _24411_ ( .A(_01574_ ), .B(_03704_ ), .C1(\exu.io_in_bits_sll ), .C2(_03705_ ), .ZN(_03706_ ) );
NAND3_X1 _24412_ ( .A1(_01399_ ), .A2(_01346_ ), .A3(_01416_ ), .ZN(_03707_ ) );
NOR2_X1 _24413_ ( .A1(_03655_ ), .A2(_01694_ ), .ZN(_03708_ ) );
AOI21_X1 _24414_ ( .A(_03706_ ), .B1(_03707_ ), .B2(_03708_ ), .ZN(_03709_ ) );
OAI221_X1 _24415_ ( .A(_01341_ ), .B1(_01823_ ), .B2(_09619_ ), .C1(_03709_ ), .C2(\exu.io_in_bits_jal ), .ZN(_03710_ ) );
AND2_X1 _24416_ ( .A1(_09617_ ), .A2(_01699_ ), .ZN(_03711_ ) );
OAI211_X1 _24417_ ( .A(_03710_ ), .B(_01989_ ), .C1(_01854_ ), .C2(_03711_ ), .ZN(_03712_ ) );
MUX2_X1 _24418_ ( .A(_03689_ ), .B(_03712_ ), .S(_01992_ ), .Z(_03713_ ) );
MUX2_X1 _24419_ ( .A(_03682_ ), .B(_03713_ ), .S(_01705_ ), .Z(_03714_ ) );
MUX2_X1 _24420_ ( .A(_03681_ ), .B(_03714_ ), .S(_01860_ ), .Z(_03715_ ) );
AOI21_X1 _24421_ ( .A(_03680_ ), .B1(_03715_ ), .B2(_01862_ ), .ZN(_03716_ ) );
AND3_X1 _24422_ ( .A1(_09161_ ), .A2(_01864_ ), .A3(\exu.andi.io_is ), .ZN(_03717_ ) );
OAI21_X1 _24423_ ( .A(_01877_ ), .B1(_03716_ ), .B2(_03717_ ), .ZN(_03718_ ) );
NAND2_X1 _24424_ ( .A1(_09163_ ), .A2(_02000_ ), .ZN(_03719_ ) );
AOI21_X1 _24425_ ( .A(_01876_ ), .B1(_03718_ ), .B2(_03719_ ), .ZN(_03720_ ) );
AND2_X1 _24426_ ( .A1(\exu.addi._io_rd_T_4 [24] ), .A2(_02003_ ), .ZN(_03721_ ) );
OAI21_X1 _24427_ ( .A(_01875_ ), .B1(_03720_ ), .B2(_03721_ ), .ZN(_03722_ ) );
OAI211_X1 _24428_ ( .A(_10845_ ), .B(\exu.csrrs.io_csr_rdata [24] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_03723_ ) );
NAND2_X1 _24429_ ( .A1(_03722_ ), .A2(_03723_ ), .ZN(\exu.io_out_bits_rd_wdata [24] ) );
OAI21_X1 _24430_ ( .A(_01536_ ), .B1(_02929_ ), .B2(_01568_ ), .ZN(_03724_ ) );
NOR2_X1 _24431_ ( .A1(_03724_ ), .A2(_01752_ ), .ZN(_03725_ ) );
OAI21_X1 _24432_ ( .A(_01515_ ), .B1(_03725_ ), .B2(_01182_ ), .ZN(_03726_ ) );
OAI21_X1 _24433_ ( .A(_01755_ ), .B1(\exu.add.io_rs1_data [23] ), .B2(\exu.addi.io_imm [23] ), .ZN(_03727_ ) );
OR3_X1 _24434_ ( .A1(_02933_ ), .A2(_01795_ ), .A3(_01797_ ), .ZN(_03728_ ) );
AOI21_X1 _24435_ ( .A(_01271_ ), .B1(_01269_ ), .B2(_01280_ ), .ZN(_03729_ ) );
AOI21_X1 _24436_ ( .A(_03729_ ), .B1(_01327_ ), .B2(_01686_ ), .ZN(_03730_ ) );
MUX2_X1 _24437_ ( .A(_03730_ ), .B(_02945_ ), .S(_01804_ ), .Z(_03731_ ) );
NAND2_X1 _24438_ ( .A1(_03731_ ), .A2(_01338_ ), .ZN(_03732_ ) );
NAND3_X1 _24439_ ( .A1(_01409_ ), .A2(_10698_ ), .A3(\exu.and_.io_is ), .ZN(_03733_ ) );
NOR2_X1 _24440_ ( .A1(_03724_ ), .A2(_01579_ ), .ZN(_03734_ ) );
OAI21_X1 _24441_ ( .A(_01448_ ), .B1(\exu.add.io_rs1_data [23] ), .B2(\exu._GEN_0 [23] ), .ZN(_03735_ ) );
NOR3_X1 _24442_ ( .A1(_02933_ ), .A2(_01794_ ), .A3(_01455_ ), .ZN(_03736_ ) );
AOI21_X1 _24443_ ( .A(_08897_ ), .B1(_01836_ ), .B2(_08758_ ), .ZN(_03737_ ) );
NOR2_X1 _24444_ ( .A1(_03737_ ), .A2(_08752_ ), .ZN(_03738_ ) );
INV_X1 _24445_ ( .A(_03738_ ), .ZN(_03739_ ) );
AND3_X1 _24446_ ( .A1(_03739_ ), .A2(_08751_ ), .A3(_08889_ ), .ZN(_03740_ ) );
AOI21_X1 _24447_ ( .A(_08751_ ), .B1(_03739_ ), .B2(_08889_ ), .ZN(_03741_ ) );
OR3_X1 _24448_ ( .A1(_03740_ ), .A2(_03741_ ), .A3(_01597_ ), .ZN(_03742_ ) );
AND4_X1 _24449_ ( .A1(\exu.addi.io_imm [23] ), .A2(_01600_ ), .A3(_01463_ ), .A4(_01603_ ), .ZN(_03743_ ) );
AOI21_X1 _24450_ ( .A(_03743_ ), .B1(_09482_ ), .B2(_01606_ ), .ZN(_03744_ ) );
OAI21_X1 _24451_ ( .A(_03742_ ), .B1(_03744_ ), .B2(\exu.io_in_bits_sub ), .ZN(_03745_ ) );
AOI21_X1 _24452_ ( .A(_03736_ ), .B1(_03745_ ), .B2(_01481_ ), .ZN(_03746_ ) );
OAI21_X1 _24453_ ( .A(_03735_ ), .B1(_03746_ ), .B2(\exu.io_in_bits_or ), .ZN(_03747_ ) );
AOI21_X1 _24454_ ( .A(_03734_ ), .B1(_03747_ ), .B2(_01613_ ), .ZN(_03748_ ) );
OAI21_X1 _24455_ ( .A(_03733_ ), .B1(_03748_ ), .B2(\exu.and_.io_is ), .ZN(_03749_ ) );
AOI221_X4 _24456_ ( .A(\exu.io_in_bits_sll ), .B1(_08751_ ), .B2(_01968_ ), .C1(_03749_ ), .C2(_01618_ ), .ZN(_03750_ ) );
NAND2_X1 _24457_ ( .A1(_03731_ ), .A2(_01441_ ), .ZN(_03751_ ) );
AOI211_X1 _24458_ ( .A(_01573_ ), .B(_03750_ ), .C1(\exu.io_in_bits_sll ), .C2(_03751_ ), .ZN(_03752_ ) );
INV_X1 _24459_ ( .A(_08752_ ), .ZN(_03753_ ) );
NOR4_X1 _24460_ ( .A1(_01391_ ), .A2(_08747_ ), .A3(_08749_ ), .A4(_01403_ ), .ZN(_03754_ ) );
OAI211_X1 _24461_ ( .A(_08757_ ), .B(_08754_ ), .C1(_03754_ ), .C2(_01407_ ), .ZN(_03755_ ) );
AOI21_X1 _24462_ ( .A(_03753_ ), .B1(_03755_ ), .B2(_01412_ ), .ZN(_03756_ ) );
OR3_X1 _24463_ ( .A1(_03756_ ), .A2(_08751_ ), .A3(_01414_ ), .ZN(_03757_ ) );
OAI21_X1 _24464_ ( .A(_08751_ ), .B1(_03756_ ), .B2(_01414_ ), .ZN(_03758_ ) );
AND3_X1 _24465_ ( .A1(_03757_ ), .A2(_01828_ ), .A3(_03758_ ), .ZN(_03759_ ) );
OAI21_X1 _24466_ ( .A(_01571_ ), .B1(_03752_ ), .B2(_03759_ ), .ZN(_03760_ ) );
OR2_X1 _24467_ ( .A1(_09485_ ), .A2(_01342_ ), .ZN(_03761_ ) );
AOI21_X1 _24468_ ( .A(\exu.io_in_bits_jalr ), .B1(_03760_ ), .B2(_03761_ ), .ZN(_03762_ ) );
NOR2_X1 _24469_ ( .A1(_09485_ ), .A2(_01855_ ), .ZN(_03763_ ) );
OAI21_X1 _24470_ ( .A(_01989_ ), .B1(_03762_ ), .B2(_03763_ ), .ZN(_03764_ ) );
MUX2_X1 _24471_ ( .A(_03732_ ), .B(_03764_ ), .S(_01505_ ), .Z(_03765_ ) );
MUX2_X1 _24472_ ( .A(_03728_ ), .B(_03765_ ), .S(_01705_ ), .Z(_03766_ ) );
MUX2_X1 _24473_ ( .A(_03727_ ), .B(_03766_ ), .S(_01860_ ), .Z(_03767_ ) );
AOI21_X1 _24474_ ( .A(_03726_ ), .B1(_03767_ ), .B2(_01862_ ), .ZN(_03768_ ) );
AND3_X1 _24475_ ( .A1(_09139_ ), .A2(_01864_ ), .A3(\exu.andi.io_is ), .ZN(_03769_ ) );
OAI21_X1 _24476_ ( .A(_01723_ ), .B1(_03768_ ), .B2(_03769_ ), .ZN(_03770_ ) );
NAND2_X1 _24477_ ( .A1(_09141_ ), .A2(_01519_ ), .ZN(_03771_ ) );
AOI21_X1 _24478_ ( .A(_01173_ ), .B1(_03770_ ), .B2(_03771_ ), .ZN(_03772_ ) );
AND2_X1 _24479_ ( .A1(\exu.addi._io_rd_T_4 [23] ), .A2(_01523_ ), .ZN(_03773_ ) );
OAI21_X1 _24480_ ( .A(_01109_ ), .B1(_03772_ ), .B2(_03773_ ), .ZN(_03774_ ) );
OAI211_X1 _24481_ ( .A(_01873_ ), .B(\exu.csrrs.io_csr_rdata [23] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_03775_ ) );
NAND2_X1 _24482_ ( .A1(_03774_ ), .A2(_03775_ ), .ZN(\exu.io_out_bits_rd_wdata [23] ) );
OAI211_X1 _24483_ ( .A(_02985_ ), .B(_01880_ ), .C1(_01881_ ), .C2(_01563_ ), .ZN(_03776_ ) );
AND3_X1 _24484_ ( .A1(_03776_ ), .A2(_01914_ ), .A3(_01537_ ), .ZN(_03777_ ) );
OAI21_X1 _24485_ ( .A(_01878_ ), .B1(_03777_ ), .B2(_01512_ ), .ZN(_03778_ ) );
OAI21_X1 _24486_ ( .A(_01755_ ), .B1(\exu.add.io_rs1_data [22] ), .B2(\exu.addi.io_imm [22] ), .ZN(_03779_ ) );
OAI21_X1 _24487_ ( .A(_03005_ ), .B1(_02435_ ), .B2(_01935_ ), .ZN(_03780_ ) );
NAND3_X1 _24488_ ( .A1(_03780_ ), .A2(_01213_ ), .A3(_02283_ ), .ZN(_03781_ ) );
NAND3_X1 _24489_ ( .A1(_01644_ ), .A2(_01308_ ), .A3(_01651_ ), .ZN(_03782_ ) );
OAI21_X1 _24490_ ( .A(_03782_ ), .B1(_01672_ ), .B2(_01308_ ), .ZN(_03783_ ) );
MUX2_X1 _24491_ ( .A(_03783_ ), .B(_03008_ ), .S(_01804_ ), .Z(_03784_ ) );
NAND2_X1 _24492_ ( .A1(_03784_ ), .A2(_01702_ ), .ZN(_03785_ ) );
NAND3_X1 _24493_ ( .A1(_01414_ ), .A2(_01575_ ), .A3(\exu.and_.io_is ), .ZN(_03786_ ) );
AND3_X1 _24494_ ( .A1(_03776_ ), .A2(_01445_ ), .A3(_01536_ ), .ZN(_03787_ ) );
OAI21_X1 _24495_ ( .A(_01581_ ), .B1(\exu.add.io_rs1_data [22] ), .B2(\exu._GEN_0 [22] ), .ZN(_03788_ ) );
AND3_X1 _24496_ ( .A1(_03780_ ), .A2(_01212_ ), .A3(_01594_ ), .ZN(_03789_ ) );
NAND2_X1 _24497_ ( .A1(_03737_ ), .A2(_08752_ ), .ZN(_03790_ ) );
NAND3_X1 _24498_ ( .A1(_03739_ ), .A2(_01478_ ), .A3(_03790_ ), .ZN(_03791_ ) );
AND4_X1 _24499_ ( .A1(\exu.addi.io_imm [22] ), .A2(_01601_ ), .A3(_01602_ ), .A4(_01604_ ), .ZN(_03792_ ) );
AOI21_X1 _24500_ ( .A(_03792_ ), .B1(_09526_ ), .B2(_01607_ ), .ZN(_03793_ ) );
OAI21_X1 _24501_ ( .A(_03791_ ), .B1(_03793_ ), .B2(\exu.io_in_bits_sub ), .ZN(_03794_ ) );
AOI21_X1 _24502_ ( .A(_03789_ ), .B1(_03794_ ), .B2(_01610_ ), .ZN(_03795_ ) );
OAI21_X1 _24503_ ( .A(_03788_ ), .B1(_03795_ ), .B2(\exu.io_in_bits_or ), .ZN(_03796_ ) );
AOI21_X1 _24504_ ( .A(_03787_ ), .B1(_03796_ ), .B2(_01614_ ), .ZN(_03797_ ) );
OAI21_X1 _24505_ ( .A(_03786_ ), .B1(_03797_ ), .B2(\exu.and_.io_is ), .ZN(_03798_ ) );
AOI221_X4 _24506_ ( .A(\exu.io_in_bits_sll ), .B1(_08752_ ), .B2(_01493_ ), .C1(_03798_ ), .C2(_01618_ ), .ZN(_03799_ ) );
NAND2_X1 _24507_ ( .A1(_03784_ ), .A2(_01689_ ), .ZN(_03800_ ) );
AOI211_X1 _24508_ ( .A(_01574_ ), .B(_03799_ ), .C1(\exu.io_in_bits_sll ), .C2(_03800_ ), .ZN(_03801_ ) );
AND3_X1 _24509_ ( .A1(_03755_ ), .A2(_03753_ ), .A3(_01412_ ), .ZN(_03802_ ) );
NOR3_X1 _24510_ ( .A1(_03756_ ), .A2(_01694_ ), .A3(_03802_ ), .ZN(_03803_ ) );
OAI21_X1 _24511_ ( .A(_01571_ ), .B1(_03801_ ), .B2(_03803_ ), .ZN(_03804_ ) );
NAND2_X1 _24512_ ( .A1(_09529_ ), .A2(_09452_ ), .ZN(_03805_ ) );
AOI21_X1 _24513_ ( .A(\exu.io_in_bits_jalr ), .B1(_03804_ ), .B2(_03805_ ), .ZN(_03806_ ) );
AND2_X1 _24514_ ( .A1(_09529_ ), .A2(_01699_ ), .ZN(_03807_ ) );
OAI21_X1 _24515_ ( .A(_01989_ ), .B1(_03806_ ), .B2(_03807_ ), .ZN(_03808_ ) );
MUX2_X1 _24516_ ( .A(_03785_ ), .B(_03808_ ), .S(_01992_ ), .Z(_03809_ ) );
MUX2_X1 _24517_ ( .A(_03781_ ), .B(_03809_ ), .S(_01994_ ), .Z(_03810_ ) );
MUX2_X1 _24518_ ( .A(_03779_ ), .B(_03810_ ), .S(_01860_ ), .Z(_03811_ ) );
AOI21_X1 _24519_ ( .A(_03778_ ), .B1(_03811_ ), .B2(_01862_ ), .ZN(_03812_ ) );
AND3_X1 _24520_ ( .A1(_09142_ ), .A2(_10844_ ), .A3(\exu.andi.io_is ), .ZN(_03813_ ) );
OAI21_X1 _24521_ ( .A(_01877_ ), .B1(_03812_ ), .B2(_03813_ ), .ZN(_03814_ ) );
NAND2_X1 _24522_ ( .A1(_09144_ ), .A2(_02000_ ), .ZN(_03815_ ) );
AOI21_X1 _24523_ ( .A(_01876_ ), .B1(_03814_ ), .B2(_03815_ ), .ZN(_03816_ ) );
NOR3_X1 _24524_ ( .A1(_09553_ ), .A2(_09514_ ), .A3(_02249_ ), .ZN(_03817_ ) );
OAI21_X1 _24525_ ( .A(_01875_ ), .B1(_03816_ ), .B2(_03817_ ), .ZN(_03818_ ) );
OAI211_X1 _24526_ ( .A(_01058_ ), .B(\exu.csrrs.io_csr_rdata [22] ), .C1(\exu.csrrs.io_is ), .C2(\exu.csrrw.io_is ), .ZN(_03819_ ) );
NAND2_X1 _24527_ ( .A1(_03818_ ), .A2(_03819_ ), .ZN(\exu.io_out_bits_rd_wdata [22] ) );
OR3_X1 _24528_ ( .A1(\exu.io_in_bits_sb ), .A2(\exu.io_in_bits_sh ), .A3(\exu.io_in_bits_sw ), .ZN(\exu.io_out_bits_wen ) );
AND2_X1 _24529_ ( .A1(_09399_ ), .A2(_09403_ ), .ZN(\ifu.io_out_bits_pc [28] ) );
AOI211_X1 _24530_ ( .A(_11580_ ), .B(_11540_ ), .C1(_11582_ ), .C2(_11584_ ), .ZN(\icache.icache_reg_1_3_$_SDFFE_PP0P__Q_E ) );
AND3_X1 _24531_ ( .A1(_11561_ ), .A2(_11562_ ), .A3(_11523_ ), .ZN(\icache.offset_buf_$_OR__A_Y_$_ANDNOT__B_Y ) );
AND2_X1 _24532_ ( .A1(\arbiter._clink_io_axi_araddr_T ), .A2(io_master_arready ), .ZN(_03820_ ) );
AND2_X1 _24533_ ( .A1(_01057_ ), .A2(_03820_ ), .ZN(_03821_ ) );
NOR3_X1 _24534_ ( .A1(_12017_ ), .A2(_12020_ ), .A3(_11495_ ), .ZN(_03822_ ) );
INV_X1 _24535_ ( .A(_03822_ ), .ZN(_03823_ ) );
NAND3_X1 _24536_ ( .A1(_03823_ ), .A2(\icache._io_out_arvalid_T ), .A3(_12048_ ), .ZN(_03824_ ) );
NAND2_X1 _24537_ ( .A1(_10992_ ), .A2(\icache._io_out_arvalid_T_2 ), .ZN(_03825_ ) );
AOI21_X1 _24538_ ( .A(_03821_ ), .B1(_03824_ ), .B2(_03825_ ), .ZN(\icache.state_$_DFF_P__Q_1_D ) );
OAI22_X1 _24539_ ( .A1(_03822_ ), .A2(_12020_ ), .B1(fanout_net_27 ), .B2(\icache._io_out_arvalid_T ), .ZN(_03826_ ) );
OAI21_X1 _24540_ ( .A(_03826_ ), .B1(fanout_net_27 ), .B2(_11944_ ), .ZN(\icache.state_$_DFF_P__Q_2_D ) );
NAND4_X1 _24541_ ( .A1(_03823_ ), .A2(\icache._io_out_arvalid_T ), .A3(_12048_ ), .A4(_03821_ ), .ZN(_03827_ ) );
NAND3_X1 _24542_ ( .A1(_12201_ ), .A2(_11892_ ), .A3(\icache._icache_reg_T ), .ZN(_03828_ ) );
NAND4_X1 _24543_ ( .A1(_01057_ ), .A2(_10922_ ), .A3(\icache._io_out_arvalid_T_2 ), .A4(_03820_ ), .ZN(_03829_ ) );
NAND3_X1 _24544_ ( .A1(_03827_ ), .A2(_03828_ ), .A3(_03829_ ), .ZN(\icache.state_$_DFF_P__Q_D ) );
AOI211_X1 _24545_ ( .A(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__A_Y ), .B(_11944_ ), .C1(_11582_ ), .C2(_11584_ ), .ZN(\icache.valid_reg_1_$_MUX__A_Y_$_OR__B_A_$_ANDNOT__A_Y ) );
AOI211_X1 _24546_ ( .A(\arbiter.io_ifu_araddr [4] ), .B(_11944_ ), .C1(_11582_ ), .C2(_11584_ ), .ZN(\icache.valid_reg_1_$_MUX__A_Y_$_OR__B_A_$_ANDNOT__A_1_Y ) );
OR2_X1 _24547_ ( .A1(_11165_ ), .A2(_11167_ ), .ZN(\idu._io_out_bits_csr_waddr_T_16 [0] ) );
INV_X1 _24548_ ( .A(_11077_ ), .ZN(\idu.io_out_bits_imm [0] ) );
INV_X1 _24549_ ( .A(_11086_ ), .ZN(\idu.io_out_bits_imm [3] ) );
INV_X1 _24550_ ( .A(_11066_ ), .ZN(\idu.io_out_bits_imm [2] ) );
NOR2_X1 _24551_ ( .A1(_11021_ ), .A2(_10583_ ), .ZN(\idu.io_out_bits_imm [5] ) );
AOI21_X1 _24552_ ( .A(_11131_ ), .B1(_11017_ ), .B2(_11020_ ), .ZN(\idu.io_out_bits_imm [7] ) );
NOR2_X1 _24553_ ( .A1(_11021_ ), .A2(_11134_ ), .ZN(\idu.io_out_bits_imm [6] ) );
OAI211_X1 _24554_ ( .A(_11035_ ), .B(_11044_ ), .C1(_11015_ ), .C2(_10588_ ), .ZN(\idu.io_out_bits_imm [14] ) );
OAI211_X1 _24555_ ( .A(_11035_ ), .B(_11043_ ), .C1(_11015_ ), .C2(_10588_ ), .ZN(\idu.io_out_bits_imm [12] ) );
AOI21_X1 _24556_ ( .A(_10588_ ), .B1(_11021_ ), .B2(_11037_ ), .ZN(\idu.io_out_bits_imm [31] ) );
AND2_X1 _24557_ ( .A1(_11034_ ), .A2(_11091_ ), .ZN(_03830_ ) );
AND2_X2 _24558_ ( .A1(_11033_ ), .A2(_03830_ ), .ZN(_03831_ ) );
OAI211_X1 _24559_ ( .A(_03831_ ), .B(_11107_ ), .C1(_10591_ ), .C2(_11037_ ), .ZN(\idu.io_out_bits_imm [30] ) );
INV_X1 _24560_ ( .A(_11093_ ), .ZN(\idu.io_out_bits_imm [29] ) );
NAND4_X1 _24561_ ( .A1(_11033_ ), .A2(_11107_ ), .A3(_03830_ ), .A4(_11109_ ), .ZN(\idu.io_out_bits_imm [28] ) );
OAI211_X1 _24562_ ( .A(_03831_ ), .B(_11107_ ), .C1(_11131_ ), .C2(_11037_ ), .ZN(\idu.io_out_bits_imm [27] ) );
NAND4_X1 _24563_ ( .A1(_11033_ ), .A2(_11107_ ), .A3(_03830_ ), .A4(_11108_ ), .ZN(\idu.io_out_bits_imm [26] ) );
NAND3_X1 _24564_ ( .A1(_03831_ ), .A2(_11107_ ), .A3(_11110_ ), .ZN(\idu.io_out_bits_imm [25] ) );
BUF_X2 _24565_ ( .A(_11050_ ), .Z(_03832_ ) );
BUF_X2 _24566_ ( .A(_03832_ ), .Z(_03833_ ) );
BUF_X2 _24567_ ( .A(_03833_ ), .Z(_03834_ ) );
BUF_X2 _24568_ ( .A(_03834_ ), .Z(_03835_ ) );
BUF_X2 _24569_ ( .A(_03835_ ), .Z(_03836_ ) );
BUF_X4 _24570_ ( .A(_03836_ ), .Z(_03837_ ) );
BUF_X2 _24571_ ( .A(_03837_ ), .Z(_03838_ ) );
OAI211_X1 _24572_ ( .A(_03831_ ), .B(_11107_ ), .C1(_03838_ ), .C2(_11037_ ), .ZN(\idu.io_out_bits_imm [24] ) );
OAI211_X1 _24573_ ( .A(_03831_ ), .B(_11107_ ), .C1(_11062_ ), .C2(_11037_ ), .ZN(\idu.io_out_bits_imm [23] ) );
OAI21_X1 _24574_ ( .A(\idu.immI [2] ), .B1(\idu.io_out_bits_lui ), .B2(\idu.io_out_bits_auipc ), .ZN(_03839_ ) );
NAND4_X1 _24575_ ( .A1(_11033_ ), .A2(_11107_ ), .A3(_03830_ ), .A4(_03839_ ), .ZN(\idu.io_out_bits_imm [22] ) );
OAI211_X1 _24576_ ( .A(_03831_ ), .B(_11107_ ), .C1(_11067_ ), .C2(_11037_ ), .ZN(\idu.io_out_bits_imm [21] ) );
OAI211_X1 _24577_ ( .A(_10694_ ), .B(\idu.immI [0] ), .C1(_10994_ ), .C2(_11036_ ), .ZN(_03840_ ) );
NAND4_X1 _24578_ ( .A1(_11033_ ), .A2(_11035_ ), .A3(_11091_ ), .A4(_03840_ ), .ZN(\idu.io_out_bits_imm [20] ) );
INV_X1 _24579_ ( .A(_11103_ ), .ZN(\idu.io_out_bits_imm [19] ) );
OAI221_X1 _24580_ ( .A(_11035_ ), .B1(_10601_ ), .B2(_11038_ ), .C1(_11015_ ), .C2(_10588_ ), .ZN(\idu.io_out_bits_imm [18] ) );
OAI221_X1 _24581_ ( .A(_11035_ ), .B1(_10598_ ), .B2(_11038_ ), .C1(_11015_ ), .C2(_10588_ ), .ZN(\idu.io_out_bits_imm [17] ) );
OAI21_X1 _24582_ ( .A(_11106_ ), .B1(_10588_ ), .B2(_11015_ ), .ZN(\idu.io_out_bits_imm [16] ) );
AND2_X1 _24583_ ( .A1(_11001_ ), .A2(_11036_ ), .ZN(_03841_ ) );
CLKBUF_X2 _24584_ ( .A(_03841_ ), .Z(_03842_ ) );
AND4_X1 _24585_ ( .A1(_10653_ ), .A2(_03842_ ), .A3(_10654_ ), .A4(_10695_ ), .ZN(\idu.io_out_bits_add ) );
AND2_X1 _24586_ ( .A1(_10995_ ), .A2(_10695_ ), .ZN(\idu.io_out_bits_addi ) );
AND4_X1 _24587_ ( .A1(_10653_ ), .A2(_03842_ ), .A3(_10654_ ), .A4(_10680_ ), .ZN(\idu.io_out_bits_and ) );
AND2_X1 _24588_ ( .A1(_10995_ ), .A2(_10680_ ), .ZN(\idu.io_out_bits_andi ) );
AND2_X1 _24589_ ( .A1(_10998_ ), .A2(_10695_ ), .ZN(\idu.io_out_bits_lb ) );
AND2_X1 _24590_ ( .A1(_10998_ ), .A2(_10671_ ), .ZN(\idu.io_out_bits_lbu ) );
AND4_X1 _24591_ ( .A1(_10624_ ), .A2(_11001_ ), .A3(_10634_ ), .A4(_10638_ ), .ZN(\idu.io_out_bits_lh ) );
AND4_X1 _24592_ ( .A1(\idu.io_in_bits_inst [14] ), .A2(_11001_ ), .A3(_10634_ ), .A4(_10638_ ), .ZN(\idu.io_out_bits_lhu ) );
AND4_X1 _24593_ ( .A1(_10653_ ), .A2(_03842_ ), .A3(_10654_ ), .A4(_10670_ ), .ZN(\idu.io_out_bits_or ) );
AND2_X1 _24594_ ( .A1(_10995_ ), .A2(_10670_ ), .ZN(\idu.io_out_bits_ori ) );
AND4_X1 _24595_ ( .A1(_10653_ ), .A2(_03842_ ), .A3(_10654_ ), .A4(_10681_ ), .ZN(\idu.io_out_bits_sll ) );
AND4_X1 _24596_ ( .A1(_10653_ ), .A2(_10995_ ), .A3(_10654_ ), .A4(_10681_ ), .ZN(\idu.io_out_bits_slli ) );
AND4_X1 _24597_ ( .A1(_10653_ ), .A2(_03842_ ), .A3(_10654_ ), .A4(_10996_ ), .ZN(\idu.io_out_bits_slt ) );
AND2_X1 _24598_ ( .A1(_10654_ ), .A2(_10653_ ), .ZN(_03843_ ) );
AND3_X1 _24599_ ( .A1(_03843_ ), .A2(_10999_ ), .A3(_03842_ ), .ZN(\idu.io_out_bits_sltu ) );
NAND3_X1 _24600_ ( .A1(_11001_ ), .A2(_10674_ ), .A3(_11036_ ), .ZN(_03844_ ) );
NOR3_X1 _24601_ ( .A1(_11011_ ), .A2(_10608_ ), .A3(_10610_ ), .ZN(_03845_ ) );
NAND2_X1 _24602_ ( .A1(_10584_ ), .A2(_03845_ ), .ZN(_03846_ ) );
NOR2_X1 _24603_ ( .A1(_03844_ ), .A2(_03846_ ), .ZN(\idu.io_out_bits_sra ) );
NAND4_X1 _24604_ ( .A1(_03842_ ), .A2(_10653_ ), .A3(_10654_ ), .A4(_10674_ ), .ZN(_03847_ ) );
INV_X1 _24605_ ( .A(_03847_ ), .ZN(\idu.io_out_bits_srl ) );
NAND3_X1 _24606_ ( .A1(_11001_ ), .A2(_10695_ ), .A3(_11036_ ), .ZN(_03848_ ) );
NOR2_X1 _24607_ ( .A1(_03848_ ), .A2(_03846_ ), .ZN(\idu.io_out_bits_sub ) );
AND3_X1 _24608_ ( .A1(_03843_ ), .A2(_10671_ ), .A3(_03841_ ), .ZN(\idu.io_out_bits_xor ) );
AND2_X1 _24609_ ( .A1(_10788_ ), .A2(_10822_ ), .ZN(_03849_ ) );
INV_X1 _24610_ ( .A(_03849_ ), .ZN(\idu.io_raw ) );
BUF_X4 _24611_ ( .A(_10574_ ), .Z(_03850_ ) );
BUF_X4 _24612_ ( .A(_03850_ ), .Z(_03851_ ) );
OAI21_X1 _24613_ ( .A(\ifu.ren_REG_$_DFF_P__Q_D_$_NAND__Y_B ), .B1(_03851_ ), .B2(\idu.io_in_valid ), .ZN(\idu.rs_reg_$_DFF_P__Q_D ) );
AND3_X1 _24614_ ( .A1(_10818_ ), .A2(\exu.io_in_bits_wen_rd ), .A3(_10819_ ), .ZN(_03852_ ) );
INV_X1 _24615_ ( .A(_03852_ ), .ZN(_03853_ ) );
AOI21_X1 _24616_ ( .A(_03853_ ), .B1(_09013_ ), .B2(_09034_ ), .ZN(_03854_ ) );
AND2_X1 _24617_ ( .A1(_10805_ ), .A2(_03854_ ), .ZN(_03855_ ) );
INV_X1 _24618_ ( .A(_03855_ ), .ZN(_03856_ ) );
BUF_X4 _24619_ ( .A(_03856_ ), .Z(_03857_ ) );
NOR2_X1 _24620_ ( .A1(_01528_ ), .A2(_03857_ ), .ZN(_03858_ ) );
BUF_X4 _24621_ ( .A(_03855_ ), .Z(_03859_ ) );
INV_X1 _24622_ ( .A(\io_master_awaddr [25] ), .ZN(_03860_ ) );
NAND2_X1 _24623_ ( .A1(_08542_ ), .A2(_08541_ ), .ZN(_03861_ ) );
AND4_X1 _24624_ ( .A1(_03860_ ), .A2(_08535_ ), .A3(_03861_ ), .A4(_08545_ ), .ZN(_03862_ ) );
NAND2_X1 _24625_ ( .A1(_03862_ ), .A2(_08556_ ), .ZN(_03863_ ) );
AND2_X1 _24626_ ( .A1(\io_master_awaddr [9] ), .A2(\io_master_awaddr [6] ), .ZN(_03864_ ) );
NAND3_X1 _24627_ ( .A1(_03864_ ), .A2(\io_master_awaddr [8] ), .A3(\io_master_awaddr [7] ), .ZN(_03865_ ) );
INV_X1 _24628_ ( .A(\io_master_awaddr [13] ), .ZN(_03866_ ) );
INV_X1 _24629_ ( .A(\io_master_awaddr [10] ), .ZN(_03867_ ) );
NOR3_X1 _24630_ ( .A1(_03865_ ), .A2(_03866_ ), .A3(_03867_ ), .ZN(_03868_ ) );
NAND3_X1 _24631_ ( .A1(_03868_ ), .A2(\io_master_awaddr [12] ), .A3(\io_master_awaddr [11] ), .ZN(_03869_ ) );
NAND4_X1 _24632_ ( .A1(\io_master_awaddr [5] ), .A2(\io_master_awaddr [4] ), .A3(\io_master_awaddr [3] ), .A4(fanout_net_16 ), .ZN(_03870_ ) );
NAND2_X1 _24633_ ( .A1(\io_master_awaddr [0] ), .A2(\io_master_awaddr [27] ), .ZN(_03871_ ) );
INV_X1 _24634_ ( .A(\io_master_awaddr [1] ), .ZN(_03872_ ) );
NOR4_X1 _24635_ ( .A1(_03870_ ), .A2(_03871_ ), .A3(_03872_ ), .A4(_08533_ ), .ZN(_03873_ ) );
AND2_X1 _24636_ ( .A1(\io_master_awaddr [25] ), .A2(\io_master_awaddr [24] ), .ZN(_03874_ ) );
NAND4_X1 _24637_ ( .A1(_03873_ ), .A2(\io_master_awaddr [23] ), .A3(\io_master_awaddr [22] ), .A4(_03874_ ), .ZN(_03875_ ) );
NAND4_X1 _24638_ ( .A1(\io_master_awaddr [17] ), .A2(\io_master_awaddr [16] ), .A3(\io_master_awaddr [15] ), .A4(\io_master_awaddr [14] ), .ZN(_03876_ ) );
NAND4_X1 _24639_ ( .A1(\io_master_awaddr [21] ), .A2(\io_master_awaddr [20] ), .A3(\io_master_awaddr [19] ), .A4(\io_master_awaddr [18] ), .ZN(_03877_ ) );
NOR4_X1 _24640_ ( .A1(_03869_ ), .A2(_03875_ ), .A3(_03876_ ), .A4(_03877_ ), .ZN(_03878_ ) );
NAND2_X1 _24641_ ( .A1(\io_master_awaddr [29] ), .A2(\io_master_awaddr [28] ), .ZN(_03879_ ) );
OAI21_X1 _24642_ ( .A(_03863_ ), .B1(_03878_ ), .B2(_03879_ ), .ZN(_03880_ ) );
AND2_X1 _24643_ ( .A1(_03880_ ), .A2(_08542_ ), .ZN(_03881_ ) );
BUF_X2 _24644_ ( .A(_03881_ ), .Z(_03882_ ) );
NOR2_X1 _24645_ ( .A1(\io_master_awaddr [1] ), .A2(\io_master_awaddr [0] ), .ZN(_03883_ ) );
NOR2_X1 _24646_ ( .A1(_03882_ ), .A2(_03883_ ), .ZN(_03884_ ) );
NOR3_X1 _24647_ ( .A1(_08547_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A3(_08560_ ), .ZN(_03885_ ) );
AOI21_X1 _24648_ ( .A(_03885_ ), .B1(_08563_ ), .B2(\io_master_rdata [31] ), .ZN(_03886_ ) );
NOR2_X1 _24649_ ( .A1(_03886_ ), .A2(_10988_ ), .ZN(_03887_ ) );
INV_X1 _24650_ ( .A(_03887_ ), .ZN(_03888_ ) );
NOR3_X1 _24651_ ( .A1(_08547_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_8_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A3(_08560_ ), .ZN(_03889_ ) );
AOI21_X1 _24652_ ( .A(_03889_ ), .B1(_08563_ ), .B2(\io_master_rdata [23] ), .ZN(_03890_ ) );
NOR2_X1 _24653_ ( .A1(_03890_ ), .A2(_10988_ ), .ZN(_03891_ ) );
INV_X1 _24654_ ( .A(_03891_ ), .ZN(_03892_ ) );
OAI221_X1 _24655_ ( .A(_03884_ ), .B1(_03888_ ), .B2(\io_master_awaddr [0] ), .C1(\io_master_awaddr [1] ), .C2(_03892_ ), .ZN(_03893_ ) );
NOR3_X1 _24656_ ( .A1(_08547_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_16_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A3(_08560_ ), .ZN(_03894_ ) );
AOI21_X1 _24657_ ( .A(_03894_ ), .B1(_08563_ ), .B2(\io_master_rdata [15] ), .ZN(_03895_ ) );
OAI22_X1 _24658_ ( .A1(_03882_ ), .A2(_03883_ ), .B1(_10988_ ), .B2(_03895_ ), .ZN(_03896_ ) );
AND2_X2 _24659_ ( .A1(_03893_ ), .A2(_03896_ ), .ZN(_03897_ ) );
AND2_X1 _24660_ ( .A1(_03897_ ), .A2(\lsu.io_in_bits_lh ), .ZN(_03898_ ) );
BUF_X4 _24661_ ( .A(_03884_ ), .Z(_03899_ ) );
INV_X1 _24662_ ( .A(\arbiter.io_lsu_arsize [1] ), .ZN(_03900_ ) );
NOR3_X1 _24663_ ( .A1(_03899_ ), .A2(_03900_ ), .A3(_03888_ ), .ZN(_03901_ ) );
OR2_X1 _24664_ ( .A1(_03898_ ), .A2(_03901_ ), .ZN(_03902_ ) );
MUX2_X1 _24665_ ( .A(_03892_ ), .B(_03888_ ), .S(\io_master_awaddr [0] ), .Z(_03903_ ) );
NAND2_X1 _24666_ ( .A1(_03903_ ), .A2(\io_master_awaddr [1] ), .ZN(_03904_ ) );
INV_X1 _24667_ ( .A(\io_master_awaddr [0] ), .ZN(_03905_ ) );
NOR2_X1 _24668_ ( .A1(_03905_ ), .A2(\io_master_awaddr [1] ), .ZN(_03906_ ) );
OAI21_X1 _24669_ ( .A(_03906_ ), .B1(_03895_ ), .B2(_10988_ ), .ZN(_03907_ ) );
AOI21_X1 _24670_ ( .A(_03882_ ), .B1(_03904_ ), .B2(_03907_ ), .ZN(_03908_ ) );
INV_X1 _24671_ ( .A(_03882_ ), .ZN(_03909_ ) );
INV_X1 _24672_ ( .A(_03883_ ), .ZN(_03910_ ) );
OR3_X1 _24673_ ( .A1(_08547_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_8_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_08560_ ), .ZN(_03911_ ) );
OAI21_X1 _24674_ ( .A(\io_master_rdata [7] ), .B1(_08547_ ), .B2(_08560_ ), .ZN(_03912_ ) );
NAND2_X1 _24675_ ( .A1(_03911_ ), .A2(_03912_ ), .ZN(_03913_ ) );
AOI22_X1 _24676_ ( .A1(_03909_ ), .A2(_03910_ ), .B1(fanout_net_1 ), .B2(_03913_ ), .ZN(_03914_ ) );
NOR2_X1 _24677_ ( .A1(_03908_ ), .A2(_03914_ ), .ZN(_03915_ ) );
AND2_X1 _24678_ ( .A1(_03915_ ), .A2(\lsu.io_in_bits_lb ), .ZN(_03916_ ) );
BUF_X4 _24679_ ( .A(_03916_ ), .Z(_03917_ ) );
OAI21_X1 _24680_ ( .A(\lsu.io_in_bits_ren ), .B1(_03902_ ), .B2(_03917_ ), .ZN(_03918_ ) );
INV_X1 _24681_ ( .A(io_master_bready ), .ZN(_03919_ ) );
NOR3_X1 _24682_ ( .A1(_08564_ ), .A2(_03919_ ), .A3(_10988_ ), .ZN(_03920_ ) );
INV_X1 _24683_ ( .A(\lsu.io_in_bits_ren ), .ZN(_03921_ ) );
AND4_X1 _24684_ ( .A1(\lsu.io_in_valid ), .A2(_03921_ ), .A3(\lsu._io_in_ready_T ), .A4(\lsu.io_in_bits_wen_rd ), .ZN(_03922_ ) );
OAI211_X1 _24685_ ( .A(_10773_ ), .B(_10755_ ), .C1(_03920_ ), .C2(_03922_ ), .ZN(_03923_ ) );
NOR2_X1 _24686_ ( .A1(_08570_ ), .A2(_03923_ ), .ZN(_03924_ ) );
BUF_X2 _24687_ ( .A(_03924_ ), .Z(_03925_ ) );
BUF_X4 _24688_ ( .A(_03921_ ), .Z(_03926_ ) );
BUF_X4 _24689_ ( .A(_03926_ ), .Z(_03927_ ) );
NAND2_X1 _24690_ ( .A1(_03927_ ), .A2(\lsu.io_in_bits_rd_wdata [31] ), .ZN(_03928_ ) );
AND3_X1 _24691_ ( .A1(_03918_ ), .A2(_03925_ ), .A3(_03928_ ), .ZN(_03929_ ) );
INV_X1 _24692_ ( .A(_03924_ ), .ZN(_03930_ ) );
BUF_X4 _24693_ ( .A(_03930_ ), .Z(_03931_ ) );
BUF_X4 _24694_ ( .A(_03931_ ), .Z(_03932_ ) );
XOR2_X1 _24695_ ( .A(\idu.io_in_bits_pc [4] ), .B(\wbu.io_in_bits_pc [4] ), .Z(_03933_ ) );
XOR2_X1 _24696_ ( .A(\idu.io_in_bits_pc [16] ), .B(\wbu.io_in_bits_pc [16] ), .Z(_03934_ ) );
INV_X1 _24697_ ( .A(\idu.io_in_bits_pc [29] ), .ZN(_03935_ ) );
NAND2_X1 _24698_ ( .A1(_03935_ ), .A2(\wbu.io_in_bits_pc [29] ), .ZN(_03936_ ) );
INV_X1 _24699_ ( .A(\wbu.io_in_bits_pc [26] ), .ZN(_03937_ ) );
OAI21_X1 _24700_ ( .A(_03936_ ), .B1(\idu.io_in_bits_pc [26] ), .B2(_03937_ ), .ZN(_03938_ ) );
INV_X1 _24701_ ( .A(\wbu.io_in_bits_pc [25] ), .ZN(_03939_ ) );
OAI22_X1 _24702_ ( .A1(_03935_ ), .A2(\wbu.io_in_bits_pc [29] ), .B1(_03939_ ), .B2(\idu.io_in_bits_pc [25] ), .ZN(_03940_ ) );
NOR4_X1 _24703_ ( .A1(_03933_ ), .A2(_03934_ ), .A3(_03938_ ), .A4(_03940_ ), .ZN(_03941_ ) );
INV_X1 _24704_ ( .A(\idu.io_in_bits_pc [21] ), .ZN(_03942_ ) );
AOI22_X1 _24705_ ( .A1(\idu.io_in_bits_pc [25] ), .A2(_03939_ ), .B1(_03942_ ), .B2(\wbu.io_in_bits_pc [21] ), .ZN(_03943_ ) );
INV_X1 _24706_ ( .A(\idu.io_in_bits_pc [11] ), .ZN(_03944_ ) );
NAND2_X1 _24707_ ( .A1(_03944_ ), .A2(\wbu.io_in_bits_pc [11] ), .ZN(_03945_ ) );
OAI211_X1 _24708_ ( .A(_03943_ ), .B(_03945_ ), .C1(_03942_ ), .C2(\wbu.io_in_bits_pc [21] ), .ZN(_03946_ ) );
INV_X1 _24709_ ( .A(\idu.io_in_bits_pc [10] ), .ZN(_03947_ ) );
NOR2_X1 _24710_ ( .A1(_03947_ ), .A2(\wbu.io_in_bits_pc [10] ), .ZN(_03948_ ) );
INV_X1 _24711_ ( .A(\wbu.io_in_bits_pc [17] ), .ZN(_03949_ ) );
AND2_X1 _24712_ ( .A1(_03949_ ), .A2(\idu.io_in_bits_pc [17] ), .ZN(_03950_ ) );
OAI22_X1 _24713_ ( .A1(\idu.io_in_bits_pc [17] ), .A2(_03949_ ), .B1(_03944_ ), .B2(\wbu.io_in_bits_pc [11] ), .ZN(_03951_ ) );
NOR4_X1 _24714_ ( .A1(_03946_ ), .A2(_03948_ ), .A3(_03950_ ), .A4(_03951_ ), .ZN(_03952_ ) );
XNOR2_X1 _24715_ ( .A(\idu.io_in_bits_pc [12] ), .B(\wbu.io_in_bits_pc [12] ), .ZN(_03953_ ) );
XNOR2_X1 _24716_ ( .A(\idu.io_in_bits_pc [8] ), .B(\wbu.io_in_bits_pc [8] ), .ZN(_03954_ ) );
XNOR2_X1 _24717_ ( .A(\idu.io_in_bits_pc [1] ), .B(\wbu.io_in_bits_pc [1] ), .ZN(_03955_ ) );
XNOR2_X1 _24718_ ( .A(\idu.io_in_bits_pc [24] ), .B(\wbu.io_in_bits_pc [24] ), .ZN(_03956_ ) );
AND4_X1 _24719_ ( .A1(_03953_ ), .A2(_03954_ ), .A3(_03955_ ), .A4(_03956_ ), .ZN(_03957_ ) );
INV_X1 _24720_ ( .A(\idu.io_in_bits_pc [20] ), .ZN(_03958_ ) );
AOI22_X1 _24721_ ( .A1(\idu.io_in_bits_pc [26] ), .A2(_03937_ ), .B1(_03958_ ), .B2(\wbu.io_in_bits_pc [20] ), .ZN(_03959_ ) );
INV_X1 _24722_ ( .A(\idu.io_in_bits_pc [28] ), .ZN(_03960_ ) );
NAND2_X1 _24723_ ( .A1(_03960_ ), .A2(\wbu.io_in_bits_pc [28] ), .ZN(_03961_ ) );
OAI211_X1 _24724_ ( .A(_03959_ ), .B(_03961_ ), .C1(_03958_ ), .C2(\wbu.io_in_bits_pc [20] ), .ZN(_03962_ ) );
XOR2_X1 _24725_ ( .A(\idu.io_in_bits_pc [2] ), .B(\wbu.io_in_bits_pc [2] ), .Z(_03963_ ) );
XOR2_X1 _24726_ ( .A(\idu.io_in_bits_pc [3] ), .B(\wbu.io_in_bits_pc [3] ), .Z(_03964_ ) );
NOR3_X1 _24727_ ( .A1(_03962_ ), .A2(_03963_ ), .A3(_03964_ ), .ZN(_03965_ ) );
AND4_X1 _24728_ ( .A1(_03941_ ), .A2(_03952_ ), .A3(_03957_ ), .A4(_03965_ ), .ZN(_03966_ ) );
XNOR2_X1 _24729_ ( .A(\idu.io_in_bits_pc [6] ), .B(\wbu.io_in_bits_pc [6] ), .ZN(_03967_ ) );
XNOR2_X1 _24730_ ( .A(\idu.io_in_bits_pc [19] ), .B(\wbu.io_in_bits_pc [19] ), .ZN(_03968_ ) );
XNOR2_X1 _24731_ ( .A(\idu.io_in_bits_pc [13] ), .B(\wbu.io_in_bits_pc [13] ), .ZN(_03969_ ) );
XNOR2_X1 _24732_ ( .A(\idu.io_in_bits_pc [9] ), .B(\wbu.io_in_bits_pc [9] ), .ZN(_03970_ ) );
AND4_X1 _24733_ ( .A1(_03967_ ), .A2(_03968_ ), .A3(_03969_ ), .A4(_03970_ ), .ZN(_03971_ ) );
XNOR2_X1 _24734_ ( .A(\idu.io_in_bits_pc [23] ), .B(\wbu.io_in_bits_pc [23] ), .ZN(_03972_ ) );
NOR2_X1 _24735_ ( .A1(_03960_ ), .A2(\wbu.io_in_bits_pc [28] ), .ZN(_03973_ ) );
AOI21_X1 _24736_ ( .A(_03973_ ), .B1(_03947_ ), .B2(\wbu.io_in_bits_pc [10] ), .ZN(_03974_ ) );
XNOR2_X1 _24737_ ( .A(\idu.io_in_bits_pc [22] ), .B(\wbu.io_in_bits_pc [22] ), .ZN(_03975_ ) );
XNOR2_X1 _24738_ ( .A(\idu.io_in_bits_pc [27] ), .B(\wbu.io_in_bits_pc [27] ), .ZN(_03976_ ) );
AND4_X1 _24739_ ( .A1(_03972_ ), .A2(_03974_ ), .A3(_03975_ ), .A4(_03976_ ), .ZN(_03977_ ) );
XNOR2_X1 _24740_ ( .A(\idu.io_in_bits_pc [7] ), .B(\wbu.io_in_bits_pc [7] ), .ZN(_03978_ ) );
XNOR2_X1 _24741_ ( .A(\idu.io_in_bits_pc [18] ), .B(\wbu.io_in_bits_pc [18] ), .ZN(_03979_ ) );
XNOR2_X1 _24742_ ( .A(\idu.io_in_bits_pc [5] ), .B(\wbu.io_in_bits_pc [5] ), .ZN(_03980_ ) );
XNOR2_X1 _24743_ ( .A(\idu.io_in_bits_pc [31] ), .B(\wbu.io_in_bits_pc [31] ), .ZN(_03981_ ) );
AND4_X1 _24744_ ( .A1(_03978_ ), .A2(_03979_ ), .A3(_03980_ ), .A4(_03981_ ), .ZN(_03982_ ) );
XNOR2_X1 _24745_ ( .A(\idu.io_in_bits_pc [15] ), .B(\wbu.io_in_bits_pc [15] ), .ZN(_03983_ ) );
XNOR2_X1 _24746_ ( .A(\idu.io_in_bits_pc [30] ), .B(\wbu.io_in_bits_pc [30] ), .ZN(_03984_ ) );
XNOR2_X1 _24747_ ( .A(\idu.io_in_bits_pc [0] ), .B(\wbu.io_in_bits_pc [0] ), .ZN(_03985_ ) );
XNOR2_X1 _24748_ ( .A(\idu.io_in_bits_pc [14] ), .B(\wbu.io_in_bits_pc [14] ), .ZN(_03986_ ) );
AND4_X1 _24749_ ( .A1(_03983_ ), .A2(_03984_ ), .A3(_03985_ ), .A4(_03986_ ), .ZN(_03987_ ) );
AND4_X1 _24750_ ( .A1(_03971_ ), .A2(_03977_ ), .A3(_03982_ ), .A4(_03987_ ), .ZN(_03988_ ) );
AND2_X2 _24751_ ( .A1(_03966_ ), .A2(_03988_ ), .ZN(_03989_ ) );
INV_X1 _24752_ ( .A(_03989_ ), .ZN(_03990_ ) );
BUF_X4 _24753_ ( .A(_03990_ ), .Z(_03991_ ) );
BUF_X2 _24754_ ( .A(_10767_ ), .Z(_03992_ ) );
BUF_X2 _24755_ ( .A(_03992_ ), .Z(_03993_ ) );
BUF_X2 _24756_ ( .A(_03993_ ), .Z(_03994_ ) );
XNOR2_X1 _24757_ ( .A(_03994_ ), .B(_08571_ ), .ZN(_03995_ ) );
AOI21_X1 _24758_ ( .A(_12978_ ), .B1(_11030_ ), .B2(\idu.io_in_bits_inst [18] ), .ZN(_03996_ ) );
NOR4_X1 _24759_ ( .A1(_13276_ ), .A2(_03995_ ), .A3(wbu_io_in_valid_REG_$_NOT__A_Y ), .A4(_03996_ ), .ZN(_03997_ ) );
BUF_X4 _24760_ ( .A(_03997_ ), .Z(_03998_ ) );
NAND3_X1 _24761_ ( .A1(_11030_ ), .A2(\idu.io_in_bits_inst [16] ), .A3(_08576_ ), .ZN(_03999_ ) );
BUF_X2 _24762_ ( .A(_10593_ ), .Z(_04000_ ) );
OAI21_X1 _24763_ ( .A(\wbu.io_in_bits_rd [1] ), .B1(_10760_ ), .B2(_04000_ ), .ZN(_04001_ ) );
NAND3_X1 _24764_ ( .A1(_11030_ ), .A2(\idu.io_in_bits_inst [15] ), .A3(_12972_ ), .ZN(_04002_ ) );
BUF_X4 _24765_ ( .A(_11030_ ), .Z(_04003_ ) );
NAND3_X1 _24766_ ( .A1(_04003_ ), .A2(\idu.io_in_bits_inst [18] ), .A3(_12978_ ), .ZN(_04004_ ) );
BUF_X4 _24767_ ( .A(_10628_ ), .Z(_04005_ ) );
OAI21_X1 _24768_ ( .A(\wbu.io_in_bits_rd [0] ), .B1(_10760_ ), .B2(_04005_ ), .ZN(_04006_ ) );
AND4_X1 _24769_ ( .A1(_04001_ ), .A2(_04002_ ), .A3(_04004_ ), .A4(_04006_ ), .ZN(_04007_ ) );
NAND3_X1 _24770_ ( .A1(_04003_ ), .A2(\idu.io_in_bits_inst [17] ), .A3(_13006_ ), .ZN(_04008_ ) );
OAI21_X1 _24771_ ( .A(\wbu.io_in_bits_rd [2] ), .B1(_11082_ ), .B2(_10596_ ), .ZN(_04009_ ) );
AND4_X2 _24772_ ( .A1(_03999_ ), .A2(_04007_ ), .A3(_04008_ ), .A4(_04009_ ), .ZN(_04010_ ) );
BUF_X4 _24773_ ( .A(_04010_ ), .Z(_04011_ ) );
NAND4_X1 _24774_ ( .A1(_03991_ ), .A2(\wbu.io_in_bits_rd_wdata [31] ), .A3(_03998_ ), .A4(_04011_ ), .ZN(_04012_ ) );
AOI211_X1 _24775_ ( .A(_03859_ ), .B(_03929_ ), .C1(_03932_ ), .C2(_04012_ ), .ZN(_04013_ ) );
OAI21_X1 _24776_ ( .A(_03850_ ), .B1(_03858_ ), .B2(_04013_ ), .ZN(_04014_ ) );
BUF_X4 _24777_ ( .A(_10595_ ), .Z(_04015_ ) );
BUF_X2 _24778_ ( .A(_10767_ ), .Z(_04016_ ) );
CLKBUF_X2 _24779_ ( .A(_04016_ ), .Z(_04017_ ) );
BUF_X2 _24780_ ( .A(_04017_ ), .Z(_04018_ ) );
BUF_X2 _24781_ ( .A(_04018_ ), .Z(_04019_ ) );
BUF_X2 _24782_ ( .A(_04019_ ), .Z(_04020_ ) );
AND3_X1 _24783_ ( .A1(_04020_ ), .A2(_10600_ ), .A3(\idu.io_in_bits_inst [17] ), .ZN(_04021_ ) );
INV_X1 _24784_ ( .A(_04021_ ), .ZN(_04022_ ) );
BUF_X4 _24785_ ( .A(_04022_ ), .Z(_04023_ ) );
AOI211_X1 _24786_ ( .A(_04015_ ), .B(_04023_ ), .C1(_04005_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04024_ ) );
NOR2_X1 _24787_ ( .A1(_10792_ ), .A2(_10629_ ), .ZN(_04025_ ) );
BUF_X2 _24788_ ( .A(_04025_ ), .Z(_04026_ ) );
AND2_X2 _24789_ ( .A1(_04026_ ), .A2(_04016_ ), .ZN(_04027_ ) );
INV_X1 _24790_ ( .A(_04027_ ), .ZN(_04028_ ) );
BUF_X2 _24791_ ( .A(_04028_ ), .Z(_04029_ ) );
CLKBUF_X2 _24792_ ( .A(_04029_ ), .Z(_04030_ ) );
AND2_X1 _24793_ ( .A1(_10597_ ), .A2(\idu.io_in_bits_inst [18] ), .ZN(_04031_ ) );
BUF_X2 _24794_ ( .A(_04031_ ), .Z(_04032_ ) );
INV_X1 _24795_ ( .A(_04032_ ), .ZN(_04033_ ) );
BUF_X2 _24796_ ( .A(_04033_ ), .Z(_04034_ ) );
NOR3_X1 _24797_ ( .A1(_04030_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04034_ ), .ZN(_04035_ ) );
BUF_X2 _24798_ ( .A(_04032_ ), .Z(_04036_ ) );
BUF_X2 _24799_ ( .A(_04026_ ), .Z(_04037_ ) );
BUF_X2 _24800_ ( .A(_04037_ ), .Z(_04038_ ) );
BUF_X2 _24801_ ( .A(_11098_ ), .Z(_04039_ ) );
BUF_X2 _24802_ ( .A(_04039_ ), .Z(_04040_ ) );
BUF_X4 _24803_ ( .A(_04040_ ), .Z(_04041_ ) );
BUF_X4 _24804_ ( .A(_04041_ ), .Z(_04042_ ) );
BUF_X2 _24805_ ( .A(_04042_ ), .Z(_04043_ ) );
NAND4_X1 _24806_ ( .A1(_04036_ ), .A2(_04038_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04043_ ), .ZN(_04044_ ) );
AND2_X2 _24807_ ( .A1(_10600_ ), .A2(_10596_ ), .ZN(_04045_ ) );
AND2_X2 _24808_ ( .A1(_10594_ ), .A2(_10628_ ), .ZN(_04046_ ) );
AND2_X1 _24809_ ( .A1(_04045_ ), .A2(_04046_ ), .ZN(_04047_ ) );
BUF_X2 _24810_ ( .A(_04047_ ), .Z(_04048_ ) );
NAND3_X1 _24811_ ( .A1(_04048_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04042_ ), .ZN(_04049_ ) );
NOR2_X1 _24812_ ( .A1(_10597_ ), .A2(_10600_ ), .ZN(_04050_ ) );
AND2_X2 _24813_ ( .A1(_04046_ ), .A2(_04050_ ), .ZN(_04051_ ) );
AND2_X1 _24814_ ( .A1(_04051_ ), .A2(_11096_ ), .ZN(_04052_ ) );
BUF_X4 _24815_ ( .A(_04052_ ), .Z(_04053_ ) );
INV_X1 _24816_ ( .A(_04053_ ), .ZN(_04054_ ) );
NOR2_X1 _24817_ ( .A1(_04054_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04055_ ) );
INV_X1 _24818_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_04056_ ) );
AND2_X2 _24819_ ( .A1(_10629_ ), .A2(_10593_ ), .ZN(_04057_ ) );
AND2_X1 _24820_ ( .A1(_04057_ ), .A2(_04050_ ), .ZN(_04058_ ) );
AND2_X1 _24821_ ( .A1(_04058_ ), .A2(_11096_ ), .ZN(_04059_ ) );
AOI21_X1 _24822_ ( .A(_04055_ ), .B1(_04056_ ), .B2(_04059_ ), .ZN(_04060_ ) );
AND2_X1 _24823_ ( .A1(_10629_ ), .A2(\idu.io_in_bits_inst [16] ), .ZN(_04061_ ) );
AND2_X1 _24824_ ( .A1(_04061_ ), .A2(_04050_ ), .ZN(_04062_ ) );
AND2_X1 _24825_ ( .A1(_04062_ ), .A2(_11096_ ), .ZN(_04063_ ) );
INV_X1 _24826_ ( .A(_04063_ ), .ZN(_04064_ ) );
OAI21_X1 _24827_ ( .A(_04060_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04064_ ), .ZN(_04065_ ) );
AND2_X2 _24828_ ( .A1(_10597_ ), .A2(_10599_ ), .ZN(_04066_ ) );
AND2_X1 _24829_ ( .A1(_04066_ ), .A2(_04025_ ), .ZN(_04067_ ) );
AND2_X2 _24830_ ( .A1(_04067_ ), .A2(_11096_ ), .ZN(_04068_ ) );
INV_X1 _24831_ ( .A(_04068_ ), .ZN(_04069_ ) );
BUF_X2 _24832_ ( .A(_04069_ ), .Z(_04070_ ) );
NOR2_X1 _24833_ ( .A1(_04070_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04071_ ) );
INV_X1 _24834_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04072_ ) );
BUF_X2 _24835_ ( .A(_04057_ ), .Z(_04073_ ) );
BUF_X2 _24836_ ( .A(_04066_ ), .Z(_04074_ ) );
AND4_X1 _24837_ ( .A1(_04072_ ), .A2(_04073_ ), .A3(_04074_ ), .A4(_04039_ ), .ZN(_04075_ ) );
NOR3_X1 _24838_ ( .A1(_04065_ ), .A2(_04071_ ), .A3(_04075_ ), .ZN(_04076_ ) );
AND2_X2 _24839_ ( .A1(_04066_ ), .A2(_04046_ ), .ZN(_04077_ ) );
BUF_X2 _24840_ ( .A(_04077_ ), .Z(_04078_ ) );
INV_X1 _24841_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04079_ ) );
BUF_X2 _24842_ ( .A(_11099_ ), .Z(_04080_ ) );
NAND3_X1 _24843_ ( .A1(_04078_ ), .A2(_04079_ ), .A3(_04080_ ), .ZN(_04081_ ) );
AND2_X1 _24844_ ( .A1(_04061_ ), .A2(_04066_ ), .ZN(_04082_ ) );
AND2_X1 _24845_ ( .A1(_04082_ ), .A2(_11097_ ), .ZN(_04083_ ) );
INV_X1 _24846_ ( .A(_04083_ ), .ZN(_04084_ ) );
BUF_X2 _24847_ ( .A(_04084_ ), .Z(_04085_ ) );
OR2_X1 _24848_ ( .A1(_04085_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04086_ ) );
AND3_X1 _24849_ ( .A1(_04076_ ), .A2(_04081_ ), .A3(_04086_ ), .ZN(_04087_ ) );
AND3_X1 _24850_ ( .A1(_10600_ ), .A2(_10596_ ), .A3(_10604_ ), .ZN(_04088_ ) );
AND2_X1 _24851_ ( .A1(_04088_ ), .A2(_04025_ ), .ZN(_04089_ ) );
INV_X1 _24852_ ( .A(_04089_ ), .ZN(_04090_ ) );
OAI21_X1 _24853_ ( .A(_04087_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04090_ ), .ZN(_04091_ ) );
AND2_X1 _24854_ ( .A1(_04088_ ), .A2(_04057_ ), .ZN(_04092_ ) );
INV_X1 _24855_ ( .A(_04092_ ), .ZN(_04093_ ) );
INV_X1 _24856_ ( .A(_04047_ ), .ZN(_04094_ ) );
BUF_X2 _24857_ ( .A(_04094_ ), .Z(_04095_ ) );
OAI22_X1 _24858_ ( .A1(_04093_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_04095_ ), .B2(_03994_ ), .ZN(_04096_ ) );
OAI21_X1 _24859_ ( .A(_04049_ ), .B1(_04091_ ), .B2(_04096_ ), .ZN(_04097_ ) );
CLKBUF_X2 _24860_ ( .A(_04061_ ), .Z(_04098_ ) );
AND2_X1 _24861_ ( .A1(_04045_ ), .A2(_04098_ ), .ZN(_04099_ ) );
AND2_X1 _24862_ ( .A1(_04099_ ), .A2(_11099_ ), .ZN(_04100_ ) );
INV_X1 _24863_ ( .A(_04100_ ), .ZN(_04101_ ) );
BUF_X2 _24864_ ( .A(_04101_ ), .Z(_04102_ ) );
OAI21_X1 _24865_ ( .A(_04097_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04102_ ), .ZN(_04103_ ) );
AND2_X2 _24866_ ( .A1(_04031_ ), .A2(_10604_ ), .ZN(_04104_ ) );
AND2_X1 _24867_ ( .A1(_04104_ ), .A2(_04025_ ), .ZN(_04105_ ) );
OAI21_X1 _24868_ ( .A(_04044_ ), .B1(_04103_ ), .B2(_04105_ ), .ZN(_04106_ ) );
BUF_X2 _24869_ ( .A(_04073_ ), .Z(_04107_ ) );
BUF_X2 _24870_ ( .A(_04107_ ), .Z(_04108_ ) );
BUF_X2 _24871_ ( .A(_04108_ ), .Z(_04109_ ) );
CLKBUF_X2 _24872_ ( .A(_04031_ ), .Z(_04110_ ) );
BUF_X2 _24873_ ( .A(_04110_ ), .Z(_04111_ ) );
INV_X1 _24874_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04112_ ) );
BUF_X4 _24875_ ( .A(_04042_ ), .Z(_04113_ ) );
BUF_X4 _24876_ ( .A(_04113_ ), .Z(_04114_ ) );
NAND4_X1 _24877_ ( .A1(_04109_ ), .A2(_04111_ ), .A3(_04112_ ), .A4(_04114_ ), .ZN(_04115_ ) );
BUF_X2 _24878_ ( .A(_04046_ ), .Z(_04116_ ) );
BUF_X2 _24879_ ( .A(_04116_ ), .Z(_04117_ ) );
BUF_X2 _24880_ ( .A(_04117_ ), .Z(_04118_ ) );
BUF_X2 _24881_ ( .A(_04118_ ), .Z(_04119_ ) );
INV_X1 _24882_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04120_ ) );
NAND4_X1 _24883_ ( .A1(_04119_ ), .A2(_04111_ ), .A3(_04120_ ), .A4(_04114_ ), .ZN(_04121_ ) );
NAND3_X1 _24884_ ( .A1(_04106_ ), .A2(_04115_ ), .A3(_04121_ ), .ZN(_04122_ ) );
INV_X1 _24885_ ( .A(_04061_ ), .ZN(_04123_ ) );
CLKBUF_X2 _24886_ ( .A(_04123_ ), .Z(_04124_ ) );
BUF_X2 _24887_ ( .A(_04124_ ), .Z(_04125_ ) );
BUF_X2 _24888_ ( .A(_04125_ ), .Z(_04126_ ) );
BUF_X2 _24889_ ( .A(_03992_ ), .Z(_04127_ ) );
CLKBUF_X2 _24890_ ( .A(_04127_ ), .Z(_04128_ ) );
BUF_X2 _24891_ ( .A(_04128_ ), .Z(_04129_ ) );
NOR4_X1 _24892_ ( .A1(_04126_ ), .A2(_04034_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04129_ ), .ZN(_04130_ ) );
BUF_X2 _24893_ ( .A(_04028_ ), .Z(_04131_ ) );
NOR4_X1 _24894_ ( .A1(_04131_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10597_ ), .A4(_10600_ ), .ZN(_04132_ ) );
NOR3_X1 _24895_ ( .A1(_04122_ ), .A2(_04130_ ), .A3(_04132_ ), .ZN(_04133_ ) );
BUF_X2 _24896_ ( .A(_04058_ ), .Z(_04134_ ) );
AND2_X1 _24897_ ( .A1(_04134_ ), .A2(_04018_ ), .ZN(_04135_ ) );
INV_X1 _24898_ ( .A(_04135_ ), .ZN(_04136_ ) );
OR2_X1 _24899_ ( .A1(_04136_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04137_ ) );
BUF_X2 _24900_ ( .A(_04127_ ), .Z(_04138_ ) );
AND2_X1 _24901_ ( .A1(_04051_ ), .A2(_04138_ ), .ZN(_04139_ ) );
INV_X1 _24902_ ( .A(_04139_ ), .ZN(_04140_ ) );
OR2_X1 _24903_ ( .A1(_04140_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04141_ ) );
NAND3_X1 _24904_ ( .A1(_04133_ ), .A2(_04137_ ), .A3(_04141_ ), .ZN(_04142_ ) );
INV_X1 _24905_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04143_ ) );
BUF_X2 _24906_ ( .A(_04098_ ), .Z(_04144_ ) );
BUF_X2 _24907_ ( .A(_04144_ ), .Z(_04145_ ) );
BUF_X2 _24908_ ( .A(_04145_ ), .Z(_04146_ ) );
BUF_X2 _24909_ ( .A(_04146_ ), .Z(_04147_ ) );
BUF_X2 _24910_ ( .A(_04050_ ), .Z(_04148_ ) );
BUF_X2 _24911_ ( .A(_04148_ ), .Z(_04149_ ) );
BUF_X2 _24912_ ( .A(_04149_ ), .Z(_04150_ ) );
BUF_X2 _24913_ ( .A(_04150_ ), .Z(_04151_ ) );
AND4_X1 _24914_ ( .A1(_04143_ ), .A2(_04147_ ), .A3(_04151_ ), .A4(_04020_ ), .ZN(_04152_ ) );
INV_X1 _24915_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04153_ ) );
BUF_X2 _24916_ ( .A(_04074_ ), .Z(_04154_ ) );
BUF_X2 _24917_ ( .A(_04154_ ), .Z(_04155_ ) );
BUF_X2 _24918_ ( .A(_04155_ ), .Z(_04156_ ) );
BUF_X2 _24919_ ( .A(_04038_ ), .Z(_04157_ ) );
CLKBUF_X2 _24920_ ( .A(_04157_ ), .Z(_04158_ ) );
CLKBUF_X2 _24921_ ( .A(_04129_ ), .Z(_04159_ ) );
AND4_X1 _24922_ ( .A1(_04153_ ), .A2(_04156_ ), .A3(_04158_ ), .A4(_04159_ ), .ZN(_04160_ ) );
NOR3_X1 _24923_ ( .A1(_04142_ ), .A2(_04152_ ), .A3(_04160_ ), .ZN(_04161_ ) );
AND2_X2 _24924_ ( .A1(_04057_ ), .A2(_04066_ ), .ZN(_04162_ ) );
BUF_X2 _24925_ ( .A(_04138_ ), .Z(_04163_ ) );
AND2_X1 _24926_ ( .A1(_04162_ ), .A2(_04163_ ), .ZN(_04164_ ) );
INV_X1 _24927_ ( .A(_04164_ ), .ZN(_04165_ ) );
OR2_X1 _24928_ ( .A1(_04165_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04166_ ) );
BUF_X2 _24929_ ( .A(_04156_ ), .Z(_04167_ ) );
BUF_X4 _24930_ ( .A(_04167_ ), .Z(_04168_ ) );
BUF_X2 _24931_ ( .A(_04117_ ), .Z(_04169_ ) );
BUF_X2 _24932_ ( .A(_04169_ ), .Z(_04170_ ) );
BUF_X2 _24933_ ( .A(_04170_ ), .Z(_04171_ ) );
INV_X1 _24934_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04172_ ) );
BUF_X2 _24935_ ( .A(_04163_ ), .Z(_04173_ ) );
BUF_X2 _24936_ ( .A(_04173_ ), .Z(_04174_ ) );
BUF_X2 _24937_ ( .A(_04174_ ), .Z(_04175_ ) );
NAND4_X1 _24938_ ( .A1(_04168_ ), .A2(_04171_ ), .A3(_04172_ ), .A4(_04175_ ), .ZN(_04176_ ) );
NAND3_X1 _24939_ ( .A1(_04161_ ), .A2(_04166_ ), .A3(_04176_ ), .ZN(_04177_ ) );
BUF_X2 _24940_ ( .A(_04126_ ), .Z(_04178_ ) );
BUF_X2 _24941_ ( .A(_04178_ ), .Z(_04179_ ) );
INV_X1 _24942_ ( .A(_04074_ ), .ZN(_04180_ ) );
BUF_X2 _24943_ ( .A(_04180_ ), .Z(_04181_ ) );
CLKBUF_X2 _24944_ ( .A(_04181_ ), .Z(_04182_ ) );
BUF_X2 _24945_ ( .A(_04114_ ), .Z(_04183_ ) );
CLKBUF_X2 _24946_ ( .A(_04183_ ), .Z(_04184_ ) );
NOR4_X1 _24947_ ( .A1(_04179_ ), .A2(_04182_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04184_ ), .ZN(_04185_ ) );
NAND2_X2 _24948_ ( .A1(_04045_ ), .A2(_04025_ ), .ZN(_04186_ ) );
BUF_X2 _24949_ ( .A(_04186_ ), .Z(_04187_ ) );
CLKBUF_X2 _24950_ ( .A(_04187_ ), .Z(_04188_ ) );
BUF_X2 _24951_ ( .A(_04113_ ), .Z(_04189_ ) );
BUF_X2 _24952_ ( .A(_04189_ ), .Z(_04190_ ) );
CLKBUF_X2 _24953_ ( .A(_04190_ ), .Z(_04191_ ) );
NOR3_X1 _24954_ ( .A1(_04188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04191_ ), .ZN(_04192_ ) );
OR3_X1 _24955_ ( .A1(_04177_ ), .A2(_04185_ ), .A3(_04192_ ), .ZN(_04193_ ) );
BUF_X4 _24956_ ( .A(_04000_ ), .Z(_04194_ ) );
NOR4_X1 _24957_ ( .A1(_11082_ ), .A2(_10599_ ), .A3(\idu.io_in_bits_inst [17] ), .A4(_10604_ ), .ZN(_04195_ ) );
BUF_X2 _24958_ ( .A(_04195_ ), .Z(_04196_ ) );
BUF_X4 _24959_ ( .A(_04196_ ), .Z(_04197_ ) );
INV_X1 _24960_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04198_ ) );
BUF_X4 _24961_ ( .A(_10756_ ), .Z(_04199_ ) );
AND4_X1 _24962_ ( .A1(_04194_ ), .A2(_04197_ ), .A3(_04198_ ), .A4(_04199_ ), .ZN(_04200_ ) );
AND2_X1 _24963_ ( .A1(_04099_ ), .A2(_04020_ ), .ZN(_04201_ ) );
INV_X1 _24964_ ( .A(_04201_ ), .ZN(_04202_ ) );
AND2_X1 _24965_ ( .A1(_04048_ ), .A2(_04159_ ), .ZN(_04203_ ) );
INV_X1 _24966_ ( .A(_04203_ ), .ZN(_04204_ ) );
OAI21_X1 _24967_ ( .A(_04202_ ), .B1(_04204_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04205_ ) );
OR3_X1 _24968_ ( .A1(_04193_ ), .A2(_04200_ ), .A3(_04205_ ), .ZN(_04206_ ) );
BUF_X2 _24969_ ( .A(_04099_ ), .Z(_04207_ ) );
BUF_X2 _24970_ ( .A(_04173_ ), .Z(_04208_ ) );
BUF_X4 _24971_ ( .A(_04208_ ), .Z(_04209_ ) );
BUF_X4 _24972_ ( .A(_04209_ ), .Z(_04210_ ) );
BUF_X4 _24973_ ( .A(_04210_ ), .Z(_04211_ ) );
BUF_X4 _24974_ ( .A(_04211_ ), .Z(_04212_ ) );
NAND3_X1 _24975_ ( .A1(_04207_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04212_ ), .ZN(_04213_ ) );
AOI21_X1 _24976_ ( .A(_04035_ ), .B1(_04206_ ), .B2(_04213_ ), .ZN(_04214_ ) );
BUF_X2 _24977_ ( .A(_04021_ ), .Z(_04215_ ) );
CLKBUF_X2 _24978_ ( .A(_04109_ ), .Z(_04216_ ) );
BUF_X2 _24979_ ( .A(_04216_ ), .Z(_04217_ ) );
AND2_X1 _24980_ ( .A1(_04215_ ), .A2(_04217_ ), .ZN(_04218_ ) );
INV_X1 _24981_ ( .A(_04218_ ), .ZN(_04219_ ) );
NAND2_X1 _24982_ ( .A1(_04214_ ), .A2(_04219_ ), .ZN(_04220_ ) );
BUF_X4 _24983_ ( .A(_04215_ ), .Z(_04221_ ) );
BUF_X4 _24984_ ( .A(_04221_ ), .Z(_04222_ ) );
BUF_X2 _24985_ ( .A(_04217_ ), .Z(_04223_ ) );
BUF_X2 _24986_ ( .A(_04223_ ), .Z(_04224_ ) );
NAND3_X1 _24987_ ( .A1(_04222_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04224_ ), .ZN(_04225_ ) );
AOI21_X1 _24988_ ( .A(_04024_ ), .B1(_04220_ ), .B2(_04225_ ), .ZN(_04226_ ) );
NAND4_X1 _24989_ ( .A1(_10793_ ), .A2(_10798_ ), .A3(_10804_ ), .A4(_03852_ ), .ZN(_04227_ ) );
NOR2_X2 _24990_ ( .A1(_04227_ ), .A2(_10816_ ), .ZN(_04228_ ) );
INV_X1 _24991_ ( .A(_04228_ ), .ZN(_04229_ ) );
OAI21_X1 _24992_ ( .A(_04229_ ), .B1(_08570_ ), .B2(_03923_ ), .ZN(_04230_ ) );
INV_X1 _24993_ ( .A(_03996_ ), .ZN(_04231_ ) );
NAND4_X1 _24994_ ( .A1(_04231_ ), .A2(_04008_ ), .A3(_04009_ ), .A4(_04004_ ), .ZN(_04232_ ) );
NAND4_X1 _24995_ ( .A1(_03999_ ), .A2(_04002_ ), .A3(_04001_ ), .A4(_04006_ ), .ZN(_04233_ ) );
NOR3_X1 _24996_ ( .A1(_04232_ ), .A2(_04233_ ), .A3(_03995_ ), .ZN(_04234_ ) );
INV_X1 _24997_ ( .A(wbu_io_in_valid_REG_$_NOT__A_Y ), .ZN(_04235_ ) );
NAND4_X1 _24998_ ( .A1(_04234_ ), .A2(_04235_ ), .A3(_12962_ ), .A4(_12963_ ), .ZN(_04236_ ) );
NOR2_X1 _24999_ ( .A1(_03989_ ), .A2(_04236_ ), .ZN(_04237_ ) );
OR2_X1 _25000_ ( .A1(_04230_ ), .A2(_04237_ ), .ZN(_04238_ ) );
AND2_X1 _25001_ ( .A1(_04238_ ), .A2(_10574_ ), .ZN(_04239_ ) );
BUF_X2 _25002_ ( .A(_04239_ ), .Z(_04240_ ) );
BUF_X2 _25003_ ( .A(_04147_ ), .Z(_04241_ ) );
BUF_X2 _25004_ ( .A(_04241_ ), .Z(_04242_ ) );
BUF_X4 _25005_ ( .A(_04242_ ), .Z(_04243_ ) );
AND3_X1 _25006_ ( .A1(_04221_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04243_ ), .ZN(_04244_ ) );
OR2_X1 _25007_ ( .A1(_04240_ ), .A2(_04244_ ), .ZN(_04245_ ) );
OAI21_X1 _25008_ ( .A(_04014_ ), .B1(_04226_ ), .B2(_04245_ ), .ZN(\idu.io_out_bits_rs1_data [31] ) );
INV_X1 _25009_ ( .A(_04240_ ), .ZN(_04246_ ) );
BUF_X4 _25010_ ( .A(_04246_ ), .Z(_04247_ ) );
INV_X1 _25011_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_04248_ ) );
AND2_X1 _25012_ ( .A1(_04021_ ), .A2(_04241_ ), .ZN(_04249_ ) );
BUF_X4 _25013_ ( .A(_04249_ ), .Z(_04250_ ) );
INV_X1 _25014_ ( .A(_04250_ ), .ZN(_04251_ ) );
AND3_X1 _25015_ ( .A1(_04027_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04167_ ), .ZN(_04252_ ) );
BUF_X2 _25016_ ( .A(_04150_ ), .Z(_04253_ ) );
BUF_X2 _25017_ ( .A(_04129_ ), .Z(_04254_ ) );
NAND4_X1 _25018_ ( .A1(_04253_ ), .A2(_04157_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04254_ ), .ZN(_04255_ ) );
OR4_X1 _25019_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04125_ ), .A3(_04033_ ), .A4(_04018_ ), .ZN(_04256_ ) );
BUF_X2 _25020_ ( .A(_04088_ ), .Z(_04257_ ) );
INV_X1 _25021_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04258_ ) );
NAND3_X1 _25022_ ( .A1(_04257_ ), .A2(_04258_ ), .A3(_04108_ ), .ZN(_04259_ ) );
INV_X1 _25023_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04260_ ) );
AND4_X1 _25024_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04046_ ), .A3(_04050_ ), .A4(_11097_ ), .ZN(_04261_ ) );
NAND2_X1 _25025_ ( .A1(_04057_ ), .A2(_04050_ ), .ZN(_04262_ ) );
CLKBUF_X2 _25026_ ( .A(_04262_ ), .Z(_04263_ ) );
OR3_X1 _25027_ ( .A1(_04263_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10766_ ), .ZN(_04264_ ) );
AOI21_X1 _25028_ ( .A(_04261_ ), .B1(_04054_ ), .B2(_04264_ ), .ZN(_04265_ ) );
MUX2_X1 _25029_ ( .A(_04260_ ), .B(_04265_ ), .S(_04064_ ), .Z(_04266_ ) );
NOR2_X1 _25030_ ( .A1(_04070_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04267_ ) );
INV_X1 _25031_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04268_ ) );
AND4_X1 _25032_ ( .A1(_04268_ ), .A2(_04057_ ), .A3(_04074_ ), .A4(_04039_ ), .ZN(_04269_ ) );
OR3_X1 _25033_ ( .A1(_04266_ ), .A2(_04267_ ), .A3(_04269_ ), .ZN(_04270_ ) );
AND2_X1 _25034_ ( .A1(_04077_ ), .A2(_11097_ ), .ZN(_04271_ ) );
INV_X1 _25035_ ( .A(_04271_ ), .ZN(_04272_ ) );
NOR2_X1 _25036_ ( .A1(_04272_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04273_ ) );
OAI21_X1 _25037_ ( .A(_04090_ ), .B1(_04085_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04274_ ) );
NOR3_X1 _25038_ ( .A1(_04270_ ), .A2(_04273_ ), .A3(_04274_ ), .ZN(_04275_ ) );
AND3_X1 _25039_ ( .A1(_04257_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04026_ ), .ZN(_04276_ ) );
OAI21_X1 _25040_ ( .A(_04259_ ), .B1(_04275_ ), .B2(_04276_ ), .ZN(_04277_ ) );
NOR3_X1 _25041_ ( .A1(_04095_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04138_ ), .ZN(_04278_ ) );
NOR2_X1 _25042_ ( .A1(_04102_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04279_ ) );
NOR3_X1 _25043_ ( .A1(_04277_ ), .A2(_04278_ ), .A3(_04279_ ), .ZN(_04280_ ) );
INV_X1 _25044_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04281_ ) );
BUF_X2 _25045_ ( .A(_04080_ ), .Z(_04282_ ) );
BUF_X2 _25046_ ( .A(_04282_ ), .Z(_04283_ ) );
NAND4_X1 _25047_ ( .A1(_04036_ ), .A2(_04038_ ), .A3(_04281_ ), .A4(_04283_ ), .ZN(_04284_ ) );
AND2_X1 _25048_ ( .A1(_04104_ ), .A2(_04073_ ), .ZN(_04285_ ) );
INV_X1 _25049_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04286_ ) );
BUF_X2 _25050_ ( .A(_04104_ ), .Z(_04287_ ) );
AOI22_X1 _25051_ ( .A1(_04285_ ), .A2(_04286_ ), .B1(_04118_ ), .B2(_04287_ ), .ZN(_04288_ ) );
AND3_X1 _25052_ ( .A1(_04280_ ), .A2(_04284_ ), .A3(_04288_ ), .ZN(_04289_ ) );
AND3_X1 _25053_ ( .A1(_04287_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04169_ ), .ZN(_04290_ ) );
OAI21_X1 _25054_ ( .A(_04256_ ), .B1(_04289_ ), .B2(_04290_ ), .ZN(_04291_ ) );
AND2_X2 _25055_ ( .A1(_04027_ ), .A2(_04149_ ), .ZN(_04292_ ) );
OAI21_X1 _25056_ ( .A(_04255_ ), .B1(_04291_ ), .B2(_04292_ ), .ZN(_04293_ ) );
BUF_X2 _25057_ ( .A(_04263_ ), .Z(_04294_ ) );
BUF_X2 _25058_ ( .A(_04043_ ), .Z(_04295_ ) );
OR3_X1 _25059_ ( .A1(_04294_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04295_ ), .ZN(_04296_ ) );
BUF_X2 _25060_ ( .A(_04119_ ), .Z(_04297_ ) );
INV_X1 _25061_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04298_ ) );
NAND4_X1 _25062_ ( .A1(_04297_ ), .A2(_04151_ ), .A3(_04298_ ), .A4(_04174_ ), .ZN(_04299_ ) );
AND3_X1 _25063_ ( .A1(_04293_ ), .A2(_04296_ ), .A3(_04299_ ), .ZN(_04300_ ) );
AND2_X1 _25064_ ( .A1(_04062_ ), .A2(_04128_ ), .ZN(_04301_ ) );
INV_X1 _25065_ ( .A(_04301_ ), .ZN(_04302_ ) );
BUF_X2 _25066_ ( .A(_04302_ ), .Z(_04303_ ) );
NOR2_X1 _25067_ ( .A1(_04303_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04304_ ) );
AND2_X1 _25068_ ( .A1(_04027_ ), .A2(_04155_ ), .ZN(_04305_ ) );
NOR2_X1 _25069_ ( .A1(_04304_ ), .A2(_04305_ ), .ZN(_04306_ ) );
AOI21_X1 _25070_ ( .A(_04252_ ), .B1(_04300_ ), .B2(_04306_ ), .ZN(_04307_ ) );
INV_X1 _25071_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04308_ ) );
CLKBUF_X2 _25072_ ( .A(_04156_ ), .Z(_04309_ ) );
CLKBUF_X2 _25073_ ( .A(_04254_ ), .Z(_04310_ ) );
AND4_X1 _25074_ ( .A1(_04308_ ), .A2(_04216_ ), .A3(_04309_ ), .A4(_04310_ ), .ZN(_04311_ ) );
INV_X1 _25075_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04312_ ) );
BUF_X2 _25076_ ( .A(_04020_ ), .Z(_04313_ ) );
AND3_X1 _25077_ ( .A1(_04078_ ), .A2(_04312_ ), .A3(_04313_ ), .ZN(_04314_ ) );
NOR3_X1 _25078_ ( .A1(_04307_ ), .A2(_04311_ ), .A3(_04314_ ), .ZN(_04315_ ) );
CLKBUF_X2 _25079_ ( .A(_04126_ ), .Z(_04316_ ) );
BUF_X2 _25080_ ( .A(_04181_ ), .Z(_04317_ ) );
CLKBUF_X2 _25081_ ( .A(_04295_ ), .Z(_04318_ ) );
OR4_X1 _25082_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04316_ ), .A3(_04317_ ), .A4(_04318_ ), .ZN(_04319_ ) );
BUF_X2 _25083_ ( .A(_04190_ ), .Z(_04320_ ) );
OR3_X1 _25084_ ( .A1(_04188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04320_ ), .ZN(_04321_ ) );
AND3_X1 _25085_ ( .A1(_04315_ ), .A2(_04319_ ), .A3(_04321_ ), .ZN(_04322_ ) );
AND2_X1 _25086_ ( .A1(_04217_ ), .A2(_04196_ ), .ZN(_04323_ ) );
INV_X1 _25087_ ( .A(_04323_ ), .ZN(_04324_ ) );
OR2_X1 _25088_ ( .A1(_04324_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04325_ ) );
CLKBUF_X2 _25089_ ( .A(_04095_ ), .Z(_04326_ ) );
BUF_X2 _25090_ ( .A(_04320_ ), .Z(_04327_ ) );
OR3_X1 _25091_ ( .A1(_04326_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04327_ ), .ZN(_04328_ ) );
NAND3_X1 _25092_ ( .A1(_04322_ ), .A2(_04325_ ), .A3(_04328_ ), .ZN(_04329_ ) );
INV_X1 _25093_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04330_ ) );
BUF_X2 _25094_ ( .A(_04045_ ), .Z(_04331_ ) );
BUF_X2 _25095_ ( .A(_04331_ ), .Z(_04332_ ) );
CLKBUF_X2 _25096_ ( .A(_04332_ ), .Z(_04333_ ) );
AND4_X1 _25097_ ( .A1(_04330_ ), .A2(_04333_ ), .A3(_04242_ ), .A4(_04210_ ), .ZN(_04334_ ) );
NOR3_X1 _25098_ ( .A1(_04030_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04034_ ), .ZN(_04335_ ) );
NOR3_X1 _25099_ ( .A1(_04329_ ), .A2(_04334_ ), .A3(_04335_ ), .ZN(_04336_ ) );
OAI21_X1 _25100_ ( .A(_04336_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04219_ ), .ZN(_04337_ ) );
AOI211_X1 _25101_ ( .A(_04015_ ), .B(_04023_ ), .C1(_04005_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04338_ ) );
OAI221_X1 _25102_ ( .A(_04247_ ), .B1(_04248_ ), .B2(_04251_ ), .C1(_04337_ ), .C2(_04338_ ), .ZN(_04339_ ) );
BUF_X4 _25103_ ( .A(_03925_ ), .Z(_04340_ ) );
INV_X1 _25104_ ( .A(_04237_ ), .ZN(_04341_ ) );
NOR3_X1 _25105_ ( .A1(_04340_ ), .A2(_13185_ ), .A3(_04341_ ), .ZN(_04342_ ) );
OR3_X1 _25106_ ( .A1(_08547_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_1_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A3(_08560_ ), .ZN(_04343_ ) );
OAI21_X1 _25107_ ( .A(\io_master_rdata [30] ), .B1(_08547_ ), .B2(_08560_ ), .ZN(_04344_ ) );
NAND2_X1 _25108_ ( .A1(_04343_ ), .A2(_04344_ ), .ZN(_04345_ ) );
AND2_X1 _25109_ ( .A1(_04345_ ), .A2(fanout_net_1 ), .ZN(_04346_ ) );
INV_X1 _25110_ ( .A(_04346_ ), .ZN(_04347_ ) );
NOR3_X1 _25111_ ( .A1(_03899_ ), .A2(_03900_ ), .A3(_04347_ ), .ZN(_04348_ ) );
OR2_X1 _25112_ ( .A1(_03898_ ), .A2(_04348_ ), .ZN(_04349_ ) );
OAI21_X1 _25113_ ( .A(\lsu.io_in_bits_ren ), .B1(_04349_ ), .B2(_03917_ ), .ZN(_04350_ ) );
BUF_X2 _25114_ ( .A(_03926_ ), .Z(_04351_ ) );
NAND2_X1 _25115_ ( .A1(_04351_ ), .A2(\lsu.io_in_bits_rd_wdata [30] ), .ZN(_04352_ ) );
NAND2_X1 _25116_ ( .A1(_04350_ ), .A2(_04352_ ), .ZN(\lsu.io_out_bits_rd_wdata [30] ) );
BUF_X4 _25117_ ( .A(_03925_ ), .Z(_04353_ ) );
AOI21_X1 _25118_ ( .A(_04342_ ), .B1(\lsu.io_out_bits_rd_wdata [30] ), .B2(_04353_ ), .ZN(_04354_ ) );
MUX2_X1 _25119_ ( .A(_04354_ ), .B(_01720_ ), .S(_04228_ ), .Z(_04355_ ) );
OAI21_X1 _25120_ ( .A(_04339_ ), .B1(_04355_ ), .B2(\idu.rs_reg ), .ZN(\idu.io_out_bits_rs1_data [30] ) );
BUF_X4 _25121_ ( .A(_04228_ ), .Z(_04356_ ) );
NAND2_X1 _25122_ ( .A1(\exu.io_out_bits_rd_wdata [21] ), .A2(_04356_ ), .ZN(_04357_ ) );
INV_X1 _25123_ ( .A(_03916_ ), .ZN(_04358_ ) );
NOR3_X1 _25124_ ( .A1(_00967_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_10_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A3(_00969_ ), .ZN(_04359_ ) );
AOI21_X1 _25125_ ( .A(_04359_ ), .B1(_08563_ ), .B2(\io_master_rdata [21] ), .ZN(_04360_ ) );
NOR2_X1 _25126_ ( .A1(_04360_ ), .A2(_10989_ ), .ZN(_04361_ ) );
INV_X1 _25127_ ( .A(_04361_ ), .ZN(_04362_ ) );
OR3_X1 _25128_ ( .A1(_08547_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_2_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A3(_08560_ ), .ZN(_04363_ ) );
OAI21_X1 _25129_ ( .A(\io_master_rdata [29] ), .B1(_00967_ ), .B2(_00969_ ), .ZN(_04364_ ) );
NAND2_X1 _25130_ ( .A1(_04363_ ), .A2(_04364_ ), .ZN(_04365_ ) );
AND2_X1 _25131_ ( .A1(_04365_ ), .A2(fanout_net_1 ), .ZN(_04366_ ) );
INV_X1 _25132_ ( .A(_04366_ ), .ZN(_04367_ ) );
MUX2_X1 _25133_ ( .A(_04362_ ), .B(_04367_ ), .S(\io_master_awaddr [0] ), .Z(_04368_ ) );
NOR2_X1 _25134_ ( .A1(_03882_ ), .A2(\io_master_awaddr [1] ), .ZN(_04369_ ) );
INV_X1 _25135_ ( .A(_04369_ ), .ZN(_04370_ ) );
OAI22_X1 _25136_ ( .A1(_04368_ ), .A2(_04370_ ), .B1(_03909_ ), .B2(_04362_ ), .ZN(_04371_ ) );
AOI22_X1 _25137_ ( .A1(_03897_ ), .A2(\lsu.io_in_bits_lh ), .B1(_04371_ ), .B2(\arbiter.io_lsu_arsize [1] ), .ZN(_04372_ ) );
AOI21_X1 _25138_ ( .A(_03927_ ), .B1(_04358_ ), .B2(_04372_ ), .ZN(_04373_ ) );
AND2_X1 _25139_ ( .A1(_03926_ ), .A2(\lsu.io_in_bits_rd_wdata [21] ), .ZN(_04374_ ) );
OR3_X1 _25140_ ( .A1(_04373_ ), .A2(_03930_ ), .A3(_04374_ ), .ZN(_04375_ ) );
NAND4_X1 _25141_ ( .A1(_03990_ ), .A2(\wbu.io_in_bits_rd_wdata [21] ), .A3(_03997_ ), .A4(_04010_ ), .ZN(_04376_ ) );
AOI21_X1 _25142_ ( .A(_03859_ ), .B1(_03931_ ), .B2(_04376_ ), .ZN(_04377_ ) );
NAND2_X1 _25143_ ( .A1(_04375_ ), .A2(_04377_ ), .ZN(_04378_ ) );
AOI21_X1 _25144_ ( .A(\idu.rs_reg ), .B1(_04357_ ), .B2(_04378_ ), .ZN(_04379_ ) );
INV_X1 _25145_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04380_ ) );
AND3_X1 _25146_ ( .A1(_04215_ ), .A2(_04380_ ), .A3(_04223_ ), .ZN(_04381_ ) );
INV_X1 _25147_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04382_ ) );
AND4_X1 _25148_ ( .A1(_04382_ ), .A2(_04216_ ), .A3(_04156_ ), .A4(_04159_ ), .ZN(_04383_ ) );
BUF_X2 _25149_ ( .A(_04073_ ), .Z(_04384_ ) );
BUF_X2 _25150_ ( .A(_04384_ ), .Z(_04385_ ) );
INV_X1 _25151_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04386_ ) );
NAND4_X1 _25152_ ( .A1(_04385_ ), .A2(_04110_ ), .A3(_04386_ ), .A4(_04283_ ), .ZN(_04387_ ) );
INV_X1 _25153_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_04388_ ) );
NAND3_X1 _25154_ ( .A1(_04058_ ), .A2(_04388_ ), .A3(_11098_ ), .ZN(_04389_ ) );
OAI21_X1 _25155_ ( .A(_04389_ ), .B1(_04054_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04390_ ) );
INV_X1 _25156_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04391_ ) );
BUF_X4 _25157_ ( .A(_04063_ ), .Z(_04392_ ) );
AOI21_X1 _25158_ ( .A(_04390_ ), .B1(_04391_ ), .B2(_04392_ ), .ZN(_04393_ ) );
OR2_X1 _25159_ ( .A1(_04070_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04394_ ) );
AND2_X2 _25160_ ( .A1(_04162_ ), .A2(_11097_ ), .ZN(_04395_ ) );
INV_X1 _25161_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04396_ ) );
AOI22_X1 _25162_ ( .A1(_04395_ ), .A2(_04396_ ), .B1(_04039_ ), .B2(_04077_ ), .ZN(_04397_ ) );
AND3_X1 _25163_ ( .A1(_04393_ ), .A2(_04394_ ), .A3(_04397_ ), .ZN(_04398_ ) );
BUF_X2 _25164_ ( .A(_11098_ ), .Z(_04399_ ) );
AND3_X1 _25165_ ( .A1(_04077_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04399_ ), .ZN(_04400_ ) );
NOR2_X1 _25166_ ( .A1(_04398_ ), .A2(_04400_ ), .ZN(_04401_ ) );
INV_X1 _25167_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04402_ ) );
CLKBUF_X2 _25168_ ( .A(_04074_ ), .Z(_04403_ ) );
AND4_X1 _25169_ ( .A1(_04402_ ), .A2(_04098_ ), .A3(_04403_ ), .A4(_04040_ ), .ZN(_04404_ ) );
NOR3_X1 _25170_ ( .A1(_04186_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03993_ ), .ZN(_04405_ ) );
NOR3_X1 _25171_ ( .A1(_04401_ ), .A2(_04404_ ), .A3(_04405_ ), .ZN(_04406_ ) );
INV_X1 _25172_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04407_ ) );
NAND3_X1 _25173_ ( .A1(_04257_ ), .A2(_04407_ ), .A3(_04384_ ), .ZN(_04408_ ) );
NAND2_X1 _25174_ ( .A1(_04406_ ), .A2(_04408_ ), .ZN(_04409_ ) );
INV_X1 _25175_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04410_ ) );
CLKBUF_X2 _25176_ ( .A(_04399_ ), .Z(_04411_ ) );
AND4_X1 _25177_ ( .A1(_04410_ ), .A2(_04331_ ), .A3(_04117_ ), .A4(_04411_ ), .ZN(_04412_ ) );
INV_X1 _25178_ ( .A(_04105_ ), .ZN(_04413_ ) );
BUF_X2 _25179_ ( .A(_04413_ ), .Z(_04414_ ) );
OAI21_X1 _25180_ ( .A(_04414_ ), .B1(_04101_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04415_ ) );
NOR3_X1 _25181_ ( .A1(_04409_ ), .A2(_04412_ ), .A3(_04415_ ), .ZN(_04416_ ) );
AND3_X1 _25182_ ( .A1(_04287_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04037_ ), .ZN(_04417_ ) );
OAI21_X1 _25183_ ( .A(_04387_ ), .B1(_04416_ ), .B2(_04417_ ), .ZN(_04418_ ) );
INV_X1 _25184_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04419_ ) );
AND3_X1 _25185_ ( .A1(_04287_ ), .A2(_04419_ ), .A3(_04118_ ), .ZN(_04420_ ) );
NOR4_X1 _25186_ ( .A1(_04125_ ), .A2(_04034_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04018_ ), .ZN(_04421_ ) );
NOR3_X1 _25187_ ( .A1(_04418_ ), .A2(_04420_ ), .A3(_04421_ ), .ZN(_04422_ ) );
INV_X1 _25188_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04423_ ) );
NAND4_X1 _25189_ ( .A1(_04150_ ), .A2(_04157_ ), .A3(_04423_ ), .A4(_04019_ ), .ZN(_04424_ ) );
INV_X1 _25190_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04425_ ) );
NAND4_X1 _25191_ ( .A1(_04109_ ), .A2(_04150_ ), .A3(_04425_ ), .A4(_04019_ ), .ZN(_04426_ ) );
AND3_X1 _25192_ ( .A1(_04422_ ), .A2(_04424_ ), .A3(_04426_ ), .ZN(_04427_ ) );
INV_X1 _25193_ ( .A(_04305_ ), .ZN(_04428_ ) );
OR2_X1 _25194_ ( .A1(_04140_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04429_ ) );
OR2_X1 _25195_ ( .A1(_04302_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04430_ ) );
NAND4_X1 _25196_ ( .A1(_04427_ ), .A2(_04428_ ), .A3(_04429_ ), .A4(_04430_ ), .ZN(_04431_ ) );
NAND4_X1 _25197_ ( .A1(_04167_ ), .A2(_04158_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04208_ ), .ZN(_04432_ ) );
AOI21_X1 _25198_ ( .A(_04383_ ), .B1(_04431_ ), .B2(_04432_ ), .ZN(_04433_ ) );
AND2_X1 _25199_ ( .A1(_04078_ ), .A2(_04019_ ), .ZN(_04434_ ) );
INV_X1 _25200_ ( .A(_04434_ ), .ZN(_04435_ ) );
OR2_X1 _25201_ ( .A1(_04435_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04436_ ) );
CLKBUF_X2 _25202_ ( .A(_04043_ ), .Z(_04437_ ) );
OR4_X1 _25203_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04126_ ), .A3(_04181_ ), .A4(_04437_ ), .ZN(_04438_ ) );
NAND3_X1 _25204_ ( .A1(_04433_ ), .A2(_04436_ ), .A3(_04438_ ), .ZN(_04439_ ) );
NOR3_X1 _25205_ ( .A1(_04187_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04320_ ), .ZN(_04440_ ) );
INV_X1 _25206_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04441_ ) );
AND4_X1 _25207_ ( .A1(_04000_ ), .A2(_04195_ ), .A3(_04441_ ), .A4(_10756_ ), .ZN(_04442_ ) );
NOR3_X1 _25208_ ( .A1(_04439_ ), .A2(_04440_ ), .A3(_04442_ ), .ZN(_04443_ ) );
BUF_X2 _25209_ ( .A(_04027_ ), .Z(_04444_ ) );
BUF_X2 _25210_ ( .A(_04111_ ), .Z(_04445_ ) );
AND2_X1 _25211_ ( .A1(_04444_ ), .A2(_04445_ ), .ZN(_04446_ ) );
INV_X1 _25212_ ( .A(_04446_ ), .ZN(_04447_ ) );
OR3_X1 _25213_ ( .A1(_04326_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04320_ ), .ZN(_04448_ ) );
OR2_X1 _25214_ ( .A1(_04202_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04449_ ) );
NAND4_X1 _25215_ ( .A1(_04443_ ), .A2(_04447_ ), .A3(_04448_ ), .A4(_04449_ ), .ZN(_04450_ ) );
BUF_X2 _25216_ ( .A(_04158_ ), .Z(_04451_ ) );
NAND4_X1 _25217_ ( .A1(_04445_ ), .A2(_04451_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04210_ ), .ZN(_04452_ ) );
AOI21_X1 _25218_ ( .A(_04381_ ), .B1(_04450_ ), .B2(_04452_ ), .ZN(_04453_ ) );
INV_X1 _25219_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04454_ ) );
BUF_X4 _25220_ ( .A(_04199_ ), .Z(_04455_ ) );
OAI211_X1 _25221_ ( .A(_04221_ ), .B(_10792_ ), .C1(_04454_ ), .C2(_04455_ ), .ZN(_04456_ ) );
AOI221_X4 _25222_ ( .A(_04240_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B2(_04250_ ), .C1(_04453_ ), .C2(_04456_ ), .ZN(_04457_ ) );
OR2_X1 _25223_ ( .A1(_04379_ ), .A2(_04457_ ), .ZN(\idu.io_out_bits_rs1_data [21] ) );
OR2_X1 _25224_ ( .A1(_04373_ ), .A2(_04374_ ), .ZN(\lsu.io_out_bits_rd_wdata [21] ) );
AOI21_X1 _25225_ ( .A(_03857_ ), .B1(_02005_ ), .B2(_02006_ ), .ZN(_04458_ ) );
BUF_X4 _25226_ ( .A(_03855_ ), .Z(_04459_ ) );
NOR2_X1 _25227_ ( .A1(_03898_ ), .A2(_03921_ ), .ZN(_04460_ ) );
INV_X1 _25228_ ( .A(_04460_ ), .ZN(_04461_ ) );
BUF_X4 _25229_ ( .A(_03882_ ), .Z(_04462_ ) );
BUF_X2 _25230_ ( .A(_00967_ ), .Z(_04463_ ) );
BUF_X2 _25231_ ( .A(_00969_ ), .Z(_04464_ ) );
NOR3_X1 _25232_ ( .A1(_04463_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_11_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A3(_04464_ ), .ZN(_04465_ ) );
AOI21_X1 _25233_ ( .A(_04465_ ), .B1(_08563_ ), .B2(\io_master_rdata [20] ), .ZN(_04466_ ) );
NOR2_X1 _25234_ ( .A1(_04466_ ), .A2(_10990_ ), .ZN(_04467_ ) );
NAND2_X1 _25235_ ( .A1(_04462_ ), .A2(_04467_ ), .ZN(_04468_ ) );
BUF_X2 _25236_ ( .A(_03905_ ), .Z(_04469_ ) );
OR3_X1 _25237_ ( .A1(_04463_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_3_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A3(_04464_ ), .ZN(_04470_ ) );
OAI21_X1 _25238_ ( .A(\io_master_rdata [28] ), .B1(_04463_ ), .B2(_00970_ ), .ZN(_04471_ ) );
AOI211_X1 _25239_ ( .A(_10990_ ), .B(_04469_ ), .C1(_04470_ ), .C2(_04471_ ), .ZN(_04472_ ) );
AOI21_X1 _25240_ ( .A(_04472_ ), .B1(_04467_ ), .B2(_04469_ ), .ZN(_04473_ ) );
OAI21_X1 _25241_ ( .A(_04468_ ), .B1(_04370_ ), .B2(_04473_ ), .ZN(_04474_ ) );
AOI211_X1 _25242_ ( .A(_04461_ ), .B(_03917_ ), .C1(\arbiter.io_lsu_arsize [1] ), .C2(_04474_ ), .ZN(_04475_ ) );
NOR2_X1 _25243_ ( .A1(\lsu.io_in_bits_ren ), .A2(\lsu.io_in_bits_rd_wdata [20] ), .ZN(_04476_ ) );
NOR2_X1 _25244_ ( .A1(_04475_ ), .A2(_04476_ ), .ZN(\lsu.io_out_bits_rd_wdata [20] ) );
NOR2_X1 _25245_ ( .A1(\lsu.io_out_bits_rd_wdata [20] ), .A2(_03931_ ), .ZN(_04477_ ) );
NAND4_X1 _25246_ ( .A1(_03991_ ), .A2(\wbu.io_in_bits_rd_wdata [20] ), .A3(_03998_ ), .A4(_04011_ ), .ZN(_04478_ ) );
AOI211_X1 _25247_ ( .A(_04459_ ), .B(_04477_ ), .C1(_03932_ ), .C2(_04478_ ), .ZN(_04479_ ) );
OAI21_X1 _25248_ ( .A(_03851_ ), .B1(_04458_ ), .B2(_04479_ ), .ZN(_04480_ ) );
BUF_X4 _25249_ ( .A(_04246_ ), .Z(_04481_ ) );
BUF_X4 _25250_ ( .A(_04243_ ), .Z(_04482_ ) );
NAND3_X1 _25251_ ( .A1(_04222_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04482_ ), .ZN(_04483_ ) );
NAND3_X1 _25252_ ( .A1(_04207_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04212_ ), .ZN(_04484_ ) );
BUF_X2 _25253_ ( .A(_04294_ ), .Z(_04485_ ) );
NOR3_X1 _25254_ ( .A1(_04485_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04318_ ), .ZN(_04486_ ) );
NOR4_X1 _25255_ ( .A1(_04126_ ), .A2(_04034_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04254_ ), .ZN(_04487_ ) );
NOR2_X1 _25256_ ( .A1(_04487_ ), .A2(_04292_ ), .ZN(_04488_ ) );
NAND3_X1 _25257_ ( .A1(_04162_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04042_ ), .ZN(_04489_ ) );
INV_X1 _25258_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04490_ ) );
INV_X1 _25259_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04491_ ) );
NAND4_X1 _25260_ ( .A1(_04116_ ), .A2(_04148_ ), .A3(_04491_ ), .A4(_04040_ ), .ZN(_04492_ ) );
INV_X1 _25261_ ( .A(_04059_ ), .ZN(_04493_ ) );
OAI21_X1 _25262_ ( .A(_04492_ ), .B1(_04493_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_04494_ ) );
MUX2_X1 _25263_ ( .A(_04490_ ), .B(_04494_ ), .S(_04064_ ), .Z(_04495_ ) );
INV_X1 _25264_ ( .A(_04395_ ), .ZN(_04496_ ) );
BUF_X2 _25265_ ( .A(_04070_ ), .Z(_04497_ ) );
OAI21_X1 _25266_ ( .A(_04496_ ), .B1(_04497_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04498_ ) );
OAI21_X1 _25267_ ( .A(_04489_ ), .B1(_04495_ ), .B2(_04498_ ), .ZN(_04499_ ) );
INV_X1 _25268_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04500_ ) );
NAND4_X1 _25269_ ( .A1(_04155_ ), .A2(_04118_ ), .A3(_04500_ ), .A4(_04283_ ), .ZN(_04501_ ) );
OR2_X1 _25270_ ( .A1(_04085_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04502_ ) );
NAND3_X1 _25271_ ( .A1(_04499_ ), .A2(_04501_ ), .A3(_04502_ ), .ZN(_04503_ ) );
BUF_X2 _25272_ ( .A(_04257_ ), .Z(_04504_ ) );
INV_X1 _25273_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04505_ ) );
AND3_X1 _25274_ ( .A1(_04504_ ), .A2(_04505_ ), .A3(_04038_ ), .ZN(_04506_ ) );
NOR2_X1 _25275_ ( .A1(_04093_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04507_ ) );
NOR3_X1 _25276_ ( .A1(_04503_ ), .A2(_04506_ ), .A3(_04507_ ), .ZN(_04508_ ) );
BUF_X2 _25277_ ( .A(_04331_ ), .Z(_04509_ ) );
INV_X1 _25278_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04510_ ) );
NAND4_X1 _25279_ ( .A1(_04509_ ), .A2(_04119_ ), .A3(_04510_ ), .A4(_04114_ ), .ZN(_04511_ ) );
INV_X1 _25280_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04512_ ) );
CLKBUF_X2 _25281_ ( .A(_04042_ ), .Z(_04513_ ) );
NAND4_X1 _25282_ ( .A1(_04509_ ), .A2(_04146_ ), .A3(_04512_ ), .A4(_04513_ ), .ZN(_04514_ ) );
NAND3_X1 _25283_ ( .A1(_04508_ ), .A2(_04511_ ), .A3(_04514_ ), .ZN(_04515_ ) );
AND2_X2 _25284_ ( .A1(_04104_ ), .A2(_04116_ ), .ZN(_04516_ ) );
NOR2_X1 _25285_ ( .A1(_04414_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04517_ ) );
NAND2_X1 _25286_ ( .A1(_04384_ ), .A2(_04032_ ), .ZN(_04518_ ) );
BUF_X2 _25287_ ( .A(_04518_ ), .Z(_04519_ ) );
NOR3_X1 _25288_ ( .A1(_04519_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04019_ ), .ZN(_04520_ ) );
NOR4_X1 _25289_ ( .A1(_04515_ ), .A2(_04516_ ), .A3(_04517_ ), .A4(_04520_ ), .ZN(_04521_ ) );
BUF_X2 _25290_ ( .A(_04036_ ), .Z(_04522_ ) );
AND4_X1 _25291_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04170_ ), .A3(_04522_ ), .A4(_04295_ ), .ZN(_04523_ ) );
OAI21_X1 _25292_ ( .A(_04488_ ), .B1(_04521_ ), .B2(_04523_ ), .ZN(_04524_ ) );
BUF_X2 _25293_ ( .A(_04253_ ), .Z(_04525_ ) );
NAND3_X1 _25294_ ( .A1(_04444_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04525_ ), .ZN(_04526_ ) );
AOI21_X1 _25295_ ( .A(_04486_ ), .B1(_04524_ ), .B2(_04526_ ), .ZN(_04527_ ) );
BUF_X2 _25296_ ( .A(_04297_ ), .Z(_04528_ ) );
BUF_X2 _25297_ ( .A(_04151_ ), .Z(_04529_ ) );
INV_X1 _25298_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04530_ ) );
NAND4_X1 _25299_ ( .A1(_04528_ ), .A2(_04529_ ), .A3(_04530_ ), .A4(_04209_ ), .ZN(_04531_ ) );
OR2_X1 _25300_ ( .A1(_04303_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04532_ ) );
AND3_X1 _25301_ ( .A1(_04527_ ), .A2(_04531_ ), .A3(_04532_ ), .ZN(_04533_ ) );
BUF_X2 _25302_ ( .A(_04317_ ), .Z(_04534_ ) );
OR3_X1 _25303_ ( .A1(_04030_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04534_ ), .ZN(_04535_ ) );
BUF_X4 _25304_ ( .A(_04168_ ), .Z(_04536_ ) );
INV_X1 _25305_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04537_ ) );
BUF_X2 _25306_ ( .A(_04175_ ), .Z(_04538_ ) );
NAND4_X1 _25307_ ( .A1(_04223_ ), .A2(_04536_ ), .A3(_04537_ ), .A4(_04538_ ), .ZN(_04539_ ) );
NAND3_X1 _25308_ ( .A1(_04533_ ), .A2(_04535_ ), .A3(_04539_ ), .ZN(_04540_ ) );
INV_X1 _25309_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04541_ ) );
BUF_X2 _25310_ ( .A(_04167_ ), .Z(_04542_ ) );
AND4_X1 _25311_ ( .A1(_04541_ ), .A2(_04542_ ), .A3(_04528_ ), .A4(_04538_ ), .ZN(_04543_ ) );
BUF_X2 _25312_ ( .A(_04179_ ), .Z(_04544_ ) );
BUF_X2 _25313_ ( .A(_04184_ ), .Z(_04545_ ) );
NOR4_X1 _25314_ ( .A1(_04544_ ), .A2(_04534_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04545_ ), .ZN(_04546_ ) );
NOR3_X1 _25315_ ( .A1(_04540_ ), .A2(_04543_ ), .A3(_04546_ ), .ZN(_04547_ ) );
CLKBUF_X2 _25316_ ( .A(_04187_ ), .Z(_04548_ ) );
CLKBUF_X2 _25317_ ( .A(_04190_ ), .Z(_04549_ ) );
BUF_X2 _25318_ ( .A(_04549_ ), .Z(_04550_ ) );
OR3_X1 _25319_ ( .A1(_04548_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04550_ ), .ZN(_04551_ ) );
BUF_X4 _25320_ ( .A(_04197_ ), .Z(_04552_ ) );
BUF_X4 _25321_ ( .A(_04194_ ), .Z(_04553_ ) );
INV_X1 _25322_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04554_ ) );
BUF_X4 _25323_ ( .A(_04199_ ), .Z(_04555_ ) );
NAND4_X1 _25324_ ( .A1(_04552_ ), .A2(_04553_ ), .A3(_04554_ ), .A4(_04555_ ), .ZN(_04556_ ) );
NAND3_X1 _25325_ ( .A1(_04547_ ), .A2(_04551_ ), .A3(_04556_ ), .ZN(_04557_ ) );
BUF_X4 _25326_ ( .A(_04202_ ), .Z(_04558_ ) );
OAI21_X1 _25327_ ( .A(_04558_ ), .B1(_04204_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04559_ ) );
OAI21_X1 _25328_ ( .A(_04484_ ), .B1(_04557_ ), .B2(_04559_ ), .ZN(_04560_ ) );
OR3_X1 _25329_ ( .A1(_04030_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04034_ ), .ZN(_04561_ ) );
BUF_X4 _25330_ ( .A(_04221_ ), .Z(_04562_ ) );
INV_X1 _25331_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04563_ ) );
NAND3_X1 _25332_ ( .A1(_04562_ ), .A2(_04563_ ), .A3(_04224_ ), .ZN(_04564_ ) );
NAND3_X1 _25333_ ( .A1(_04560_ ), .A2(_04561_ ), .A3(_04564_ ), .ZN(_04565_ ) );
BUF_X4 _25334_ ( .A(_04015_ ), .Z(_04566_ ) );
BUF_X4 _25335_ ( .A(_04023_ ), .Z(_04567_ ) );
BUF_X4 _25336_ ( .A(_04005_ ), .Z(_04568_ ) );
AOI211_X1 _25337_ ( .A(_04566_ ), .B(_04567_ ), .C1(_04568_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04569_ ) );
OAI211_X1 _25338_ ( .A(_04481_ ), .B(_04483_ ), .C1(_04565_ ), .C2(_04569_ ), .ZN(_04570_ ) );
NAND2_X1 _25339_ ( .A1(_04480_ ), .A2(_04570_ ), .ZN(\idu.io_out_bits_rs1_data [20] ) );
BUF_X4 _25340_ ( .A(_04221_ ), .Z(_04571_ ) );
NAND3_X1 _25341_ ( .A1(_04571_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04243_ ), .ZN(_04572_ ) );
NOR2_X1 _25342_ ( .A1(_04165_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04573_ ) );
INV_X1 _25343_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04574_ ) );
AND4_X1 _25344_ ( .A1(_04574_ ), .A2(_04147_ ), .A3(_04151_ ), .A4(_04020_ ), .ZN(_04575_ ) );
AOI21_X1 _25345_ ( .A(_04575_ ), .B1(_04209_ ), .B2(_04067_ ), .ZN(_04576_ ) );
NOR3_X1 _25346_ ( .A1(_04485_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04183_ ), .ZN(_04577_ ) );
AND2_X1 _25347_ ( .A1(_04104_ ), .A2(_04144_ ), .ZN(_04578_ ) );
INV_X1 _25348_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04579_ ) );
AOI21_X1 _25349_ ( .A(_04292_ ), .B1(_04578_ ), .B2(_04579_ ), .ZN(_04580_ ) );
OR3_X1 _25350_ ( .A1(_04263_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10767_ ), .ZN(_04581_ ) );
MUX2_X1 _25351_ ( .A(_04581_ ), .B(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(_04053_ ), .Z(_04582_ ) );
OR2_X1 _25352_ ( .A1(_04064_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04583_ ) );
INV_X1 _25353_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04584_ ) );
AOI22_X1 _25354_ ( .A1(_04068_ ), .A2(_04584_ ), .B1(_04040_ ), .B2(_04162_ ), .ZN(_04585_ ) );
NAND3_X1 _25355_ ( .A1(_04582_ ), .A2(_04583_ ), .A3(_04585_ ), .ZN(_04586_ ) );
NAND3_X1 _25356_ ( .A1(_04162_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04041_ ), .ZN(_04587_ ) );
AOI21_X1 _25357_ ( .A(_04271_ ), .B1(_04586_ ), .B2(_04587_ ), .ZN(_04588_ ) );
AND3_X1 _25358_ ( .A1(_04078_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04041_ ), .ZN(_04589_ ) );
NOR2_X1 _25359_ ( .A1(_04588_ ), .A2(_04589_ ), .ZN(_04590_ ) );
NOR2_X1 _25360_ ( .A1(_04085_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04591_ ) );
BUF_X2 _25361_ ( .A(_04186_ ), .Z(_04592_ ) );
NOR3_X1 _25362_ ( .A1(_04592_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03994_ ), .ZN(_04593_ ) );
NOR3_X1 _25363_ ( .A1(_04590_ ), .A2(_04591_ ), .A3(_04593_ ), .ZN(_04594_ ) );
INV_X1 _25364_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04595_ ) );
NAND3_X1 _25365_ ( .A1(_04504_ ), .A2(_04595_ ), .A3(_04385_ ), .ZN(_04596_ ) );
INV_X1 _25366_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04597_ ) );
CLKBUF_X2 _25367_ ( .A(_04041_ ), .Z(_04598_ ) );
NAND4_X1 _25368_ ( .A1(_04331_ ), .A2(_04118_ ), .A3(_04597_ ), .A4(_04598_ ), .ZN(_04599_ ) );
AND3_X1 _25369_ ( .A1(_04594_ ), .A2(_04596_ ), .A3(_04599_ ), .ZN(_04600_ ) );
OR2_X1 _25370_ ( .A1(_04102_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04601_ ) );
OR2_X1 _25371_ ( .A1(_04414_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04602_ ) );
NAND3_X1 _25372_ ( .A1(_04600_ ), .A2(_04601_ ), .A3(_04602_ ), .ZN(_04603_ ) );
NOR3_X1 _25373_ ( .A1(_04519_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04019_ ), .ZN(_04604_ ) );
NOR3_X1 _25374_ ( .A1(_04603_ ), .A2(_04516_ ), .A3(_04604_ ), .ZN(_04605_ ) );
BUF_X2 _25375_ ( .A(_04287_ ), .Z(_04606_ ) );
AND3_X1 _25376_ ( .A1(_04606_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04170_ ), .ZN(_04607_ ) );
OAI21_X1 _25377_ ( .A(_04580_ ), .B1(_04605_ ), .B2(_04607_ ), .ZN(_04608_ ) );
NAND3_X1 _25378_ ( .A1(_04027_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04525_ ), .ZN(_04609_ ) );
AOI211_X1 _25379_ ( .A(_04139_ ), .B(_04577_ ), .C1(_04608_ ), .C2(_04609_ ), .ZN(_04610_ ) );
AND4_X1 _25380_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04171_ ), .A3(_04525_ ), .A4(_04208_ ), .ZN(_04611_ ) );
OAI21_X1 _25381_ ( .A(_04576_ ), .B1(_04610_ ), .B2(_04611_ ), .ZN(_04612_ ) );
NAND3_X1 _25382_ ( .A1(_04444_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04542_ ), .ZN(_04613_ ) );
AOI21_X1 _25383_ ( .A(_04573_ ), .B1(_04612_ ), .B2(_04613_ ), .ZN(_04614_ ) );
BUF_X2 _25384_ ( .A(_04171_ ), .Z(_04615_ ) );
INV_X1 _25385_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04616_ ) );
NAND4_X1 _25386_ ( .A1(_04536_ ), .A2(_04615_ ), .A3(_04616_ ), .A4(_04210_ ), .ZN(_04617_ ) );
OR4_X1 _25387_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04316_ ), .A3(_04182_ ), .A4(_04184_ ), .ZN(_04618_ ) );
AND3_X1 _25388_ ( .A1(_04614_ ), .A2(_04617_ ), .A3(_04618_ ), .ZN(_04619_ ) );
BUF_X2 _25389_ ( .A(_04333_ ), .Z(_04620_ ) );
BUF_X2 _25390_ ( .A(_04451_ ), .Z(_04621_ ) );
INV_X1 _25391_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04622_ ) );
CLKBUF_X2 _25392_ ( .A(_04310_ ), .Z(_04623_ ) );
CLKBUF_X2 _25393_ ( .A(_04623_ ), .Z(_04624_ ) );
NAND4_X1 _25394_ ( .A1(_04620_ ), .A2(_04621_ ), .A3(_04622_ ), .A4(_04624_ ), .ZN(_04625_ ) );
INV_X1 _25395_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04626_ ) );
NAND4_X1 _25396_ ( .A1(_04197_ ), .A2(_04194_ ), .A3(_04626_ ), .A4(_04199_ ), .ZN(_04627_ ) );
NAND3_X1 _25397_ ( .A1(_04619_ ), .A2(_04625_ ), .A3(_04627_ ), .ZN(_04628_ ) );
INV_X1 _25398_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04629_ ) );
AND4_X1 _25399_ ( .A1(_04629_ ), .A2(_04333_ ), .A3(_04615_ ), .A4(_04624_ ), .ZN(_04630_ ) );
NOR2_X1 _25400_ ( .A1(_04558_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04631_ ) );
NOR3_X1 _25401_ ( .A1(_04628_ ), .A2(_04630_ ), .A3(_04631_ ), .ZN(_04632_ ) );
BUF_X2 _25402_ ( .A(_04445_ ), .Z(_04633_ ) );
INV_X1 _25403_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04634_ ) );
NAND4_X1 _25404_ ( .A1(_04633_ ), .A2(_04621_ ), .A3(_04634_ ), .A4(_04212_ ), .ZN(_04635_ ) );
CLKBUF_X2 _25405_ ( .A(_04519_ ), .Z(_04636_ ) );
CLKBUF_X2 _25406_ ( .A(_04545_ ), .Z(_04637_ ) );
OR3_X1 _25407_ ( .A1(_04636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04637_ ), .ZN(_04638_ ) );
NAND3_X1 _25408_ ( .A1(_04632_ ), .A2(_04635_ ), .A3(_04638_ ), .ZN(_04639_ ) );
AOI211_X1 _25409_ ( .A(_04015_ ), .B(_04023_ ), .C1(_04005_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04640_ ) );
OAI211_X1 _25410_ ( .A(_04247_ ), .B(_04572_ ), .C1(_04639_ ), .C2(_04640_ ), .ZN(_04641_ ) );
INV_X1 _25411_ ( .A(_03898_ ), .ZN(_04642_ ) );
NOR3_X1 _25412_ ( .A1(_00967_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_12_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A3(_00969_ ), .ZN(_04643_ ) );
AOI21_X1 _25413_ ( .A(_04643_ ), .B1(_08563_ ), .B2(\io_master_rdata [19] ), .ZN(_04644_ ) );
NOR2_X1 _25414_ ( .A1(_04644_ ), .A2(_10990_ ), .ZN(_04645_ ) );
OR3_X1 _25415_ ( .A1(_00967_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_4_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A3(_00969_ ), .ZN(_04646_ ) );
OAI21_X1 _25416_ ( .A(\io_master_rdata [27] ), .B1(_00967_ ), .B2(_00969_ ), .ZN(_04647_ ) );
NAND2_X1 _25417_ ( .A1(_04646_ ), .A2(_04647_ ), .ZN(_04648_ ) );
AND2_X1 _25418_ ( .A1(_04648_ ), .A2(fanout_net_1 ), .ZN(_04649_ ) );
MUX2_X1 _25419_ ( .A(_04645_ ), .B(_04649_ ), .S(\io_master_awaddr [0] ), .Z(_04650_ ) );
AOI22_X1 _25420_ ( .A1(_04650_ ), .A2(_04369_ ), .B1(_04462_ ), .B2(_04645_ ), .ZN(_04651_ ) );
OAI21_X1 _25421_ ( .A(_04642_ ), .B1(_03900_ ), .B2(_04651_ ), .ZN(_04652_ ) );
OAI21_X1 _25422_ ( .A(\lsu.io_in_bits_ren ), .B1(_04652_ ), .B2(_03917_ ), .ZN(_04653_ ) );
NAND2_X1 _25423_ ( .A1(_04351_ ), .A2(\lsu.io_in_bits_rd_wdata [19] ), .ZN(_04654_ ) );
NAND2_X1 _25424_ ( .A1(_04653_ ), .A2(_04654_ ), .ZN(\lsu.io_out_bits_rd_wdata [19] ) );
NAND2_X1 _25425_ ( .A1(\lsu.io_out_bits_rd_wdata [19] ), .A2(_04353_ ), .ZN(_04655_ ) );
BUF_X4 _25426_ ( .A(_04237_ ), .Z(_04656_ ) );
BUF_X4 _25427_ ( .A(_08570_ ), .Z(_04657_ ) );
BUF_X4 _25428_ ( .A(_03923_ ), .Z(_04658_ ) );
OAI211_X1 _25429_ ( .A(\wbu.io_in_bits_rd_wdata [19] ), .B(_04656_ ), .C1(_04657_ ), .C2(_04658_ ), .ZN(_04659_ ) );
AOI21_X1 _25430_ ( .A(_04228_ ), .B1(_04655_ ), .B2(_04659_ ), .ZN(_04660_ ) );
AOI21_X1 _25431_ ( .A(_04660_ ), .B1(\exu.io_out_bits_rd_wdata [19] ), .B2(_04459_ ), .ZN(_04661_ ) );
OAI21_X1 _25432_ ( .A(_04641_ ), .B1(_04661_ ), .B2(\idu.rs_reg ), .ZN(\idu.io_out_bits_rs1_data [19] ) );
AND2_X1 _25433_ ( .A1(\exu.io_out_bits_rd_wdata [18] ), .A2(_04356_ ), .ZN(_04662_ ) );
OR3_X1 _25434_ ( .A1(_04463_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_5_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A3(_04464_ ), .ZN(_04663_ ) );
OAI21_X1 _25435_ ( .A(\io_master_rdata [26] ), .B1(_00968_ ), .B2(_00970_ ), .ZN(_04664_ ) );
AOI211_X1 _25436_ ( .A(_10990_ ), .B(_04469_ ), .C1(_04663_ ), .C2(_04664_ ), .ZN(_04665_ ) );
NOR3_X1 _25437_ ( .A1(_04463_ ), .A2(lsu_io_out_bits_rd_wdata_$_MUX__Y_13_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A3(_04464_ ), .ZN(_04666_ ) );
AOI21_X1 _25438_ ( .A(_04666_ ), .B1(_08563_ ), .B2(\io_master_rdata [18] ), .ZN(_04667_ ) );
NOR2_X1 _25439_ ( .A1(_04667_ ), .A2(_10990_ ), .ZN(_04668_ ) );
AOI21_X1 _25440_ ( .A(_04665_ ), .B1(_04668_ ), .B2(_04469_ ), .ZN(_04669_ ) );
NOR3_X1 _25441_ ( .A1(_04669_ ), .A2(\io_master_awaddr [1] ), .A3(_03882_ ), .ZN(_04670_ ) );
AND2_X1 _25442_ ( .A1(_03882_ ), .A2(_04668_ ), .ZN(_04671_ ) );
OAI21_X1 _25443_ ( .A(\arbiter.io_lsu_arsize [1] ), .B1(_04670_ ), .B2(_04671_ ), .ZN(_04672_ ) );
NAND2_X1 _25444_ ( .A1(_04642_ ), .A2(_04672_ ), .ZN(_04673_ ) );
OAI21_X1 _25445_ ( .A(\lsu.io_in_bits_ren ), .B1(_04673_ ), .B2(_03917_ ), .ZN(_04674_ ) );
NAND2_X1 _25446_ ( .A1(_04351_ ), .A2(\lsu.io_in_bits_rd_wdata [18] ), .ZN(_04675_ ) );
NAND2_X1 _25447_ ( .A1(_04674_ ), .A2(_04675_ ), .ZN(\lsu.io_out_bits_rd_wdata [18] ) );
NAND2_X1 _25448_ ( .A1(\lsu.io_out_bits_rd_wdata [18] ), .A2(_04353_ ), .ZN(_04676_ ) );
OAI211_X1 _25449_ ( .A(\wbu.io_in_bits_rd_wdata [18] ), .B(_04656_ ), .C1(_04657_ ), .C2(_04658_ ), .ZN(_04677_ ) );
AOI21_X1 _25450_ ( .A(_04356_ ), .B1(_04676_ ), .B2(_04677_ ), .ZN(_04678_ ) );
OAI21_X1 _25451_ ( .A(_03851_ ), .B1(_04662_ ), .B2(_04678_ ), .ZN(_04679_ ) );
NAND3_X1 _25452_ ( .A1(_04222_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04482_ ), .ZN(_04680_ ) );
NAND4_X1 _25453_ ( .A1(_04150_ ), .A2(_04038_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04129_ ), .ZN(_04681_ ) );
NAND3_X1 _25454_ ( .A1(_04287_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04117_ ), .ZN(_04682_ ) );
INV_X1 _25455_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04683_ ) );
AND4_X1 _25456_ ( .A1(_04683_ ), .A2(_04045_ ), .A3(_04098_ ), .A4(_04040_ ), .ZN(_04684_ ) );
OR3_X1 _25457_ ( .A1(_04263_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10766_ ), .ZN(_04685_ ) );
OAI21_X1 _25458_ ( .A(_04685_ ), .B1(_04054_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04686_ ) );
NOR2_X1 _25459_ ( .A1(_04069_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04687_ ) );
INV_X1 _25460_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04688_ ) );
AND4_X1 _25461_ ( .A1(_04688_ ), .A2(_04061_ ), .A3(_04050_ ), .A4(_11096_ ), .ZN(_04689_ ) );
NOR3_X1 _25462_ ( .A1(_04686_ ), .A2(_04687_ ), .A3(_04689_ ), .ZN(_04690_ ) );
OAI21_X1 _25463_ ( .A(_04690_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04496_ ), .ZN(_04691_ ) );
INV_X1 _25464_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04692_ ) );
AND3_X1 _25465_ ( .A1(_04077_ ), .A2(_04692_ ), .A3(_11097_ ), .ZN(_04693_ ) );
INV_X1 _25466_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04694_ ) );
AND4_X1 _25467_ ( .A1(_04694_ ), .A2(_04061_ ), .A3(_04066_ ), .A4(_11097_ ), .ZN(_04695_ ) );
OR3_X1 _25468_ ( .A1(_04691_ ), .A2(_04693_ ), .A3(_04695_ ), .ZN(_04696_ ) );
NOR3_X1 _25469_ ( .A1(_04186_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10767_ ), .ZN(_04697_ ) );
OAI22_X1 _25470_ ( .A1(_04093_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_04094_ ), .B2(_10767_ ), .ZN(_04698_ ) );
OR3_X1 _25471_ ( .A1(_04696_ ), .A2(_04697_ ), .A3(_04698_ ), .ZN(_04699_ ) );
NAND3_X1 _25472_ ( .A1(_04047_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04041_ ), .ZN(_04700_ ) );
AOI21_X1 _25473_ ( .A(_04684_ ), .B1(_04699_ ), .B2(_04700_ ), .ZN(_04701_ ) );
OAI21_X1 _25474_ ( .A(_04701_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04414_ ), .ZN(_04702_ ) );
INV_X1 _25475_ ( .A(_04516_ ), .ZN(_04703_ ) );
INV_X1 _25476_ ( .A(_04285_ ), .ZN(_04704_ ) );
OAI21_X1 _25477_ ( .A(_04703_ ), .B1(_04704_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04705_ ) );
OAI21_X1 _25478_ ( .A(_04682_ ), .B1(_04702_ ), .B2(_04705_ ), .ZN(_04706_ ) );
INV_X1 _25479_ ( .A(_04578_ ), .ZN(_04707_ ) );
OAI21_X1 _25480_ ( .A(_04706_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04707_ ), .ZN(_04708_ ) );
OAI21_X1 _25481_ ( .A(_04681_ ), .B1(_04708_ ), .B2(_04292_ ), .ZN(_04709_ ) );
MUX2_X1 _25482_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_04709_ ), .S(_04136_ ), .Z(_04710_ ) );
BUF_X2 _25483_ ( .A(_04140_ ), .Z(_04711_ ) );
OR2_X1 _25484_ ( .A1(_04711_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04712_ ) );
OR2_X1 _25485_ ( .A1(_04303_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04713_ ) );
AND3_X1 _25486_ ( .A1(_04710_ ), .A2(_04712_ ), .A3(_04713_ ), .ZN(_04714_ ) );
INV_X1 _25487_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04715_ ) );
NAND4_X1 _25488_ ( .A1(_04168_ ), .A2(_04451_ ), .A3(_04715_ ), .A4(_04313_ ), .ZN(_04716_ ) );
INV_X1 _25489_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04717_ ) );
NAND4_X1 _25490_ ( .A1(_04217_ ), .A2(_04309_ ), .A3(_04717_ ), .A4(_04313_ ), .ZN(_04718_ ) );
NAND3_X1 _25491_ ( .A1(_04714_ ), .A2(_04716_ ), .A3(_04718_ ), .ZN(_04719_ ) );
NOR2_X1 _25492_ ( .A1(_04435_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04720_ ) );
INV_X1 _25493_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04721_ ) );
AND4_X1 _25494_ ( .A1(_04721_ ), .A2(_04241_ ), .A3(_04167_ ), .A4(_04310_ ), .ZN(_04722_ ) );
NOR3_X1 _25495_ ( .A1(_04719_ ), .A2(_04720_ ), .A3(_04722_ ), .ZN(_04723_ ) );
OR3_X1 _25496_ ( .A1(_04188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04191_ ), .ZN(_04724_ ) );
AND3_X1 _25497_ ( .A1(_04723_ ), .A2(_04324_ ), .A3(_04724_ ), .ZN(_04725_ ) );
AOI21_X1 _25498_ ( .A(_04725_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04323_ ), .ZN(_04726_ ) );
INV_X1 _25499_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04727_ ) );
BUF_X2 _25500_ ( .A(_04615_ ), .Z(_04728_ ) );
AND4_X1 _25501_ ( .A1(_04727_ ), .A2(_04620_ ), .A3(_04728_ ), .A4(_04624_ ), .ZN(_04729_ ) );
NOR2_X1 _25502_ ( .A1(_04558_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04730_ ) );
NOR3_X1 _25503_ ( .A1(_04726_ ), .A2(_04729_ ), .A3(_04730_ ), .ZN(_04731_ ) );
OR3_X1 _25504_ ( .A1(_04030_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04034_ ), .ZN(_04732_ ) );
INV_X1 _25505_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04733_ ) );
NAND3_X1 _25506_ ( .A1(_04562_ ), .A2(_04733_ ), .A3(_04224_ ), .ZN(_04734_ ) );
NAND3_X1 _25507_ ( .A1(_04731_ ), .A2(_04732_ ), .A3(_04734_ ), .ZN(_04735_ ) );
AOI211_X1 _25508_ ( .A(_04566_ ), .B(_04567_ ), .C1(_04568_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04736_ ) );
OAI211_X1 _25509_ ( .A(_04481_ ), .B(_04680_ ), .C1(_04735_ ), .C2(_04736_ ), .ZN(_04737_ ) );
NAND2_X1 _25510_ ( .A1(_04679_ ), .A2(_04737_ ), .ZN(\idu.io_out_bits_rs1_data [18] ) );
BUF_X4 _25511_ ( .A(_04229_ ), .Z(_04738_ ) );
NOR2_X1 _25512_ ( .A1(_02254_ ), .A2(_04738_ ), .ZN(_04739_ ) );
INV_X1 _25513_ ( .A(\io_master_awaddr [7] ), .ZN(_04740_ ) );
INV_X1 _25514_ ( .A(\io_master_awaddr [28] ), .ZN(_04741_ ) );
AND4_X1 _25515_ ( .A1(_08538_ ), .A2(_04741_ ), .A3(_08534_ ), .A4(\io_master_awaddr [25] ), .ZN(_04742_ ) );
AND4_X1 _25516_ ( .A1(_04740_ ), .A2(_08556_ ), .A3(_08537_ ), .A4(_04742_ ), .ZN(_04743_ ) );
NOR4_X1 _25517_ ( .A1(\io_master_awaddr [11] ), .A2(\io_master_awaddr [8] ), .A3(\io_master_awaddr [27] ), .A4(\io_master_awaddr [26] ), .ZN(_04744_ ) );
INV_X1 _25518_ ( .A(\io_master_awaddr [9] ), .ZN(_04745_ ) );
NAND4_X1 _25519_ ( .A1(_04744_ ), .A2(_03867_ ), .A3(_04745_ ), .A4(_03883_ ), .ZN(_04746_ ) );
INV_X1 _25520_ ( .A(\io_master_awaddr [6] ), .ZN(_04747_ ) );
NAND4_X1 _25521_ ( .A1(_08543_ ), .A2(_08544_ ), .A3(_04747_ ), .A4(_08536_ ), .ZN(_04748_ ) );
NOR3_X1 _25522_ ( .A1(_04746_ ), .A2(_03861_ ), .A3(_04748_ ), .ZN(_04749_ ) );
AND2_X1 _25523_ ( .A1(_04743_ ), .A2(_04749_ ), .ZN(_04750_ ) );
INV_X1 _25524_ ( .A(_04750_ ), .ZN(_04751_ ) );
AOI21_X1 _25525_ ( .A(_10989_ ), .B1(_04751_ ), .B2(_11627_ ), .ZN(_04752_ ) );
NAND4_X1 _25526_ ( .A1(_04743_ ), .A2(_04749_ ), .A3(fanout_net_1 ), .A4(lsu_io_out_bits_rd_wdata_$_MUX__Y_14_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .ZN(_04753_ ) );
NAND4_X1 _25527_ ( .A1(_04752_ ), .A2(_08542_ ), .A3(_03880_ ), .A4(_04753_ ), .ZN(_04754_ ) );
AND3_X1 _25528_ ( .A1(_04752_ ), .A2(_04469_ ), .A3(_04753_ ), .ZN(_04755_ ) );
OAI21_X1 _25529_ ( .A(fanout_net_1 ), .B1(_04750_ ), .B2(\io_master_rdata [25] ), .ZN(_04756_ ) );
AND4_X1 _25530_ ( .A1(fanout_net_1 ), .A2(_04743_ ), .A3(_04749_ ), .A4(lsu_io_out_bits_rd_wdata_$_MUX__Y_6_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .ZN(_04757_ ) );
NOR2_X1 _25531_ ( .A1(_04756_ ), .A2(_04757_ ), .ZN(_04758_ ) );
AOI21_X1 _25532_ ( .A(_04755_ ), .B1(\io_master_awaddr [0] ), .B2(_04758_ ), .ZN(_04759_ ) );
OAI21_X1 _25533_ ( .A(_04754_ ), .B1(_04759_ ), .B2(_04370_ ), .ZN(_04760_ ) );
AOI22_X1 _25534_ ( .A1(_03897_ ), .A2(\lsu.io_in_bits_lh ), .B1(\arbiter.io_lsu_arsize [1] ), .B2(_04760_ ), .ZN(_04761_ ) );
AOI21_X1 _25535_ ( .A(_04351_ ), .B1(_04358_ ), .B2(_04761_ ), .ZN(_04762_ ) );
AND2_X1 _25536_ ( .A1(_04351_ ), .A2(\lsu.io_in_bits_rd_wdata [17] ), .ZN(_04763_ ) );
OAI21_X1 _25537_ ( .A(_04353_ ), .B1(_04762_ ), .B2(_04763_ ), .ZN(_04764_ ) );
OAI211_X1 _25538_ ( .A(\wbu.io_in_bits_rd_wdata [17] ), .B(_04656_ ), .C1(_04657_ ), .C2(_04658_ ), .ZN(_04765_ ) );
AOI21_X1 _25539_ ( .A(_04228_ ), .B1(_04764_ ), .B2(_04765_ ), .ZN(_04766_ ) );
OAI21_X1 _25540_ ( .A(_03850_ ), .B1(_04739_ ), .B2(_04766_ ), .ZN(_04767_ ) );
AND3_X1 _25541_ ( .A1(_04444_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04633_ ), .ZN(_04768_ ) );
AND3_X1 _25542_ ( .A1(_04606_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04170_ ), .ZN(_04769_ ) );
OR2_X1 _25543_ ( .A1(_04070_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04770_ ) );
NOR3_X1 _25544_ ( .A1(_04294_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_03992_ ), .ZN(_04771_ ) );
INV_X1 _25545_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04772_ ) );
AOI21_X1 _25546_ ( .A(_04771_ ), .B1(_04053_ ), .B2(_04772_ ), .ZN(_04773_ ) );
INV_X1 _25547_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04774_ ) );
NAND4_X1 _25548_ ( .A1(_04144_ ), .A2(_04149_ ), .A3(_04774_ ), .A4(_04080_ ), .ZN(_04775_ ) );
AND3_X1 _25549_ ( .A1(_04770_ ), .A2(_04773_ ), .A3(_04775_ ), .ZN(_04776_ ) );
OAI21_X1 _25550_ ( .A(_04776_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04496_ ), .ZN(_04777_ ) );
INV_X1 _25551_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04778_ ) );
AND3_X1 _25552_ ( .A1(_04078_ ), .A2(_04778_ ), .A3(_04282_ ), .ZN(_04779_ ) );
NOR4_X1 _25553_ ( .A1(_04125_ ), .A2(_04180_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04017_ ), .ZN(_04780_ ) );
NOR3_X1 _25554_ ( .A1(_04777_ ), .A2(_04779_ ), .A3(_04780_ ), .ZN(_04781_ ) );
OR3_X1 _25555_ ( .A1(_04592_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04138_ ), .ZN(_04782_ ) );
INV_X1 _25556_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04783_ ) );
AOI22_X1 _25557_ ( .A1(_04783_ ), .A2(_04092_ ), .B1(_04048_ ), .B2(_04283_ ), .ZN(_04784_ ) );
AND3_X1 _25558_ ( .A1(_04781_ ), .A2(_04782_ ), .A3(_04784_ ), .ZN(_04785_ ) );
AND3_X1 _25559_ ( .A1(_04048_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04043_ ), .ZN(_04786_ ) );
OAI221_X1 _25560_ ( .A(_04414_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04102_ ), .C1(_04785_ ), .C2(_04786_ ), .ZN(_04787_ ) );
NAND4_X1 _25561_ ( .A1(_04445_ ), .A2(_04157_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04437_ ), .ZN(_04788_ ) );
NAND2_X1 _25562_ ( .A1(_04787_ ), .A2(_04788_ ), .ZN(_04789_ ) );
NOR3_X1 _25563_ ( .A1(_04519_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04254_ ), .ZN(_04790_ ) );
NOR2_X1 _25564_ ( .A1(_04516_ ), .A2(_04790_ ), .ZN(_04791_ ) );
AOI21_X1 _25565_ ( .A(_04769_ ), .B1(_04789_ ), .B2(_04791_ ), .ZN(_04792_ ) );
INV_X1 _25566_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04793_ ) );
AND4_X1 _25567_ ( .A1(_04793_ ), .A2(_04147_ ), .A3(_04445_ ), .A4(_04183_ ), .ZN(_04794_ ) );
NOR4_X1 _25568_ ( .A1(_04029_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10597_ ), .A4(_10600_ ), .ZN(_04795_ ) );
NOR3_X1 _25569_ ( .A1(_04792_ ), .A2(_04794_ ), .A3(_04795_ ), .ZN(_04796_ ) );
OR3_X1 _25570_ ( .A1(_04485_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04318_ ), .ZN(_04797_ ) );
OR2_X1 _25571_ ( .A1(_04711_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04798_ ) );
NAND3_X1 _25572_ ( .A1(_04796_ ), .A2(_04797_ ), .A3(_04798_ ), .ZN(_04799_ ) );
NOR2_X1 _25573_ ( .A1(_04303_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04800_ ) );
INV_X1 _25574_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04801_ ) );
AND4_X1 _25575_ ( .A1(_04801_ ), .A2(_04309_ ), .A3(_04158_ ), .A4(_04313_ ), .ZN(_04802_ ) );
NOR3_X1 _25576_ ( .A1(_04799_ ), .A2(_04800_ ), .A3(_04802_ ), .ZN(_04803_ ) );
INV_X1 _25577_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04804_ ) );
NAND4_X1 _25578_ ( .A1(_04223_ ), .A2(_04536_ ), .A3(_04804_ ), .A4(_04210_ ), .ZN(_04805_ ) );
OR2_X1 _25579_ ( .A1(_04435_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04806_ ) );
NAND3_X1 _25580_ ( .A1(_04803_ ), .A2(_04805_ ), .A3(_04806_ ), .ZN(_04807_ ) );
INV_X1 _25581_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04808_ ) );
AND4_X1 _25582_ ( .A1(_04808_ ), .A2(_04242_ ), .A3(_04542_ ), .A4(_04538_ ), .ZN(_04809_ ) );
NOR3_X1 _25583_ ( .A1(_04548_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04550_ ), .ZN(_04810_ ) );
NOR3_X1 _25584_ ( .A1(_04807_ ), .A2(_04809_ ), .A3(_04810_ ), .ZN(_04811_ ) );
INV_X1 _25585_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04812_ ) );
NAND4_X1 _25586_ ( .A1(_04552_ ), .A2(_04553_ ), .A3(_04812_ ), .A4(_04555_ ), .ZN(_04813_ ) );
OR3_X1 _25587_ ( .A1(_04326_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04550_ ), .ZN(_04814_ ) );
AND3_X1 _25588_ ( .A1(_04811_ ), .A2(_04813_ ), .A3(_04814_ ), .ZN(_04815_ ) );
NOR2_X1 _25589_ ( .A1(_04558_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04816_ ) );
NOR2_X1 _25590_ ( .A1(_04816_ ), .A2(_04446_ ), .ZN(_04817_ ) );
AOI21_X1 _25591_ ( .A(_04768_ ), .B1(_04815_ ), .B2(_04817_ ), .ZN(_04818_ ) );
CLKBUF_X2 _25592_ ( .A(_04320_ ), .Z(_04819_ ) );
CLKBUF_X2 _25593_ ( .A(_04819_ ), .Z(_04820_ ) );
NOR3_X1 _25594_ ( .A1(_04636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04820_ ), .ZN(_04821_ ) );
AOI211_X1 _25595_ ( .A(_04015_ ), .B(_04023_ ), .C1(_04005_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04822_ ) );
NOR3_X1 _25596_ ( .A1(_04818_ ), .A2(_04821_ ), .A3(_04822_ ), .ZN(_04823_ ) );
INV_X1 _25597_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_04824_ ) );
OAI21_X1 _25598_ ( .A(_04247_ ), .B1(_04824_ ), .B2(_04251_ ), .ZN(_04825_ ) );
OAI21_X1 _25599_ ( .A(_04767_ ), .B1(_04823_ ), .B2(_04825_ ), .ZN(\idu.io_out_bits_rs1_data [17] ) );
OR2_X1 _25600_ ( .A1(_04762_ ), .A2(_04763_ ), .ZN(\lsu.io_out_bits_rd_wdata [17] ) );
AOI21_X1 _25601_ ( .A(_03857_ ), .B1(_02326_ ), .B2(_02327_ ), .ZN(_04826_ ) );
OR4_X1 _25602_ ( .A1(_10988_ ), .A2(_00967_ ), .A3(lsu_io_out_bits_rd_wdata_$_MUX__Y_7_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A4(_00969_ ), .ZN(_04827_ ) );
OAI211_X1 _25603_ ( .A(fanout_net_1 ), .B(\io_master_rdata [24] ), .C1(_04463_ ), .C2(_04464_ ), .ZN(_04828_ ) );
AND2_X1 _25604_ ( .A1(_04827_ ), .A2(_04828_ ), .ZN(_04829_ ) );
AOI21_X1 _25605_ ( .A(_10989_ ), .B1(_04751_ ), .B2(_11636_ ), .ZN(_04830_ ) );
NAND4_X1 _25606_ ( .A1(_04743_ ), .A2(_04749_ ), .A3(fanout_net_1 ), .A4(lsu_io_out_bits_rd_wdata_$_MUX__Y_15_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .ZN(_04831_ ) );
NAND2_X1 _25607_ ( .A1(_04830_ ), .A2(_04831_ ), .ZN(_04832_ ) );
MUX2_X1 _25608_ ( .A(_04829_ ), .B(_04832_ ), .S(_04469_ ), .Z(_04833_ ) );
OAI22_X1 _25609_ ( .A1(_04833_ ), .A2(_04370_ ), .B1(_03909_ ), .B2(_04832_ ), .ZN(_04834_ ) );
AOI211_X1 _25610_ ( .A(_04461_ ), .B(_03916_ ), .C1(\arbiter.io_lsu_arsize [1] ), .C2(_04834_ ), .ZN(_04835_ ) );
NOR2_X1 _25611_ ( .A1(\lsu.io_in_bits_ren ), .A2(\lsu.io_in_bits_rd_wdata [16] ), .ZN(_04836_ ) );
NOR2_X1 _25612_ ( .A1(_04835_ ), .A2(_04836_ ), .ZN(\lsu.io_out_bits_rd_wdata [16] ) );
NOR2_X1 _25613_ ( .A1(\lsu.io_out_bits_rd_wdata [16] ), .A2(_03931_ ), .ZN(_04837_ ) );
NAND4_X1 _25614_ ( .A1(_03991_ ), .A2(\wbu.io_in_bits_rd_wdata [16] ), .A3(_03998_ ), .A4(_04011_ ), .ZN(_04838_ ) );
AOI211_X1 _25615_ ( .A(_04459_ ), .B(_04837_ ), .C1(_03932_ ), .C2(_04838_ ), .ZN(_04839_ ) );
OAI21_X1 _25616_ ( .A(_03851_ ), .B1(_04826_ ), .B2(_04839_ ), .ZN(_04840_ ) );
NAND3_X1 _25617_ ( .A1(_04222_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04482_ ), .ZN(_04841_ ) );
BUF_X2 _25618_ ( .A(_04310_ ), .Z(_04842_ ) );
NAND3_X1 _25619_ ( .A1(_04062_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04842_ ), .ZN(_04843_ ) );
OR3_X1 _25620_ ( .A1(_04519_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04129_ ), .ZN(_04844_ ) );
AND2_X1 _25621_ ( .A1(_04047_ ), .A2(_04041_ ), .ZN(_04845_ ) );
INV_X1 _25622_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04846_ ) );
AOI22_X1 _25623_ ( .A1(_04845_ ), .A2(_04846_ ), .B1(_04283_ ), .B2(_04099_ ), .ZN(_04847_ ) );
NAND4_X1 _25624_ ( .A1(_04384_ ), .A2(_04154_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04041_ ), .ZN(_04848_ ) );
NAND4_X1 _25625_ ( .A1(_04098_ ), .A2(_04148_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04399_ ), .ZN(_04849_ ) );
INV_X1 _25626_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04850_ ) );
NAND3_X1 _25627_ ( .A1(_04051_ ), .A2(_04850_ ), .A3(_11099_ ), .ZN(_04851_ ) );
OAI21_X1 _25628_ ( .A(_04851_ ), .B1(_04493_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_04852_ ) );
OAI21_X1 _25629_ ( .A(_04849_ ), .B1(_04852_ ), .B2(_04392_ ), .ZN(_04853_ ) );
OAI21_X1 _25630_ ( .A(_04853_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04497_ ), .ZN(_04854_ ) );
OAI21_X1 _25631_ ( .A(_04848_ ), .B1(_04854_ ), .B2(_04395_ ), .ZN(_04855_ ) );
INV_X1 _25632_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04856_ ) );
NAND3_X1 _25633_ ( .A1(_04078_ ), .A2(_04856_ ), .A3(_11101_ ), .ZN(_04857_ ) );
BUF_X2 _25634_ ( .A(_04403_ ), .Z(_04858_ ) );
INV_X1 _25635_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04859_ ) );
NAND4_X1 _25636_ ( .A1(_04145_ ), .A2(_04858_ ), .A3(_04859_ ), .A4(_04282_ ), .ZN(_04860_ ) );
NAND3_X1 _25637_ ( .A1(_04855_ ), .A2(_04857_ ), .A3(_04860_ ), .ZN(_04861_ ) );
NOR3_X1 _25638_ ( .A1(_04592_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03994_ ), .ZN(_04862_ ) );
NOR3_X1 _25639_ ( .A1(_04861_ ), .A2(_04092_ ), .A3(_04862_ ), .ZN(_04863_ ) );
AND3_X1 _25640_ ( .A1(_04504_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04108_ ), .ZN(_04864_ ) );
OAI21_X1 _25641_ ( .A(_04847_ ), .B1(_04863_ ), .B2(_04864_ ), .ZN(_04865_ ) );
NAND3_X1 _25642_ ( .A1(_04099_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04513_ ), .ZN(_04866_ ) );
AOI21_X1 _25643_ ( .A(_04105_ ), .B1(_04865_ ), .B2(_04866_ ), .ZN(_04867_ ) );
AND3_X1 _25644_ ( .A1(_04606_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04157_ ), .ZN(_04868_ ) );
OAI21_X1 _25645_ ( .A(_04844_ ), .B1(_04867_ ), .B2(_04868_ ), .ZN(_04869_ ) );
INV_X1 _25646_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04870_ ) );
AND4_X1 _25647_ ( .A1(_04870_ ), .A2(_04119_ ), .A3(_04111_ ), .A4(_04189_ ), .ZN(_04871_ ) );
NOR4_X1 _25648_ ( .A1(_04126_ ), .A2(_04034_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04173_ ), .ZN(_04872_ ) );
NOR3_X1 _25649_ ( .A1(_04869_ ), .A2(_04871_ ), .A3(_04872_ ), .ZN(_04873_ ) );
OR4_X1 _25650_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04131_ ), .A3(_10597_ ), .A4(_10600_ ), .ZN(_04874_ ) );
AND2_X1 _25651_ ( .A1(_04873_ ), .A2(_04874_ ), .ZN(_04875_ ) );
OAI21_X1 _25652_ ( .A(_04875_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04136_ ), .ZN(_04876_ ) );
OAI21_X1 _25653_ ( .A(_04303_ ), .B1(_04711_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04877_ ) );
OAI21_X1 _25654_ ( .A(_04843_ ), .B1(_04876_ ), .B2(_04877_ ), .ZN(_04878_ ) );
INV_X1 _25655_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04879_ ) );
NAND4_X1 _25656_ ( .A1(_04536_ ), .A2(_04451_ ), .A3(_04879_ ), .A4(_04538_ ), .ZN(_04880_ ) );
INV_X1 _25657_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04881_ ) );
NAND4_X1 _25658_ ( .A1(_04223_ ), .A2(_04542_ ), .A3(_04881_ ), .A4(_04538_ ), .ZN(_04882_ ) );
NAND3_X1 _25659_ ( .A1(_04878_ ), .A2(_04880_ ), .A3(_04882_ ), .ZN(_04883_ ) );
NOR2_X1 _25660_ ( .A1(_04435_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04884_ ) );
NOR4_X1 _25661_ ( .A1(_04179_ ), .A2(_04534_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04545_ ), .ZN(_04885_ ) );
NOR3_X1 _25662_ ( .A1(_04883_ ), .A2(_04884_ ), .A3(_04885_ ), .ZN(_04886_ ) );
INV_X1 _25663_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04887_ ) );
NAND4_X1 _25664_ ( .A1(_04620_ ), .A2(_04621_ ), .A3(_04887_ ), .A4(_04211_ ), .ZN(_04888_ ) );
INV_X1 _25665_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04889_ ) );
NAND4_X1 _25666_ ( .A1(_04552_ ), .A2(_04553_ ), .A3(_04889_ ), .A4(_04555_ ), .ZN(_04890_ ) );
NAND3_X1 _25667_ ( .A1(_04886_ ), .A2(_04888_ ), .A3(_04890_ ), .ZN(_04891_ ) );
NOR3_X1 _25668_ ( .A1(_04326_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04820_ ), .ZN(_04892_ ) );
INV_X1 _25669_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04893_ ) );
AND4_X1 _25670_ ( .A1(_04893_ ), .A2(_04333_ ), .A3(_04242_ ), .A4(_04624_ ), .ZN(_04894_ ) );
NOR3_X1 _25671_ ( .A1(_04891_ ), .A2(_04892_ ), .A3(_04894_ ), .ZN(_04895_ ) );
OR3_X1 _25672_ ( .A1(_04030_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04034_ ), .ZN(_04896_ ) );
OR3_X1 _25673_ ( .A1(_04636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04820_ ), .ZN(_04897_ ) );
NAND3_X1 _25674_ ( .A1(_04895_ ), .A2(_04896_ ), .A3(_04897_ ), .ZN(_04898_ ) );
AOI211_X1 _25675_ ( .A(_04566_ ), .B(_04567_ ), .C1(_04568_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04899_ ) );
OAI211_X1 _25676_ ( .A(_04481_ ), .B(_04841_ ), .C1(_04898_ ), .C2(_04899_ ), .ZN(_04900_ ) );
NAND2_X1 _25677_ ( .A1(_04840_ ), .A2(_04900_ ), .ZN(\idu.io_out_bits_rs1_data [16] ) );
AOI21_X1 _25678_ ( .A(_03857_ ), .B1(_02405_ ), .B2(_02406_ ), .ZN(_04901_ ) );
NOR2_X1 _25679_ ( .A1(\lsu.io_in_bits_lh ), .A2(\lsu.io_in_bits_lhu ), .ZN(_04902_ ) );
AND2_X1 _25680_ ( .A1(_04902_ ), .A2(_03900_ ), .ZN(_04903_ ) );
INV_X1 _25681_ ( .A(_04903_ ), .ZN(_04904_ ) );
AOI221_X4 _25682_ ( .A(_03921_ ), .B1(_03897_ ), .B2(_04904_ ), .C1(_03915_ ), .C2(\lsu.io_in_bits_lb ), .ZN(_04905_ ) );
NOR2_X1 _25683_ ( .A1(\lsu.io_in_bits_ren ), .A2(\lsu.io_in_bits_rd_wdata [15] ), .ZN(_04906_ ) );
NOR2_X1 _25684_ ( .A1(_04905_ ), .A2(_04906_ ), .ZN(\lsu.io_out_bits_rd_wdata [15] ) );
NOR2_X1 _25685_ ( .A1(\lsu.io_out_bits_rd_wdata [15] ), .A2(_03930_ ), .ZN(_04907_ ) );
NAND4_X1 _25686_ ( .A1(_03991_ ), .A2(\wbu.io_in_bits_rd_wdata [15] ), .A3(_03998_ ), .A4(_04011_ ), .ZN(_04908_ ) );
AOI211_X1 _25687_ ( .A(_03859_ ), .B(_04907_ ), .C1(_03932_ ), .C2(_04908_ ), .ZN(_04909_ ) );
OAI21_X1 _25688_ ( .A(_03850_ ), .B1(_04901_ ), .B2(_04909_ ), .ZN(_04910_ ) );
NAND3_X1 _25689_ ( .A1(_04444_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04633_ ), .ZN(_04911_ ) );
OR3_X1 _25690_ ( .A1(_04029_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04317_ ), .ZN(_04912_ ) );
OAI21_X1 _25691_ ( .A(_04303_ ), .B1(_04711_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04913_ ) );
NAND4_X1 _25692_ ( .A1(_04403_ ), .A2(_04025_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04039_ ), .ZN(_04914_ ) );
NAND4_X1 _25693_ ( .A1(_04046_ ), .A2(_04148_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_11098_ ), .ZN(_04915_ ) );
NOR3_X1 _25694_ ( .A1(_04263_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10766_ ), .ZN(_04916_ ) );
OAI21_X1 _25695_ ( .A(_04915_ ), .B1(_04053_ ), .B2(_04916_ ), .ZN(_04917_ ) );
INV_X1 _25696_ ( .A(_04050_ ), .ZN(_04918_ ) );
OR4_X1 _25697_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04123_ ), .A3(_04918_ ), .A4(_10766_ ), .ZN(_04919_ ) );
NAND2_X1 _25698_ ( .A1(_04917_ ), .A2(_04919_ ), .ZN(_04920_ ) );
OAI21_X1 _25699_ ( .A(_04914_ ), .B1(_04920_ ), .B2(_04068_ ), .ZN(_04921_ ) );
INV_X1 _25700_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04922_ ) );
NAND4_X1 _25701_ ( .A1(_04073_ ), .A2(_04403_ ), .A3(_04922_ ), .A4(_04399_ ), .ZN(_04923_ ) );
OR2_X1 _25702_ ( .A1(_04272_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04924_ ) );
AND3_X1 _25703_ ( .A1(_04921_ ), .A2(_04923_ ), .A3(_04924_ ), .ZN(_04925_ ) );
MUX2_X1 _25704_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_04925_ ), .S(_04085_ ), .Z(_04926_ ) );
OR3_X1 _25705_ ( .A1(_04592_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04017_ ), .ZN(_04927_ ) );
OR2_X1 _25706_ ( .A1(_04093_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04928_ ) );
AND3_X1 _25707_ ( .A1(_04926_ ), .A2(_04927_ ), .A3(_04928_ ), .ZN(_04929_ ) );
INV_X1 _25708_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04930_ ) );
NAND4_X1 _25709_ ( .A1(_04509_ ), .A2(_04169_ ), .A3(_04930_ ), .A4(_04043_ ), .ZN(_04931_ ) );
INV_X1 _25710_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04932_ ) );
NAND4_X1 _25711_ ( .A1(_04509_ ), .A2(_04146_ ), .A3(_04932_ ), .A4(_04113_ ), .ZN(_04933_ ) );
AND3_X1 _25712_ ( .A1(_04929_ ), .A2(_04931_ ), .A3(_04933_ ), .ZN(_04934_ ) );
OR2_X1 _25713_ ( .A1(_04414_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04935_ ) );
BUF_X2 _25714_ ( .A(_04385_ ), .Z(_04936_ ) );
INV_X1 _25715_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04937_ ) );
NAND4_X1 _25716_ ( .A1(_04936_ ), .A2(_04522_ ), .A3(_04937_ ), .A4(_04189_ ), .ZN(_04938_ ) );
NAND3_X1 _25717_ ( .A1(_04934_ ), .A2(_04935_ ), .A3(_04938_ ), .ZN(_04939_ ) );
INV_X1 _25718_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04940_ ) );
AND4_X1 _25719_ ( .A1(_04940_ ), .A2(_04119_ ), .A3(_04522_ ), .A4(_04189_ ), .ZN(_04941_ ) );
NAND2_X1 _25720_ ( .A1(_04144_ ), .A2(_04032_ ), .ZN(_04942_ ) );
BUF_X2 _25721_ ( .A(_04942_ ), .Z(_04943_ ) );
NOR3_X1 _25722_ ( .A1(_04943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04254_ ), .ZN(_04944_ ) );
NOR3_X1 _25723_ ( .A1(_04939_ ), .A2(_04941_ ), .A3(_04944_ ), .ZN(_04945_ ) );
BUF_X2 _25724_ ( .A(_04918_ ), .Z(_04946_ ) );
BUF_X2 _25725_ ( .A(_04946_ ), .Z(_04947_ ) );
OR3_X1 _25726_ ( .A1(_04029_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04947_ ), .ZN(_04948_ ) );
NAND3_X1 _25727_ ( .A1(_04945_ ), .A2(_04136_ ), .A3(_04948_ ), .ZN(_04949_ ) );
NAND3_X1 _25728_ ( .A1(_04134_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04313_ ), .ZN(_04950_ ) );
AOI21_X1 _25729_ ( .A(_04913_ ), .B1(_04949_ ), .B2(_04950_ ), .ZN(_04951_ ) );
AND3_X1 _25730_ ( .A1(_04062_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04175_ ), .ZN(_04952_ ) );
OAI21_X1 _25731_ ( .A(_04912_ ), .B1(_04951_ ), .B2(_04952_ ), .ZN(_04953_ ) );
INV_X1 _25732_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04954_ ) );
AND3_X1 _25733_ ( .A1(_04162_ ), .A2(_04954_ ), .A3(_04842_ ), .ZN(_04955_ ) );
INV_X1 _25734_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04956_ ) );
AND4_X1 _25735_ ( .A1(_04956_ ), .A2(_04168_ ), .A3(_04171_ ), .A4(_04209_ ), .ZN(_04957_ ) );
NOR3_X1 _25736_ ( .A1(_04953_ ), .A2(_04955_ ), .A3(_04957_ ), .ZN(_04958_ ) );
OR4_X1 _25737_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04179_ ), .A3(_04182_ ), .A4(_04191_ ), .ZN(_04959_ ) );
OR3_X1 _25738_ ( .A1(_04188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04549_ ), .ZN(_04960_ ) );
AND3_X1 _25739_ ( .A1(_04958_ ), .A2(_04959_ ), .A3(_04960_ ), .ZN(_04961_ ) );
INV_X1 _25740_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04962_ ) );
NAND4_X1 _25741_ ( .A1(_04552_ ), .A2(_04553_ ), .A3(_04962_ ), .A4(_04555_ ), .ZN(_04963_ ) );
INV_X1 _25742_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04964_ ) );
NAND4_X1 _25743_ ( .A1(_04620_ ), .A2(_04728_ ), .A3(_04964_ ), .A4(_04211_ ), .ZN(_04965_ ) );
NAND3_X1 _25744_ ( .A1(_04961_ ), .A2(_04963_ ), .A3(_04965_ ), .ZN(_04966_ ) );
OAI21_X1 _25745_ ( .A(_04447_ ), .B1(_04558_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04967_ ) );
OAI21_X1 _25746_ ( .A(_04911_ ), .B1(_04966_ ), .B2(_04967_ ), .ZN(_04968_ ) );
INV_X1 _25747_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04969_ ) );
NAND3_X1 _25748_ ( .A1(_04562_ ), .A2(_04969_ ), .A3(_04224_ ), .ZN(_04970_ ) );
INV_X1 _25749_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04971_ ) );
OAI211_X1 _25750_ ( .A(_04562_ ), .B(_10792_ ), .C1(_04971_ ), .C2(_04555_ ), .ZN(_04972_ ) );
AND3_X1 _25751_ ( .A1(_04968_ ), .A2(_04970_ ), .A3(_04972_ ), .ZN(_04973_ ) );
NAND3_X1 _25752_ ( .A1(_04222_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04482_ ), .ZN(_04974_ ) );
NAND2_X1 _25753_ ( .A1(_04481_ ), .A2(_04974_ ), .ZN(_04975_ ) );
OAI21_X1 _25754_ ( .A(_04910_ ), .B1(_04973_ ), .B2(_04975_ ), .ZN(\idu.io_out_bits_rs1_data [15] ) );
AOI21_X1 _25755_ ( .A(_04738_ ), .B1(_02471_ ), .B2(_02472_ ), .ZN(_04976_ ) );
INV_X1 _25756_ ( .A(_03899_ ), .ZN(_04977_ ) );
OR4_X1 _25757_ ( .A1(_10988_ ), .A2(_00967_ ), .A3(lsu_io_out_bits_rd_wdata_$_MUX__Y_17_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A4(_00969_ ), .ZN(_04978_ ) );
OAI211_X1 _25758_ ( .A(fanout_net_1 ), .B(\io_master_rdata [14] ), .C1(_04463_ ), .C2(_04464_ ), .ZN(_04979_ ) );
AND2_X1 _25759_ ( .A1(_04978_ ), .A2(_04979_ ), .ZN(_04980_ ) );
AOI21_X1 _25760_ ( .A(_10989_ ), .B1(_04751_ ), .B2(_11886_ ), .ZN(_04981_ ) );
CLKBUF_X2 _25761_ ( .A(_04743_ ), .Z(_04982_ ) );
CLKBUF_X2 _25762_ ( .A(_04749_ ), .Z(_04983_ ) );
NAND4_X1 _25763_ ( .A1(_04982_ ), .A2(_04983_ ), .A3(fanout_net_1 ), .A4(lsu_io_out_bits_rd_wdata_$_MUX__Y_9_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .ZN(_04984_ ) );
NAND3_X1 _25764_ ( .A1(_04981_ ), .A2(_03872_ ), .A3(_04984_ ), .ZN(_04985_ ) );
AOI221_X4 _25765_ ( .A(_03883_ ), .B1(_08542_ ), .B2(_03880_ ), .C1(_04346_ ), .C2(_03905_ ), .ZN(_04986_ ) );
AOI221_X4 _25766_ ( .A(_04903_ ), .B1(_04977_ ), .B2(_04980_ ), .C1(_04985_ ), .C2(_04986_ ), .ZN(_04987_ ) );
AOI211_X1 _25767_ ( .A(_03926_ ), .B(_04987_ ), .C1(_03915_ ), .C2(\lsu.io_in_bits_lb ), .ZN(_04988_ ) );
NOR2_X1 _25768_ ( .A1(\lsu.io_in_bits_ren ), .A2(\lsu.io_in_bits_rd_wdata [14] ), .ZN(_04989_ ) );
OR3_X1 _25769_ ( .A1(_04988_ ), .A2(_03930_ ), .A3(_04989_ ), .ZN(_04990_ ) );
OAI211_X1 _25770_ ( .A(\wbu.io_in_bits_rd_wdata [14] ), .B(_04656_ ), .C1(_04657_ ), .C2(_04658_ ), .ZN(_04991_ ) );
AOI21_X1 _25771_ ( .A(_04356_ ), .B1(_04990_ ), .B2(_04991_ ), .ZN(_04992_ ) );
OAI21_X1 _25772_ ( .A(_03851_ ), .B1(_04976_ ), .B2(_04992_ ), .ZN(_04993_ ) );
NAND3_X1 _25773_ ( .A1(_04222_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04482_ ), .ZN(_04994_ ) );
NAND3_X1 _25774_ ( .A1(_04162_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04623_ ), .ZN(_04995_ ) );
AND3_X1 _25775_ ( .A1(_04082_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04411_ ), .ZN(_04996_ ) );
INV_X1 _25776_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04997_ ) );
AND4_X1 _25777_ ( .A1(_04997_ ), .A2(_04107_ ), .A3(_04154_ ), .A4(_04080_ ), .ZN(_04998_ ) );
NAND4_X1 _25778_ ( .A1(_04116_ ), .A2(_04148_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04399_ ), .ZN(_04999_ ) );
NOR3_X1 _25779_ ( .A1(_04294_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_03992_ ), .ZN(_05000_ ) );
OAI21_X1 _25780_ ( .A(_04999_ ), .B1(_04053_ ), .B2(_05000_ ), .ZN(_05001_ ) );
OAI211_X1 _25781_ ( .A(_05001_ ), .B(_04497_ ), .C1(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_04064_ ), .ZN(_05002_ ) );
NAND4_X1 _25782_ ( .A1(_04858_ ), .A2(_04026_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04041_ ), .ZN(_05003_ ) );
AOI21_X1 _25783_ ( .A(_04998_ ), .B1(_05002_ ), .B2(_05003_ ), .ZN(_05004_ ) );
NOR2_X1 _25784_ ( .A1(_04272_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05005_ ) );
NOR2_X1 _25785_ ( .A1(_05005_ ), .A2(_04083_ ), .ZN(_05006_ ) );
AOI21_X1 _25786_ ( .A(_04996_ ), .B1(_05004_ ), .B2(_05006_ ), .ZN(_05007_ ) );
INV_X1 _25787_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05008_ ) );
AND3_X1 _25788_ ( .A1(_04257_ ), .A2(_05008_ ), .A3(_04037_ ), .ZN(_05009_ ) );
NAND2_X1 _25789_ ( .A1(_04057_ ), .A2(_04045_ ), .ZN(_05010_ ) );
BUF_X2 _25790_ ( .A(_05010_ ), .Z(_05011_ ) );
NOR3_X1 _25791_ ( .A1(_05011_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04138_ ), .ZN(_05012_ ) );
NOR3_X1 _25792_ ( .A1(_05007_ ), .A2(_05009_ ), .A3(_05012_ ), .ZN(_05013_ ) );
INV_X1 _25793_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05014_ ) );
NAND4_X1 _25794_ ( .A1(_04509_ ), .A2(_04169_ ), .A3(_05014_ ), .A4(_04113_ ), .ZN(_05015_ ) );
OR2_X1 _25795_ ( .A1(_04102_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05016_ ) );
NAND3_X1 _25796_ ( .A1(_05013_ ), .A2(_05015_ ), .A3(_05016_ ), .ZN(_05017_ ) );
NOR2_X1 _25797_ ( .A1(_04414_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05018_ ) );
CLKBUF_X2 _25798_ ( .A(_04703_ ), .Z(_05019_ ) );
OAI21_X1 _25799_ ( .A(_05019_ ), .B1(_04704_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05020_ ) );
NOR3_X1 _25800_ ( .A1(_05017_ ), .A2(_05018_ ), .A3(_05020_ ), .ZN(_05021_ ) );
AND3_X1 _25801_ ( .A1(_04606_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04169_ ), .ZN(_05022_ ) );
NOR2_X1 _25802_ ( .A1(_05021_ ), .A2(_05022_ ), .ZN(_05023_ ) );
INV_X1 _25803_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05024_ ) );
AND4_X1 _25804_ ( .A1(_05024_ ), .A2(_04147_ ), .A3(_04111_ ), .A4(_04189_ ), .ZN(_05025_ ) );
NOR3_X1 _25805_ ( .A1(_04131_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04946_ ), .ZN(_05026_ ) );
NOR3_X1 _25806_ ( .A1(_05023_ ), .A2(_05025_ ), .A3(_05026_ ), .ZN(_05027_ ) );
INV_X1 _25807_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05028_ ) );
NAND4_X1 _25808_ ( .A1(_04216_ ), .A2(_04525_ ), .A3(_05028_ ), .A4(_04208_ ), .ZN(_05029_ ) );
INV_X1 _25809_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05030_ ) );
NAND4_X1 _25810_ ( .A1(_04297_ ), .A2(_04151_ ), .A3(_05030_ ), .A4(_04208_ ), .ZN(_05031_ ) );
AND3_X1 _25811_ ( .A1(_05027_ ), .A2(_05029_ ), .A3(_05031_ ), .ZN(_05032_ ) );
OAI21_X1 _25812_ ( .A(_05032_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04303_ ), .ZN(_05033_ ) );
OAI21_X1 _25813_ ( .A(_04165_ ), .B1(_04428_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05034_ ) );
OAI21_X1 _25814_ ( .A(_04995_ ), .B1(_05033_ ), .B2(_05034_ ), .ZN(_05035_ ) );
INV_X1 _25815_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05036_ ) );
NAND4_X1 _25816_ ( .A1(_04536_ ), .A2(_04615_ ), .A3(_05036_ ), .A4(_04210_ ), .ZN(_05037_ ) );
AND2_X1 _25817_ ( .A1(_04082_ ), .A2(_04310_ ), .ZN(_05038_ ) );
INV_X1 _25818_ ( .A(_05038_ ), .ZN(_05039_ ) );
OR2_X1 _25819_ ( .A1(_05039_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05040_ ) );
AND3_X1 _25820_ ( .A1(_05035_ ), .A2(_05037_ ), .A3(_05040_ ), .ZN(_05041_ ) );
OR3_X1 _25821_ ( .A1(_04548_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04550_ ), .ZN(_05042_ ) );
INV_X1 _25822_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05043_ ) );
NAND4_X1 _25823_ ( .A1(_04552_ ), .A2(_04553_ ), .A3(_05043_ ), .A4(_04555_ ), .ZN(_05044_ ) );
NAND3_X1 _25824_ ( .A1(_05041_ ), .A2(_05042_ ), .A3(_05044_ ), .ZN(_05045_ ) );
INV_X1 _25825_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05046_ ) );
AND4_X1 _25826_ ( .A1(_05046_ ), .A2(_04620_ ), .A3(_04728_ ), .A4(_04624_ ), .ZN(_05047_ ) );
NOR2_X1 _25827_ ( .A1(_04558_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05048_ ) );
NOR3_X1 _25828_ ( .A1(_05045_ ), .A2(_05047_ ), .A3(_05048_ ), .ZN(_05049_ ) );
OR3_X1 _25829_ ( .A1(_04030_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04034_ ), .ZN(_05050_ ) );
INV_X1 _25830_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05051_ ) );
NAND3_X1 _25831_ ( .A1(_04562_ ), .A2(_05051_ ), .A3(_04224_ ), .ZN(_05052_ ) );
NAND3_X1 _25832_ ( .A1(_05049_ ), .A2(_05050_ ), .A3(_05052_ ), .ZN(_05053_ ) );
AOI211_X1 _25833_ ( .A(_04566_ ), .B(_04567_ ), .C1(_04568_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05054_ ) );
OAI211_X1 _25834_ ( .A(_04481_ ), .B(_04994_ ), .C1(_05053_ ), .C2(_05054_ ), .ZN(_05055_ ) );
NAND2_X1 _25835_ ( .A1(_04993_ ), .A2(_05055_ ), .ZN(\idu.io_out_bits_rs1_data [14] ) );
NOR2_X1 _25836_ ( .A1(_04988_ ), .A2(_04989_ ), .ZN(\lsu.io_out_bits_rd_wdata [14] ) );
NAND2_X1 _25837_ ( .A1(\exu.io_out_bits_rd_wdata [13] ), .A2(_04356_ ), .ZN(_05056_ ) );
OR4_X1 _25838_ ( .A1(_10988_ ), .A2(_00967_ ), .A3(lsu_io_out_bits_rd_wdata_$_MUX__Y_18_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A4(_00969_ ), .ZN(_05057_ ) );
OAI211_X1 _25839_ ( .A(fanout_net_1 ), .B(\io_master_rdata [13] ), .C1(_04463_ ), .C2(_04464_ ), .ZN(_05058_ ) );
AND2_X1 _25840_ ( .A1(_05057_ ), .A2(_05058_ ), .ZN(_05059_ ) );
OR3_X1 _25841_ ( .A1(_04360_ ), .A2(_10990_ ), .A3(\io_master_awaddr [1] ), .ZN(_05060_ ) );
AOI221_X4 _25842_ ( .A(_03883_ ), .B1(_08542_ ), .B2(_03880_ ), .C1(_04366_ ), .C2(_03905_ ), .ZN(_05061_ ) );
AOI221_X4 _25843_ ( .A(_04903_ ), .B1(_04977_ ), .B2(_05059_ ), .C1(_05060_ ), .C2(_05061_ ), .ZN(_05062_ ) );
AOI211_X1 _25844_ ( .A(_03927_ ), .B(_05062_ ), .C1(_03915_ ), .C2(\lsu.io_in_bits_lb ), .ZN(_05063_ ) );
NOR2_X1 _25845_ ( .A1(\lsu.io_in_bits_ren ), .A2(\lsu.io_in_bits_rd_wdata [13] ), .ZN(_05064_ ) );
NOR3_X1 _25846_ ( .A1(_05063_ ), .A2(_03930_ ), .A3(_05064_ ), .ZN(_05065_ ) );
NOR3_X1 _25847_ ( .A1(_04340_ ), .A2(_13629_ ), .A3(_04341_ ), .ZN(_05066_ ) );
OAI21_X1 _25848_ ( .A(_04738_ ), .B1(_05065_ ), .B2(_05066_ ), .ZN(_05067_ ) );
AOI21_X1 _25849_ ( .A(\idu.rs_reg ), .B1(_05056_ ), .B2(_05067_ ), .ZN(_05068_ ) );
INV_X1 _25850_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05069_ ) );
NAND3_X1 _25851_ ( .A1(_04078_ ), .A2(_05069_ ), .A3(_11100_ ), .ZN(_05070_ ) );
INV_X1 _25852_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05071_ ) );
NAND3_X1 _25853_ ( .A1(_04051_ ), .A2(_05071_ ), .A3(_04039_ ), .ZN(_05072_ ) );
OAI21_X1 _25854_ ( .A(_05072_ ), .B1(_04493_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_05073_ ) );
NOR2_X1 _25855_ ( .A1(_04070_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05074_ ) );
INV_X1 _25856_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05075_ ) );
AND4_X1 _25857_ ( .A1(_05075_ ), .A2(_04098_ ), .A3(_04148_ ), .A4(_11098_ ), .ZN(_05076_ ) );
NOR4_X1 _25858_ ( .A1(_05073_ ), .A2(_05074_ ), .A3(_04395_ ), .A4(_05076_ ), .ZN(_05077_ ) );
AND4_X1 _25859_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04073_ ), .A3(_04403_ ), .A4(_04399_ ), .ZN(_05078_ ) );
OAI21_X1 _25860_ ( .A(_05070_ ), .B1(_05077_ ), .B2(_05078_ ), .ZN(_05079_ ) );
NOR4_X1 _25861_ ( .A1(_04124_ ), .A2(_04180_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04016_ ), .ZN(_05080_ ) );
NOR3_X1 _25862_ ( .A1(_04186_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03993_ ), .ZN(_05081_ ) );
NOR3_X1 _25863_ ( .A1(_05079_ ), .A2(_05080_ ), .A3(_05081_ ), .ZN(_05082_ ) );
INV_X1 _25864_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05083_ ) );
NAND3_X1 _25865_ ( .A1(_04257_ ), .A2(_05083_ ), .A3(_04108_ ), .ZN(_05084_ ) );
OR3_X1 _25866_ ( .A1(_04095_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04127_ ), .ZN(_05085_ ) );
NAND3_X1 _25867_ ( .A1(_05082_ ), .A2(_05084_ ), .A3(_05085_ ), .ZN(_05086_ ) );
NOR2_X1 _25868_ ( .A1(_04102_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05087_ ) );
NAND2_X1 _25869_ ( .A1(_04031_ ), .A2(_04026_ ), .ZN(_05088_ ) );
NOR3_X1 _25870_ ( .A1(_05088_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04138_ ), .ZN(_05089_ ) );
NOR3_X1 _25871_ ( .A1(_05086_ ), .A2(_05087_ ), .A3(_05089_ ), .ZN(_05090_ ) );
INV_X1 _25872_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05091_ ) );
NAND4_X1 _25873_ ( .A1(_04385_ ), .A2(_04036_ ), .A3(_05091_ ), .A4(_04283_ ), .ZN(_05092_ ) );
OR2_X1 _25874_ ( .A1(_05019_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05093_ ) );
NAND3_X1 _25875_ ( .A1(_05090_ ), .A2(_05092_ ), .A3(_05093_ ), .ZN(_05094_ ) );
INV_X1 _25876_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05095_ ) );
AND4_X1 _25877_ ( .A1(_05095_ ), .A2(_04146_ ), .A3(_04110_ ), .A4(_04283_ ), .ZN(_05096_ ) );
NOR3_X1 _25878_ ( .A1(_04028_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04918_ ), .ZN(_05097_ ) );
NOR3_X1 _25879_ ( .A1(_05094_ ), .A2(_05096_ ), .A3(_05097_ ), .ZN(_05098_ ) );
INV_X1 _25880_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05099_ ) );
NAND4_X1 _25881_ ( .A1(_04936_ ), .A2(_04253_ ), .A3(_05099_ ), .A4(_04173_ ), .ZN(_05100_ ) );
INV_X1 _25882_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05101_ ) );
NAND4_X1 _25883_ ( .A1(_04119_ ), .A2(_04253_ ), .A3(_05101_ ), .A4(_04173_ ), .ZN(_05102_ ) );
NAND3_X1 _25884_ ( .A1(_05098_ ), .A2(_05100_ ), .A3(_05102_ ), .ZN(_05103_ ) );
NOR4_X1 _25885_ ( .A1(_04126_ ), .A2(_04946_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04189_ ), .ZN(_05104_ ) );
INV_X1 _25886_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05105_ ) );
AND4_X1 _25887_ ( .A1(_05105_ ), .A2(_04155_ ), .A3(_04157_ ), .A4(_04019_ ), .ZN(_05106_ ) );
NOR3_X1 _25888_ ( .A1(_05103_ ), .A2(_05104_ ), .A3(_05106_ ), .ZN(_05107_ ) );
OR2_X1 _25889_ ( .A1(_04165_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05108_ ) );
INV_X1 _25890_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05109_ ) );
NAND4_X1 _25891_ ( .A1(_04167_ ), .A2(_04297_ ), .A3(_05109_ ), .A4(_04174_ ), .ZN(_05110_ ) );
NAND3_X1 _25892_ ( .A1(_05107_ ), .A2(_05108_ ), .A3(_05110_ ), .ZN(_05111_ ) );
NOR4_X1 _25893_ ( .A1(_04178_ ), .A2(_04317_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04183_ ), .ZN(_05112_ ) );
INV_X1 _25894_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05113_ ) );
AND4_X1 _25895_ ( .A1(_05113_ ), .A2(_04332_ ), .A3(_04158_ ), .A4(_04174_ ), .ZN(_05114_ ) );
NOR3_X1 _25896_ ( .A1(_05111_ ), .A2(_05112_ ), .A3(_05114_ ), .ZN(_05115_ ) );
INV_X1 _25897_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05116_ ) );
NAND4_X1 _25898_ ( .A1(_04196_ ), .A2(_04000_ ), .A3(_05116_ ), .A4(_10756_ ), .ZN(_05117_ ) );
INV_X1 _25899_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05118_ ) );
AOI22_X1 _25900_ ( .A1(_04203_ ), .A2(_05118_ ), .B1(_04175_ ), .B2(_04207_ ), .ZN(_05119_ ) );
AND3_X1 _25901_ ( .A1(_05115_ ), .A2(_05117_ ), .A3(_05119_ ), .ZN(_05120_ ) );
AND3_X1 _25902_ ( .A1(_04207_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04842_ ), .ZN(_05121_ ) );
NOR2_X1 _25903_ ( .A1(_05120_ ), .A2(_05121_ ), .ZN(_05122_ ) );
INV_X1 _25904_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05123_ ) );
AND4_X1 _25905_ ( .A1(_05123_ ), .A2(_04445_ ), .A3(_04451_ ), .A4(_04623_ ), .ZN(_05124_ ) );
NOR3_X1 _25906_ ( .A1(_04519_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04327_ ), .ZN(_05125_ ) );
NOR3_X1 _25907_ ( .A1(_05122_ ), .A2(_05124_ ), .A3(_05125_ ), .ZN(_05126_ ) );
NOR4_X1 _25908_ ( .A1(_04023_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04015_ ), .A4(_04199_ ), .ZN(_05127_ ) );
NOR2_X1 _25909_ ( .A1(_05127_ ), .A2(_04249_ ), .ZN(_05128_ ) );
AOI221_X4 _25910_ ( .A(_04240_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B2(_04250_ ), .C1(_05126_ ), .C2(_05128_ ), .ZN(_05129_ ) );
OR2_X1 _25911_ ( .A1(_05068_ ), .A2(_05129_ ), .ZN(\idu.io_out_bits_rs1_data [13] ) );
NOR2_X1 _25912_ ( .A1(_05063_ ), .A2(_05064_ ), .ZN(\lsu.io_out_bits_rd_wdata [13] ) );
NAND2_X1 _25913_ ( .A1(\exu.io_out_bits_rd_wdata [12] ), .A2(_04459_ ), .ZN(_05130_ ) );
NAND2_X1 _25914_ ( .A1(_04470_ ), .A2(_04471_ ), .ZN(_05131_ ) );
AND3_X1 _25915_ ( .A1(_05131_ ), .A2(fanout_net_1 ), .A3(_04469_ ), .ZN(_05132_ ) );
NOR3_X1 _25916_ ( .A1(_04466_ ), .A2(_10990_ ), .A3(\io_master_awaddr [1] ), .ZN(_05133_ ) );
OAI211_X1 _25917_ ( .A(_03910_ ), .B(_03909_ ), .C1(_05132_ ), .C2(_05133_ ), .ZN(_05134_ ) );
INV_X1 _25918_ ( .A(_05134_ ), .ZN(_05135_ ) );
OR4_X1 _25919_ ( .A1(_10989_ ), .A2(_04463_ ), .A3(lsu_io_out_bits_rd_wdata_$_MUX__Y_19_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A4(_04464_ ), .ZN(_05136_ ) );
OAI211_X1 _25920_ ( .A(fanout_net_1 ), .B(\io_master_rdata [12] ), .C1(_00968_ ), .C2(_00970_ ), .ZN(_05137_ ) );
AOI22_X1 _25921_ ( .A1(_03909_ ), .A2(_03910_ ), .B1(_05136_ ), .B2(_05137_ ), .ZN(_05138_ ) );
OAI21_X1 _25922_ ( .A(_04904_ ), .B1(_05135_ ), .B2(_05138_ ), .ZN(_05139_ ) );
AND3_X1 _25923_ ( .A1(_04358_ ), .A2(\lsu.io_in_bits_ren ), .A3(_05139_ ), .ZN(_05140_ ) );
NOR2_X1 _25924_ ( .A1(\lsu.io_in_bits_ren ), .A2(\lsu.io_in_bits_rd_wdata [12] ), .ZN(_05141_ ) );
OAI21_X1 _25925_ ( .A(_04340_ ), .B1(_05140_ ), .B2(_05141_ ), .ZN(_05142_ ) );
AND4_X1 _25926_ ( .A1(\wbu.io_in_bits_rd_wdata [12] ), .A2(_03990_ ), .A3(_03997_ ), .A4(_04010_ ), .ZN(_05143_ ) );
OAI211_X1 _25927_ ( .A(_05142_ ), .B(_03856_ ), .C1(_04353_ ), .C2(_05143_ ), .ZN(_05144_ ) );
AOI21_X1 _25928_ ( .A(\idu.rs_reg ), .B1(_05130_ ), .B2(_05144_ ), .ZN(_05145_ ) );
AND3_X1 _25929_ ( .A1(_04221_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04242_ ), .ZN(_05146_ ) );
INV_X1 _25930_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_05147_ ) );
NAND3_X1 _25931_ ( .A1(_04058_ ), .A2(_05147_ ), .A3(_11098_ ), .ZN(_05148_ ) );
OAI21_X1 _25932_ ( .A(_05148_ ), .B1(_04054_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05149_ ) );
INV_X1 _25933_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05150_ ) );
AOI21_X1 _25934_ ( .A(_05149_ ), .B1(_05150_ ), .B2(_04392_ ), .ZN(_05151_ ) );
OR2_X1 _25935_ ( .A1(_04069_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05152_ ) );
INV_X1 _25936_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05153_ ) );
AOI22_X1 _25937_ ( .A1(_04395_ ), .A2(_05153_ ), .B1(_04039_ ), .B2(_04077_ ), .ZN(_05154_ ) );
AND3_X1 _25938_ ( .A1(_05151_ ), .A2(_05152_ ), .A3(_05154_ ), .ZN(_05155_ ) );
AND3_X1 _25939_ ( .A1(_04077_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04399_ ), .ZN(_05156_ ) );
NOR2_X1 _25940_ ( .A1(_05155_ ), .A2(_05156_ ), .ZN(_05157_ ) );
INV_X1 _25941_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05158_ ) );
AND4_X1 _25942_ ( .A1(_05158_ ), .A2(_04098_ ), .A3(_04403_ ), .A4(_04399_ ), .ZN(_05159_ ) );
NOR3_X1 _25943_ ( .A1(_04186_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03993_ ), .ZN(_05160_ ) );
NOR3_X1 _25944_ ( .A1(_05157_ ), .A2(_05159_ ), .A3(_05160_ ), .ZN(_05161_ ) );
INV_X1 _25945_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05162_ ) );
NAND3_X1 _25946_ ( .A1(_04257_ ), .A2(_05162_ ), .A3(_04384_ ), .ZN(_05163_ ) );
INV_X1 _25947_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05164_ ) );
NAND4_X1 _25948_ ( .A1(_04331_ ), .A2(_04117_ ), .A3(_05164_ ), .A4(_04411_ ), .ZN(_05165_ ) );
NAND3_X1 _25949_ ( .A1(_05161_ ), .A2(_05163_ ), .A3(_05165_ ), .ZN(_05166_ ) );
NOR2_X1 _25950_ ( .A1(_04102_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05167_ ) );
NOR3_X1 _25951_ ( .A1(_05088_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04017_ ), .ZN(_05168_ ) );
NOR3_X1 _25952_ ( .A1(_05166_ ), .A2(_05167_ ), .A3(_05168_ ), .ZN(_05169_ ) );
OR3_X1 _25953_ ( .A1(_04518_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03994_ ), .ZN(_05170_ ) );
OR2_X1 _25954_ ( .A1(_05019_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05171_ ) );
NAND3_X1 _25955_ ( .A1(_05169_ ), .A2(_05170_ ), .A3(_05171_ ), .ZN(_05172_ ) );
INV_X1 _25956_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05173_ ) );
AND4_X1 _25957_ ( .A1(_05173_ ), .A2(_04145_ ), .A3(_04110_ ), .A4(_04598_ ), .ZN(_05174_ ) );
INV_X1 _25958_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05175_ ) );
AND4_X1 _25959_ ( .A1(_05175_ ), .A2(_04149_ ), .A3(_04037_ ), .A4(_04128_ ), .ZN(_05176_ ) );
NOR3_X1 _25960_ ( .A1(_05172_ ), .A2(_05174_ ), .A3(_05176_ ), .ZN(_05177_ ) );
OR3_X1 _25961_ ( .A1(_04294_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04113_ ), .ZN(_05178_ ) );
INV_X1 _25962_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05179_ ) );
NAND4_X1 _25963_ ( .A1(_04119_ ), .A2(_04150_ ), .A3(_05179_ ), .A4(_04129_ ), .ZN(_05180_ ) );
NAND3_X1 _25964_ ( .A1(_05177_ ), .A2(_05178_ ), .A3(_05180_ ), .ZN(_05181_ ) );
INV_X1 _25965_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05182_ ) );
AND4_X1 _25966_ ( .A1(_05182_ ), .A2(_04146_ ), .A3(_04150_ ), .A4(_04129_ ), .ZN(_05183_ ) );
NOR3_X1 _25967_ ( .A1(_04131_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04180_ ), .ZN(_05184_ ) );
NOR3_X1 _25968_ ( .A1(_05181_ ), .A2(_05183_ ), .A3(_05184_ ), .ZN(_05185_ ) );
OR2_X1 _25969_ ( .A1(_04165_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05186_ ) );
INV_X1 _25970_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05187_ ) );
NAND4_X1 _25971_ ( .A1(_04156_ ), .A2(_04170_ ), .A3(_05187_ ), .A4(_04020_ ), .ZN(_05188_ ) );
NAND3_X1 _25972_ ( .A1(_05185_ ), .A2(_05186_ ), .A3(_05188_ ), .ZN(_05189_ ) );
NOR4_X1 _25973_ ( .A1(_04178_ ), .A2(_04181_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04183_ ), .ZN(_05190_ ) );
INV_X1 _25974_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05191_ ) );
AND4_X1 _25975_ ( .A1(_05191_ ), .A2(_04332_ ), .A3(_04157_ ), .A4(_04159_ ), .ZN(_05192_ ) );
NOR3_X1 _25976_ ( .A1(_05189_ ), .A2(_05190_ ), .A3(_05192_ ), .ZN(_05193_ ) );
INV_X1 _25977_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05194_ ) );
NAND4_X1 _25978_ ( .A1(_04196_ ), .A2(_04000_ ), .A3(_05194_ ), .A4(_10756_ ), .ZN(_05195_ ) );
NAND3_X1 _25979_ ( .A1(_05193_ ), .A2(_04204_ ), .A3(_05195_ ), .ZN(_05196_ ) );
NAND3_X1 _25980_ ( .A1(_04048_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04842_ ), .ZN(_05197_ ) );
AOI21_X1 _25981_ ( .A(_04201_ ), .B1(_05196_ ), .B2(_05197_ ), .ZN(_05198_ ) );
AND4_X1 _25982_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04332_ ), .A3(_04241_ ), .A4(_04842_ ), .ZN(_05199_ ) );
NOR2_X1 _25983_ ( .A1(_05198_ ), .A2(_05199_ ), .ZN(_05200_ ) );
CLKBUF_X2 _25984_ ( .A(_05088_ ), .Z(_05201_ ) );
BUF_X2 _25985_ ( .A(_05201_ ), .Z(_05202_ ) );
NOR3_X1 _25986_ ( .A1(_05202_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04327_ ), .ZN(_05203_ ) );
NOR3_X1 _25987_ ( .A1(_04519_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04327_ ), .ZN(_05204_ ) );
NOR3_X1 _25988_ ( .A1(_05200_ ), .A2(_05203_ ), .A3(_05204_ ), .ZN(_05205_ ) );
AND2_X1 _25989_ ( .A1(_04021_ ), .A2(_04528_ ), .ZN(_05206_ ) );
INV_X1 _25990_ ( .A(_05206_ ), .ZN(_05207_ ) );
MUX2_X1 _25991_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B(_05205_ ), .S(_05207_ ), .Z(_05208_ ) );
AOI211_X1 _25992_ ( .A(_04240_ ), .B(_05146_ ), .C1(_05208_ ), .C2(_04251_ ), .ZN(_05209_ ) );
OR2_X1 _25993_ ( .A1(_05145_ ), .A2(_05209_ ), .ZN(\idu.io_out_bits_rs1_data [12] ) );
NOR2_X1 _25994_ ( .A1(_05140_ ), .A2(_05141_ ), .ZN(\lsu.io_out_bits_rd_wdata [12] ) );
NOR2_X1 _25995_ ( .A1(_02660_ ), .A2(_03857_ ), .ZN(_05210_ ) );
NOR3_X1 _25996_ ( .A1(_03899_ ), .A2(_03900_ ), .A3(_04367_ ), .ZN(_05211_ ) );
OR2_X1 _25997_ ( .A1(_03898_ ), .A2(_05211_ ), .ZN(_05212_ ) );
OAI21_X1 _25998_ ( .A(\lsu.io_in_bits_ren ), .B1(_05212_ ), .B2(_03917_ ), .ZN(_05213_ ) );
NAND2_X1 _25999_ ( .A1(_03927_ ), .A2(\lsu.io_in_bits_rd_wdata [29] ), .ZN(_05214_ ) );
AND3_X1 _26000_ ( .A1(_05213_ ), .A2(_03925_ ), .A3(_05214_ ), .ZN(_05215_ ) );
NAND4_X1 _26001_ ( .A1(_03991_ ), .A2(\wbu.io_in_bits_rd_wdata [29] ), .A3(_03998_ ), .A4(_04011_ ), .ZN(_05216_ ) );
AOI211_X1 _26002_ ( .A(_03859_ ), .B(_05215_ ), .C1(_03932_ ), .C2(_05216_ ), .ZN(_05217_ ) );
OAI21_X1 _26003_ ( .A(_03850_ ), .B1(_05210_ ), .B2(_05217_ ), .ZN(_05218_ ) );
OAI21_X1 _26004_ ( .A(_04447_ ), .B1(_04558_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05219_ ) );
AND3_X1 _26005_ ( .A1(_04104_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04026_ ), .ZN(_05220_ ) );
NAND3_X1 _26006_ ( .A1(_04088_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04025_ ), .ZN(_05221_ ) );
AND4_X1 _26007_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04066_ ), .A3(_04025_ ), .A4(_11097_ ), .ZN(_05222_ ) );
OR3_X1 _26008_ ( .A1(_04262_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10605_ ), .ZN(_05223_ ) );
MUX2_X1 _26009_ ( .A(_05223_ ), .B(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(_04052_ ), .Z(_05224_ ) );
MUX2_X1 _26010_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_05224_ ), .S(_04064_ ), .Z(_05225_ ) );
AOI21_X1 _26011_ ( .A(_05222_ ), .B1(_05225_ ), .B2(_04069_ ), .ZN(_05226_ ) );
INV_X1 _26012_ ( .A(_04162_ ), .ZN(_05227_ ) );
AOI211_X1 _26013_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_05227_ ), .C1(\idu.io_in_bits_inst [19] ), .C2(_10646_ ), .ZN(_05228_ ) );
INV_X1 _26014_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05229_ ) );
AND4_X1 _26015_ ( .A1(_05229_ ), .A2(_04074_ ), .A3(_04046_ ), .A4(_11097_ ), .ZN(_05230_ ) );
OR3_X1 _26016_ ( .A1(_05226_ ), .A2(_05228_ ), .A3(_05230_ ), .ZN(_05231_ ) );
OAI21_X1 _26017_ ( .A(_04090_ ), .B1(_04085_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05232_ ) );
OAI21_X1 _26018_ ( .A(_05221_ ), .B1(_05231_ ), .B2(_05232_ ), .ZN(_05233_ ) );
OR3_X1 _26019_ ( .A1(_05010_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03992_ ), .ZN(_05234_ ) );
INV_X1 _26020_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05235_ ) );
NAND4_X1 _26021_ ( .A1(_04045_ ), .A2(_04116_ ), .A3(_05235_ ), .A4(_04040_ ), .ZN(_05236_ ) );
AND3_X1 _26022_ ( .A1(_05233_ ), .A2(_05234_ ), .A3(_05236_ ), .ZN(_05237_ ) );
INV_X1 _26023_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05238_ ) );
AOI22_X1 _26024_ ( .A1(_04100_ ), .A2(_05238_ ), .B1(_04026_ ), .B2(_04104_ ), .ZN(_05239_ ) );
AOI21_X1 _26025_ ( .A(_05220_ ), .B1(_05237_ ), .B2(_05239_ ), .ZN(_05240_ ) );
INV_X1 _26026_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05241_ ) );
AND4_X1 _26027_ ( .A1(_05241_ ), .A2(_04384_ ), .A3(_04032_ ), .A4(_04411_ ), .ZN(_05242_ ) );
INV_X1 _26028_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05243_ ) );
AND4_X1 _26029_ ( .A1(_05243_ ), .A2(_04116_ ), .A3(_04032_ ), .A4(_04411_ ), .ZN(_05244_ ) );
NOR3_X1 _26030_ ( .A1(_05240_ ), .A2(_05242_ ), .A3(_05244_ ), .ZN(_05245_ ) );
OR3_X1 _26031_ ( .A1(_04942_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03994_ ), .ZN(_05246_ ) );
OR3_X1 _26032_ ( .A1(_04028_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04918_ ), .ZN(_05247_ ) );
NAND3_X1 _26033_ ( .A1(_05245_ ), .A2(_05246_ ), .A3(_05247_ ), .ZN(_05248_ ) );
INV_X1 _26034_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05249_ ) );
AND4_X1 _26035_ ( .A1(_05249_ ), .A2(_04385_ ), .A3(_04149_ ), .A4(_04128_ ), .ZN(_05250_ ) );
INV_X1 _26036_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05251_ ) );
AND4_X1 _26037_ ( .A1(_05251_ ), .A2(_04117_ ), .A3(_04149_ ), .A4(_04128_ ), .ZN(_05252_ ) );
NOR3_X1 _26038_ ( .A1(_05248_ ), .A2(_05250_ ), .A3(_05252_ ), .ZN(_05253_ ) );
MUX2_X1 _26039_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_05253_ ), .S(_04302_ ), .Z(_05254_ ) );
MUX2_X1 _26040_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_05254_ ), .S(_04428_ ), .Z(_05255_ ) );
INV_X1 _26041_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05256_ ) );
NAND4_X1 _26042_ ( .A1(_04217_ ), .A2(_04168_ ), .A3(_05256_ ), .A4(_04209_ ), .ZN(_05257_ ) );
OR2_X1 _26043_ ( .A1(_04435_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05258_ ) );
AND3_X1 _26044_ ( .A1(_05255_ ), .A2(_05257_ ), .A3(_05258_ ), .ZN(_05259_ ) );
OR4_X1 _26045_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04316_ ), .A3(_04182_ ), .A4(_04184_ ), .ZN(_05260_ ) );
OR3_X1 _26046_ ( .A1(_04188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04191_ ), .ZN(_05261_ ) );
AND3_X1 _26047_ ( .A1(_05259_ ), .A2(_05260_ ), .A3(_05261_ ), .ZN(_05262_ ) );
INV_X1 _26048_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05263_ ) );
NAND4_X1 _26049_ ( .A1(_04197_ ), .A2(_04194_ ), .A3(_05263_ ), .A4(_04199_ ), .ZN(_05264_ ) );
NAND3_X1 _26050_ ( .A1(_05262_ ), .A2(_04204_ ), .A3(_05264_ ), .ZN(_05265_ ) );
NAND3_X1 _26051_ ( .A1(_04048_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04211_ ), .ZN(_05266_ ) );
AOI21_X1 _26052_ ( .A(_05219_ ), .B1(_05265_ ), .B2(_05266_ ), .ZN(_05267_ ) );
AND3_X1 _26053_ ( .A1(_04444_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04633_ ), .ZN(_05268_ ) );
OAI221_X1 _26054_ ( .A(_05207_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04219_ ), .C1(_05267_ ), .C2(_05268_ ), .ZN(_05269_ ) );
NAND3_X1 _26055_ ( .A1(_04222_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04728_ ), .ZN(_05270_ ) );
AOI21_X1 _26056_ ( .A(_04250_ ), .B1(_05269_ ), .B2(_05270_ ), .ZN(_05271_ ) );
INV_X1 _26057_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_05272_ ) );
OAI21_X1 _26058_ ( .A(_04247_ ), .B1(_05272_ ), .B2(_04251_ ), .ZN(_05273_ ) );
OAI21_X1 _26059_ ( .A(_05218_ ), .B1(_05271_ ), .B2(_05273_ ), .ZN(\idu.io_out_bits_rs1_data [29] ) );
NOR3_X1 _26060_ ( .A1(_03925_ ), .A2(_13719_ ), .A3(_04341_ ), .ZN(_05274_ ) );
OR3_X1 _26061_ ( .A1(_04644_ ), .A2(_10990_ ), .A3(\io_master_awaddr [1] ), .ZN(_05275_ ) );
NAND3_X1 _26062_ ( .A1(_04648_ ), .A2(fanout_net_1 ), .A3(_04469_ ), .ZN(_05276_ ) );
NAND3_X1 _26063_ ( .A1(_03899_ ), .A2(_05275_ ), .A3(_05276_ ), .ZN(_05277_ ) );
OR4_X1 _26064_ ( .A1(_10989_ ), .A2(_00968_ ), .A3(lsu_io_out_bits_rd_wdata_$_MUX__Y_20_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A4(_04464_ ), .ZN(_05278_ ) );
OAI211_X1 _26065_ ( .A(fanout_net_1 ), .B(\io_master_rdata [11] ), .C1(_00968_ ), .C2(_00970_ ), .ZN(_05279_ ) );
AND2_X1 _26066_ ( .A1(_05278_ ), .A2(_05279_ ), .ZN(_05280_ ) );
OAI21_X1 _26067_ ( .A(_05280_ ), .B1(_03882_ ), .B2(_03883_ ), .ZN(_05281_ ) );
NAND3_X1 _26068_ ( .A1(_05277_ ), .A2(_04904_ ), .A3(_05281_ ), .ZN(_05282_ ) );
INV_X1 _26069_ ( .A(_03915_ ), .ZN(_05283_ ) );
INV_X1 _26070_ ( .A(\lsu.io_in_bits_lb ), .ZN(_05284_ ) );
OAI211_X1 _26071_ ( .A(\lsu.io_in_bits_ren ), .B(_05282_ ), .C1(_05283_ ), .C2(_05284_ ), .ZN(_05285_ ) );
OR2_X1 _26072_ ( .A1(\lsu.io_in_bits_ren ), .A2(\lsu.io_in_bits_rd_wdata [11] ), .ZN(_05286_ ) );
AND2_X1 _26073_ ( .A1(_05285_ ), .A2(_05286_ ), .ZN(\lsu.io_out_bits_rd_wdata [11] ) );
AOI21_X1 _26074_ ( .A(_05274_ ), .B1(\lsu.io_out_bits_rd_wdata [11] ), .B2(_04353_ ), .ZN(_05287_ ) );
MUX2_X1 _26075_ ( .A(_05287_ ), .B(_02730_ ), .S(_04228_ ), .Z(_05288_ ) );
INV_X1 _26076_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05289_ ) );
INV_X1 _26077_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05290_ ) );
AND3_X1 _26078_ ( .A1(_04088_ ), .A2(_05290_ ), .A3(_04026_ ), .ZN(_05291_ ) );
OR3_X1 _26079_ ( .A1(_04263_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10766_ ), .ZN(_05292_ ) );
BUF_X2 _26080_ ( .A(_04054_ ), .Z(_05293_ ) );
OAI21_X1 _26081_ ( .A(_05292_ ), .B1(_05293_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05294_ ) );
NOR2_X1 _26082_ ( .A1(_04070_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05295_ ) );
INV_X1 _26083_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05296_ ) );
AND4_X1 _26084_ ( .A1(_05296_ ), .A2(_04098_ ), .A3(_04050_ ), .A4(_11098_ ), .ZN(_05297_ ) );
NOR4_X1 _26085_ ( .A1(_05294_ ), .A2(_05295_ ), .A3(_04395_ ), .A4(_05297_ ), .ZN(_05298_ ) );
AND4_X1 _26086_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04073_ ), .A3(_04403_ ), .A4(_11099_ ), .ZN(_05299_ ) );
OAI221_X1 _26087_ ( .A(_04085_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04272_ ), .C1(_05298_ ), .C2(_05299_ ), .ZN(_05300_ ) );
NAND4_X1 _26088_ ( .A1(_04144_ ), .A2(_04154_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_11100_ ), .ZN(_05301_ ) );
AOI21_X1 _26089_ ( .A(_05291_ ), .B1(_05300_ ), .B2(_05301_ ), .ZN(_05302_ ) );
OR3_X1 _26090_ ( .A1(_05011_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03993_ ), .ZN(_05303_ ) );
INV_X1 _26091_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05304_ ) );
NAND4_X1 _26092_ ( .A1(_04331_ ), .A2(_04117_ ), .A3(_05304_ ), .A4(_04282_ ), .ZN(_05305_ ) );
NAND3_X1 _26093_ ( .A1(_05302_ ), .A2(_05303_ ), .A3(_05305_ ), .ZN(_05306_ ) );
NOR2_X1 _26094_ ( .A1(_04102_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05307_ ) );
OAI21_X1 _26095_ ( .A(_04704_ ), .B1(_04414_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05308_ ) );
NOR3_X1 _26096_ ( .A1(_05306_ ), .A2(_05307_ ), .A3(_05308_ ), .ZN(_05309_ ) );
AND3_X1 _26097_ ( .A1(_04287_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04108_ ), .ZN(_05310_ ) );
NOR2_X1 _26098_ ( .A1(_05309_ ), .A2(_05310_ ), .ZN(_05311_ ) );
INV_X1 _26099_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05312_ ) );
AND4_X1 _26100_ ( .A1(_05312_ ), .A2(_04118_ ), .A3(_04110_ ), .A4(_04598_ ), .ZN(_05313_ ) );
NOR3_X1 _26101_ ( .A1(_04943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04163_ ), .ZN(_05314_ ) );
NOR3_X1 _26102_ ( .A1(_05311_ ), .A2(_05313_ ), .A3(_05314_ ), .ZN(_05315_ ) );
OR3_X1 _26103_ ( .A1(_04028_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04918_ ), .ZN(_05316_ ) );
INV_X1 _26104_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05317_ ) );
NAND4_X1 _26105_ ( .A1(_04109_ ), .A2(_04150_ ), .A3(_05317_ ), .A4(_04019_ ), .ZN(_05318_ ) );
AND3_X1 _26106_ ( .A1(_05315_ ), .A2(_05316_ ), .A3(_05318_ ), .ZN(_05319_ ) );
OR2_X1 _26107_ ( .A1(_04140_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05320_ ) );
INV_X1 _26108_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05321_ ) );
NAND4_X1 _26109_ ( .A1(_04147_ ), .A2(_04253_ ), .A3(_05321_ ), .A4(_04159_ ), .ZN(_05322_ ) );
NAND3_X1 _26110_ ( .A1(_05319_ ), .A2(_05320_ ), .A3(_05322_ ), .ZN(_05323_ ) );
MUX2_X1 _26111_ ( .A(_05289_ ), .B(_05323_ ), .S(_04428_ ), .Z(_05324_ ) );
BUF_X2 _26112_ ( .A(_05227_ ), .Z(_05325_ ) );
NOR3_X1 _26113_ ( .A1(_05325_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04320_ ), .ZN(_05326_ ) );
INV_X1 _26114_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05327_ ) );
AND4_X1 _26115_ ( .A1(_05327_ ), .A2(_04309_ ), .A3(_04171_ ), .A4(_04310_ ), .ZN(_05328_ ) );
OR3_X1 _26116_ ( .A1(_05324_ ), .A2(_05326_ ), .A3(_05328_ ), .ZN(_05329_ ) );
NOR4_X1 _26117_ ( .A1(_04544_ ), .A2(_04534_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04545_ ), .ZN(_05330_ ) );
NOR3_X1 _26118_ ( .A1(_04548_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04819_ ), .ZN(_05331_ ) );
NOR3_X1 _26119_ ( .A1(_05329_ ), .A2(_05330_ ), .A3(_05331_ ), .ZN(_05332_ ) );
INV_X1 _26120_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05333_ ) );
NAND4_X1 _26121_ ( .A1(_04197_ ), .A2(_04194_ ), .A3(_05333_ ), .A4(_04455_ ), .ZN(_05334_ ) );
OR3_X1 _26122_ ( .A1(_04326_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04819_ ), .ZN(_05335_ ) );
AND3_X1 _26123_ ( .A1(_05332_ ), .A2(_05334_ ), .A3(_05335_ ), .ZN(_05336_ ) );
INV_X1 _26124_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05337_ ) );
NAND4_X1 _26125_ ( .A1(_04620_ ), .A2(_04243_ ), .A3(_05337_ ), .A4(_04212_ ), .ZN(_05338_ ) );
OR3_X1 _26126_ ( .A1(_05202_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04637_ ), .ZN(_05339_ ) );
NAND3_X1 _26127_ ( .A1(_05336_ ), .A2(_05338_ ), .A3(_05339_ ), .ZN(_05340_ ) );
NOR3_X1 _26128_ ( .A1(_04636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04820_ ), .ZN(_05341_ ) );
AOI211_X1 _26129_ ( .A(_04015_ ), .B(_04023_ ), .C1(_04005_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05342_ ) );
NOR3_X1 _26130_ ( .A1(_05340_ ), .A2(_05341_ ), .A3(_05342_ ), .ZN(_05343_ ) );
INV_X1 _26131_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_05344_ ) );
OAI21_X1 _26132_ ( .A(_04246_ ), .B1(_05344_ ), .B2(_04251_ ), .ZN(_05345_ ) );
OAI22_X1 _26133_ ( .A1(_05288_ ), .A2(\idu.rs_reg ), .B1(_05343_ ), .B2(_05345_ ), .ZN(\idu.io_out_bits_rs1_data [11] ) );
NAND2_X1 _26134_ ( .A1(\exu.io_out_bits_rd_wdata [10] ), .A2(_04459_ ), .ZN(_05346_ ) );
OR3_X1 _26135_ ( .A1(_04667_ ), .A2(_10990_ ), .A3(\io_master_awaddr [1] ), .ZN(_05347_ ) );
NAND2_X1 _26136_ ( .A1(_04663_ ), .A2(_04664_ ), .ZN(_05348_ ) );
NAND3_X1 _26137_ ( .A1(_05348_ ), .A2(fanout_net_1 ), .A3(_04469_ ), .ZN(_05349_ ) );
NAND3_X1 _26138_ ( .A1(_03899_ ), .A2(_05347_ ), .A3(_05349_ ), .ZN(_05350_ ) );
OR4_X1 _26139_ ( .A1(_10989_ ), .A2(_04463_ ), .A3(lsu_io_out_bits_rd_wdata_$_MUX__Y_21_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A4(_04464_ ), .ZN(_05351_ ) );
OAI211_X1 _26140_ ( .A(fanout_net_1 ), .B(\io_master_rdata [10] ), .C1(_00968_ ), .C2(_00970_ ), .ZN(_05352_ ) );
AND2_X1 _26141_ ( .A1(_05351_ ), .A2(_05352_ ), .ZN(_05353_ ) );
AOI21_X1 _26142_ ( .A(_04903_ ), .B1(_04977_ ), .B2(_05353_ ), .ZN(_05354_ ) );
AOI221_X4 _26143_ ( .A(_03921_ ), .B1(_05350_ ), .B2(_05354_ ), .C1(_03915_ ), .C2(\lsu.io_in_bits_lb ), .ZN(_05355_ ) );
NOR2_X1 _26144_ ( .A1(\lsu.io_in_bits_ren ), .A2(\lsu.io_in_bits_rd_wdata [10] ), .ZN(_05356_ ) );
OAI21_X1 _26145_ ( .A(_04340_ ), .B1(_05355_ ), .B2(_05356_ ), .ZN(_05357_ ) );
AND4_X1 _26146_ ( .A1(\wbu.io_in_bits_rd_wdata [10] ), .A2(_03990_ ), .A3(_03997_ ), .A4(_04010_ ), .ZN(_05358_ ) );
OAI211_X1 _26147_ ( .A(_05357_ ), .B(_03856_ ), .C1(_04353_ ), .C2(_05358_ ), .ZN(_05359_ ) );
AOI21_X1 _26148_ ( .A(\idu.rs_reg ), .B1(_05346_ ), .B2(_05359_ ), .ZN(_05360_ ) );
NAND4_X1 _26149_ ( .A1(_04332_ ), .A2(_04241_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04842_ ), .ZN(_05361_ ) );
AND3_X1 _26150_ ( .A1(_04287_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04117_ ), .ZN(_05362_ ) );
INV_X1 _26151_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_05363_ ) );
NAND3_X1 _26152_ ( .A1(_04134_ ), .A2(_05363_ ), .A3(_11098_ ), .ZN(_05364_ ) );
MUX2_X1 _26153_ ( .A(_05364_ ), .B(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(_04053_ ), .Z(_05365_ ) );
INV_X1 _26154_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05366_ ) );
NAND4_X1 _26155_ ( .A1(_04098_ ), .A2(_04148_ ), .A3(_05366_ ), .A4(_11099_ ), .ZN(_05367_ ) );
OR2_X1 _26156_ ( .A1(_04069_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05368_ ) );
AND3_X1 _26157_ ( .A1(_05365_ ), .A2(_05367_ ), .A3(_05368_ ), .ZN(_05369_ ) );
INV_X1 _26158_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05370_ ) );
NAND4_X1 _26159_ ( .A1(_04107_ ), .A2(_04403_ ), .A3(_05370_ ), .A4(_04080_ ), .ZN(_05371_ ) );
INV_X1 _26160_ ( .A(_04077_ ), .ZN(_05372_ ) );
OR3_X1 _26161_ ( .A1(_05372_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03992_ ), .ZN(_05373_ ) );
NAND3_X1 _26162_ ( .A1(_05369_ ), .A2(_05371_ ), .A3(_05373_ ), .ZN(_05374_ ) );
INV_X1 _26163_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05375_ ) );
AND4_X1 _26164_ ( .A1(_05375_ ), .A2(_04144_ ), .A3(_04403_ ), .A4(_04040_ ), .ZN(_05376_ ) );
NOR3_X1 _26165_ ( .A1(_04186_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03993_ ), .ZN(_05377_ ) );
NOR3_X1 _26166_ ( .A1(_05374_ ), .A2(_05376_ ), .A3(_05377_ ), .ZN(_05378_ ) );
OR3_X1 _26167_ ( .A1(_05011_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03993_ ), .ZN(_05379_ ) );
OR3_X1 _26168_ ( .A1(_04095_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03993_ ), .ZN(_05380_ ) );
NAND3_X1 _26169_ ( .A1(_05378_ ), .A2(_05379_ ), .A3(_05380_ ), .ZN(_05381_ ) );
NOR2_X1 _26170_ ( .A1(_04102_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05382_ ) );
INV_X1 _26171_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05383_ ) );
AND4_X1 _26172_ ( .A1(_05383_ ), .A2(_04032_ ), .A3(_04037_ ), .A4(_04411_ ), .ZN(_05384_ ) );
NOR3_X1 _26173_ ( .A1(_05381_ ), .A2(_05382_ ), .A3(_05384_ ), .ZN(_05385_ ) );
INV_X1 _26174_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05386_ ) );
AOI22_X1 _26175_ ( .A1(_04285_ ), .A2(_05386_ ), .B1(_04118_ ), .B2(_04287_ ), .ZN(_05387_ ) );
AOI21_X1 _26176_ ( .A(_05362_ ), .B1(_05385_ ), .B2(_05387_ ), .ZN(_05388_ ) );
NOR3_X1 _26177_ ( .A1(_04943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04163_ ), .ZN(_05389_ ) );
INV_X1 _26178_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05390_ ) );
AND3_X1 _26179_ ( .A1(_04027_ ), .A2(_05390_ ), .A3(_04150_ ), .ZN(_05391_ ) );
NOR3_X1 _26180_ ( .A1(_05388_ ), .A2(_05389_ ), .A3(_05391_ ), .ZN(_05392_ ) );
INV_X1 _26181_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05393_ ) );
NAND4_X1 _26182_ ( .A1(_04936_ ), .A2(_04150_ ), .A3(_05393_ ), .A4(_04173_ ), .ZN(_05394_ ) );
OR2_X1 _26183_ ( .A1(_04140_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05395_ ) );
NAND3_X1 _26184_ ( .A1(_05392_ ), .A2(_05394_ ), .A3(_05395_ ), .ZN(_05396_ ) );
NOR4_X1 _26185_ ( .A1(_04126_ ), .A2(_04946_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04114_ ), .ZN(_05397_ ) );
NOR3_X1 _26186_ ( .A1(_04131_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04181_ ), .ZN(_05398_ ) );
NOR3_X1 _26187_ ( .A1(_05396_ ), .A2(_05397_ ), .A3(_05398_ ), .ZN(_05399_ ) );
OR3_X1 _26188_ ( .A1(_05325_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04295_ ), .ZN(_05400_ ) );
INV_X1 _26189_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05401_ ) );
NAND4_X1 _26190_ ( .A1(_04167_ ), .A2(_04297_ ), .A3(_05401_ ), .A4(_04174_ ), .ZN(_05402_ ) );
NAND3_X1 _26191_ ( .A1(_05399_ ), .A2(_05400_ ), .A3(_05402_ ), .ZN(_05403_ ) );
INV_X1 _26192_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05404_ ) );
AND4_X1 _26193_ ( .A1(_05404_ ), .A2(_04147_ ), .A3(_04156_ ), .A4(_04174_ ), .ZN(_05405_ ) );
NOR3_X1 _26194_ ( .A1(_04187_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04190_ ), .ZN(_05406_ ) );
NOR3_X1 _26195_ ( .A1(_05403_ ), .A2(_05405_ ), .A3(_05406_ ), .ZN(_05407_ ) );
INV_X1 _26196_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05408_ ) );
NAND4_X1 _26197_ ( .A1(_04196_ ), .A2(_04000_ ), .A3(_05408_ ), .A4(_10756_ ), .ZN(_05409_ ) );
INV_X1 _26198_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05410_ ) );
NAND4_X1 _26199_ ( .A1(_04332_ ), .A2(_04171_ ), .A3(_05410_ ), .A4(_04209_ ), .ZN(_05411_ ) );
NAND3_X1 _26200_ ( .A1(_05407_ ), .A2(_05409_ ), .A3(_05411_ ), .ZN(_05412_ ) );
OAI21_X1 _26201_ ( .A(_05361_ ), .B1(_05412_ ), .B2(_04201_ ), .ZN(_05413_ ) );
OR3_X1 _26202_ ( .A1(_05201_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04549_ ), .ZN(_05414_ ) );
INV_X1 _26203_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05415_ ) );
NAND3_X1 _26204_ ( .A1(_04215_ ), .A2(_05415_ ), .A3(_04223_ ), .ZN(_05416_ ) );
AND3_X1 _26205_ ( .A1(_05413_ ), .A2(_05414_ ), .A3(_05416_ ), .ZN(_05417_ ) );
INV_X1 _26206_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05418_ ) );
OAI211_X1 _26207_ ( .A(_04221_ ), .B(_10792_ ), .C1(_05418_ ), .C2(_04455_ ), .ZN(_05419_ ) );
AOI221_X4 _26208_ ( .A(_04240_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B2(_04250_ ), .C1(_05417_ ), .C2(_05419_ ), .ZN(_05420_ ) );
OR2_X1 _26209_ ( .A1(_05360_ ), .A2(_05420_ ), .ZN(\idu.io_out_bits_rs1_data [10] ) );
NOR2_X1 _26210_ ( .A1(_05355_ ), .A2(_05356_ ), .ZN(\lsu.io_out_bits_rd_wdata [10] ) );
NAND2_X1 _26211_ ( .A1(\exu.io_out_bits_rd_wdata [9] ), .A2(_04356_ ), .ZN(_05421_ ) );
NAND3_X1 _26212_ ( .A1(_04752_ ), .A2(_03872_ ), .A3(_04753_ ), .ZN(_05422_ ) );
OR3_X1 _26213_ ( .A1(_04756_ ), .A2(\io_master_awaddr [0] ), .A3(_04757_ ), .ZN(_05423_ ) );
NAND3_X1 _26214_ ( .A1(_03899_ ), .A2(_05422_ ), .A3(_05423_ ), .ZN(_05424_ ) );
OR4_X1 _26215_ ( .A1(_10989_ ), .A2(_00968_ ), .A3(lsu_io_out_bits_rd_wdata_$_MUX__Y_22_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A4(_00970_ ), .ZN(_05425_ ) );
OAI211_X1 _26216_ ( .A(fanout_net_1 ), .B(\io_master_rdata [9] ), .C1(_00968_ ), .C2(_00970_ ), .ZN(_05426_ ) );
AND2_X1 _26217_ ( .A1(_05425_ ), .A2(_05426_ ), .ZN(_05427_ ) );
OAI21_X1 _26218_ ( .A(_05427_ ), .B1(_04462_ ), .B2(_03883_ ), .ZN(_05428_ ) );
NAND3_X1 _26219_ ( .A1(_05424_ ), .A2(_04904_ ), .A3(_05428_ ), .ZN(_05429_ ) );
OAI211_X1 _26220_ ( .A(\lsu.io_in_bits_ren ), .B(_05429_ ), .C1(_05283_ ), .C2(_05284_ ), .ZN(_05430_ ) );
OR2_X1 _26221_ ( .A1(\lsu.io_in_bits_ren ), .A2(\lsu.io_in_bits_rd_wdata [9] ), .ZN(_05431_ ) );
NAND3_X1 _26222_ ( .A1(_05430_ ), .A2(_04340_ ), .A3(_05431_ ), .ZN(_05432_ ) );
OAI211_X1 _26223_ ( .A(\wbu.io_in_bits_rd_wdata [9] ), .B(_04656_ ), .C1(_04657_ ), .C2(_04658_ ), .ZN(_05433_ ) );
NAND2_X1 _26224_ ( .A1(_05432_ ), .A2(_05433_ ), .ZN(_05434_ ) );
NAND2_X1 _26225_ ( .A1(_05434_ ), .A2(_04738_ ), .ZN(_05435_ ) );
AOI21_X1 _26226_ ( .A(\idu.rs_reg ), .B1(_05421_ ), .B2(_05435_ ), .ZN(_05436_ ) );
INV_X1 _26227_ ( .A(_04045_ ), .ZN(_05437_ ) );
OR4_X1 _26228_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_05437_ ), .A3(_04124_ ), .A4(_04017_ ), .ZN(_05438_ ) );
NAND4_X1 _26229_ ( .A1(_04107_ ), .A2(_04154_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_11100_ ), .ZN(_05439_ ) );
OR4_X1 _26230_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A2(_04051_ ), .A3(_10766_ ), .A4(_04263_ ), .ZN(_05440_ ) );
OAI21_X1 _26231_ ( .A(_05440_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05293_ ), .ZN(_05441_ ) );
INV_X1 _26232_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05442_ ) );
AOI21_X1 _26233_ ( .A(_05441_ ), .B1(_05442_ ), .B2(_04392_ ), .ZN(_05443_ ) );
OR2_X1 _26234_ ( .A1(_04070_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05444_ ) );
NAND2_X1 _26235_ ( .A1(_05443_ ), .A2(_05444_ ), .ZN(_05445_ ) );
OAI21_X1 _26236_ ( .A(_05439_ ), .B1(_05445_ ), .B2(_04395_ ), .ZN(_05446_ ) );
INV_X1 _26237_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05447_ ) );
NAND3_X1 _26238_ ( .A1(_04078_ ), .A2(_05447_ ), .A3(_04411_ ), .ZN(_05448_ ) );
OR4_X1 _26239_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04123_ ), .A3(_04180_ ), .A4(_04016_ ), .ZN(_05449_ ) );
NAND3_X1 _26240_ ( .A1(_05446_ ), .A2(_05448_ ), .A3(_05449_ ), .ZN(_05450_ ) );
NOR3_X1 _26241_ ( .A1(_04186_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04017_ ), .ZN(_05451_ ) );
INV_X1 _26242_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05452_ ) );
AND3_X1 _26243_ ( .A1(_04257_ ), .A2(_05452_ ), .A3(_04107_ ), .ZN(_05453_ ) );
NOR4_X1 _26244_ ( .A1(_05450_ ), .A2(_04845_ ), .A3(_05451_ ), .A4(_05453_ ), .ZN(_05454_ ) );
AND4_X1 _26245_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04331_ ), .A3(_04117_ ), .A4(_11101_ ), .ZN(_05455_ ) );
OAI21_X1 _26246_ ( .A(_05438_ ), .B1(_05454_ ), .B2(_05455_ ), .ZN(_05456_ ) );
INV_X1 _26247_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05457_ ) );
AND4_X1 _26248_ ( .A1(_05457_ ), .A2(_04110_ ), .A3(_04038_ ), .A4(_04598_ ), .ZN(_05458_ ) );
NOR3_X1 _26249_ ( .A1(_04519_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04018_ ), .ZN(_05459_ ) );
NOR3_X1 _26250_ ( .A1(_05456_ ), .A2(_05458_ ), .A3(_05459_ ), .ZN(_05460_ ) );
OR2_X1 _26251_ ( .A1(_05019_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05461_ ) );
OR3_X1 _26252_ ( .A1(_04943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04163_ ), .ZN(_05462_ ) );
NAND3_X1 _26253_ ( .A1(_05460_ ), .A2(_05461_ ), .A3(_05462_ ), .ZN(_05463_ ) );
NOR3_X1 _26254_ ( .A1(_04131_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04946_ ), .ZN(_05464_ ) );
NOR3_X1 _26255_ ( .A1(_04294_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04189_ ), .ZN(_05465_ ) );
NOR3_X1 _26256_ ( .A1(_05463_ ), .A2(_05464_ ), .A3(_05465_ ), .ZN(_05466_ ) );
INV_X1 _26257_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05467_ ) );
NAND4_X1 _26258_ ( .A1(_04170_ ), .A2(_04151_ ), .A3(_05467_ ), .A4(_04020_ ), .ZN(_05468_ ) );
INV_X1 _26259_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05469_ ) );
NAND4_X1 _26260_ ( .A1(_04241_ ), .A2(_04151_ ), .A3(_05469_ ), .A4(_04020_ ), .ZN(_05470_ ) );
NAND3_X1 _26261_ ( .A1(_05466_ ), .A2(_05468_ ), .A3(_05470_ ), .ZN(_05471_ ) );
NOR3_X1 _26262_ ( .A1(_04029_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04317_ ), .ZN(_05472_ ) );
INV_X1 _26263_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05473_ ) );
AND4_X1 _26264_ ( .A1(_05473_ ), .A2(_04216_ ), .A3(_04156_ ), .A4(_04159_ ), .ZN(_05474_ ) );
NOR3_X1 _26265_ ( .A1(_05471_ ), .A2(_05472_ ), .A3(_05474_ ), .ZN(_05475_ ) );
INV_X1 _26266_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05476_ ) );
NAND4_X1 _26267_ ( .A1(_04168_ ), .A2(_04171_ ), .A3(_05476_ ), .A4(_04313_ ), .ZN(_05477_ ) );
OR4_X1 _26268_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04178_ ), .A3(_04181_ ), .A4(_04437_ ), .ZN(_05478_ ) );
NAND3_X1 _26269_ ( .A1(_05475_ ), .A2(_05477_ ), .A3(_05478_ ), .ZN(_05479_ ) );
NOR3_X1 _26270_ ( .A1(_04188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04320_ ), .ZN(_05480_ ) );
NOR3_X1 _26271_ ( .A1(_05011_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04320_ ), .ZN(_05481_ ) );
NOR3_X1 _26272_ ( .A1(_05479_ ), .A2(_05480_ ), .A3(_05481_ ), .ZN(_05482_ ) );
OR3_X1 _26273_ ( .A1(_04326_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04191_ ), .ZN(_05483_ ) );
INV_X1 _26274_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05484_ ) );
NAND4_X1 _26275_ ( .A1(_04333_ ), .A2(_04242_ ), .A3(_05484_ ), .A4(_04538_ ), .ZN(_05485_ ) );
NAND3_X1 _26276_ ( .A1(_05482_ ), .A2(_05483_ ), .A3(_05485_ ), .ZN(_05486_ ) );
NOR3_X1 _26277_ ( .A1(_05202_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04819_ ), .ZN(_05487_ ) );
INV_X1 _26278_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05488_ ) );
AND3_X1 _26279_ ( .A1(_04215_ ), .A2(_05488_ ), .A3(_04223_ ), .ZN(_05489_ ) );
NOR3_X1 _26280_ ( .A1(_05486_ ), .A2(_05487_ ), .A3(_05489_ ), .ZN(_05490_ ) );
INV_X1 _26281_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05491_ ) );
OAI211_X1 _26282_ ( .A(_04215_ ), .B(_10792_ ), .C1(_05491_ ), .C2(_04455_ ), .ZN(_05492_ ) );
AOI221_X4 _26283_ ( .A(_04240_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B2(_04250_ ), .C1(_05490_ ), .C2(_05492_ ), .ZN(_05493_ ) );
OR2_X1 _26284_ ( .A1(_05436_ ), .A2(_05493_ ), .ZN(\idu.io_out_bits_rs1_data [9] ) );
AND2_X1 _26285_ ( .A1(_05430_ ), .A2(_05431_ ), .ZN(\lsu.io_out_bits_rd_wdata [9] ) );
AOI21_X1 _26286_ ( .A(_03857_ ), .B1(_02916_ ), .B2(_02917_ ), .ZN(_05494_ ) );
OAI211_X1 _26287_ ( .A(fanout_net_1 ), .B(\io_master_rdata [8] ), .C1(_00968_ ), .C2(_00970_ ), .ZN(_05495_ ) );
OR4_X1 _26288_ ( .A1(_10989_ ), .A2(_00968_ ), .A3(lsu_io_out_bits_rd_wdata_$_MUX__Y_23_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ), .A4(_00970_ ), .ZN(_05496_ ) );
AND3_X1 _26289_ ( .A1(_04977_ ), .A2(_05495_ ), .A3(_05496_ ), .ZN(_05497_ ) );
BUF_X2 _26290_ ( .A(_04977_ ), .Z(_05498_ ) );
AOI21_X1 _26291_ ( .A(\io_master_awaddr [0] ), .B1(_04827_ ), .B2(_04828_ ), .ZN(_05499_ ) );
AND3_X1 _26292_ ( .A1(_04830_ ), .A2(_03872_ ), .A3(_04831_ ), .ZN(_05500_ ) );
NOR3_X1 _26293_ ( .A1(_05498_ ), .A2(_05499_ ), .A3(_05500_ ), .ZN(_05501_ ) );
NOR3_X1 _26294_ ( .A1(_05497_ ), .A2(_05501_ ), .A3(_04903_ ), .ZN(_05502_ ) );
AOI211_X1 _26295_ ( .A(_03926_ ), .B(_05502_ ), .C1(_03915_ ), .C2(\lsu.io_in_bits_lb ), .ZN(_05503_ ) );
NOR2_X1 _26296_ ( .A1(\lsu.io_in_bits_ren ), .A2(\lsu.io_in_bits_rd_wdata [8] ), .ZN(_05504_ ) );
NOR2_X1 _26297_ ( .A1(_05503_ ), .A2(_05504_ ), .ZN(\lsu.io_out_bits_rd_wdata [8] ) );
NOR2_X1 _26298_ ( .A1(\lsu.io_out_bits_rd_wdata [8] ), .A2(_03931_ ), .ZN(_05505_ ) );
NAND4_X1 _26299_ ( .A1(_03991_ ), .A2(\wbu.io_in_bits_rd_wdata [8] ), .A3(_03998_ ), .A4(_04011_ ), .ZN(_05506_ ) );
AOI211_X1 _26300_ ( .A(_04459_ ), .B(_05505_ ), .C1(_03932_ ), .C2(_05506_ ), .ZN(_05507_ ) );
OAI21_X1 _26301_ ( .A(_03851_ ), .B1(_05494_ ), .B2(_05507_ ), .ZN(_05508_ ) );
NAND3_X1 _26302_ ( .A1(_04571_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04482_ ), .ZN(_05509_ ) );
OR3_X1 _26303_ ( .A1(_04943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04173_ ), .ZN(_05510_ ) );
NOR3_X1 _26304_ ( .A1(_04592_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03994_ ), .ZN(_05511_ ) );
OR3_X1 _26305_ ( .A1(_04263_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10767_ ), .ZN(_05512_ ) );
OAI21_X1 _26306_ ( .A(_05512_ ), .B1(_05293_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05513_ ) );
NOR4_X1 _26307_ ( .A1(_04123_ ), .A2(_04918_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_10767_ ), .ZN(_05514_ ) );
NOR2_X1 _26308_ ( .A1(_05513_ ), .A2(_05514_ ), .ZN(_05515_ ) );
OAI21_X1 _26309_ ( .A(_05515_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04497_ ), .ZN(_05516_ ) );
AOI211_X1 _26310_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_05325_ ), .C1(\idu.io_in_bits_inst [19] ), .C2(_11030_ ), .ZN(_05517_ ) );
OAI21_X1 _26311_ ( .A(_04085_ ), .B1(_04272_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05518_ ) );
OR3_X1 _26312_ ( .A1(_05516_ ), .A2(_05517_ ), .A3(_05518_ ), .ZN(_05519_ ) );
NAND3_X1 _26313_ ( .A1(_04082_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04042_ ), .ZN(_05520_ ) );
AOI21_X1 _26314_ ( .A(_05511_ ), .B1(_05519_ ), .B2(_05520_ ), .ZN(_05521_ ) );
INV_X1 _26315_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05522_ ) );
NAND3_X1 _26316_ ( .A1(_04504_ ), .A2(_05522_ ), .A3(_04385_ ), .ZN(_05523_ ) );
INV_X1 _26317_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05524_ ) );
NAND4_X1 _26318_ ( .A1(_04331_ ), .A2(_04118_ ), .A3(_05524_ ), .A4(_04598_ ), .ZN(_05525_ ) );
AND3_X1 _26319_ ( .A1(_05521_ ), .A2(_05523_ ), .A3(_05525_ ), .ZN(_05526_ ) );
OR4_X1 _26320_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_05437_ ), .A3(_04125_ ), .A4(_04128_ ), .ZN(_05527_ ) );
OR3_X1 _26321_ ( .A1(_05201_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04018_ ), .ZN(_05528_ ) );
NAND4_X1 _26322_ ( .A1(_05526_ ), .A2(_04704_ ), .A3(_05527_ ), .A4(_05528_ ), .ZN(_05529_ ) );
NAND4_X1 _26323_ ( .A1(_04936_ ), .A2(_04522_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04295_ ), .ZN(_05530_ ) );
AOI21_X1 _26324_ ( .A(_04516_ ), .B1(_05529_ ), .B2(_05530_ ), .ZN(_05531_ ) );
AND3_X1 _26325_ ( .A1(_04606_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04170_ ), .ZN(_05532_ ) );
OAI21_X1 _26326_ ( .A(_05510_ ), .B1(_05531_ ), .B2(_05532_ ), .ZN(_05533_ ) );
NOR3_X1 _26327_ ( .A1(_04029_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04947_ ), .ZN(_05534_ ) );
NOR3_X1 _26328_ ( .A1(_04485_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04190_ ), .ZN(_05535_ ) );
OR3_X1 _26329_ ( .A1(_05533_ ), .A2(_05534_ ), .A3(_05535_ ), .ZN(_05536_ ) );
INV_X1 _26330_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05537_ ) );
AND4_X1 _26331_ ( .A1(_05537_ ), .A2(_04171_ ), .A3(_04529_ ), .A4(_04313_ ), .ZN(_05538_ ) );
NOR4_X1 _26332_ ( .A1(_04179_ ), .A2(_04947_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04318_ ), .ZN(_05539_ ) );
NOR3_X1 _26333_ ( .A1(_05536_ ), .A2(_05538_ ), .A3(_05539_ ), .ZN(_05540_ ) );
INV_X1 _26334_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05541_ ) );
NAND4_X1 _26335_ ( .A1(_04536_ ), .A2(_04451_ ), .A3(_05541_ ), .A4(_04538_ ), .ZN(_05542_ ) );
OR3_X1 _26336_ ( .A1(_05325_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04549_ ), .ZN(_05543_ ) );
NAND3_X1 _26337_ ( .A1(_05540_ ), .A2(_05542_ ), .A3(_05543_ ), .ZN(_05544_ ) );
INV_X1 _26338_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05545_ ) );
AND4_X1 _26339_ ( .A1(_05545_ ), .A2(_04542_ ), .A3(_04528_ ), .A4(_04623_ ), .ZN(_05546_ ) );
NOR4_X1 _26340_ ( .A1(_04179_ ), .A2(_04534_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04545_ ), .ZN(_05547_ ) );
NOR3_X1 _26341_ ( .A1(_05544_ ), .A2(_05546_ ), .A3(_05547_ ), .ZN(_05548_ ) );
OR3_X1 _26342_ ( .A1(_04548_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04819_ ), .ZN(_05549_ ) );
OR3_X1 _26343_ ( .A1(_05011_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04819_ ), .ZN(_05550_ ) );
NAND3_X1 _26344_ ( .A1(_05548_ ), .A2(_05549_ ), .A3(_05550_ ), .ZN(_05551_ ) );
INV_X1 _26345_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05552_ ) );
AND4_X1 _26346_ ( .A1(_05552_ ), .A2(_04333_ ), .A3(_04728_ ), .A4(_04624_ ), .ZN(_05553_ ) );
BUF_X2 _26347_ ( .A(_05437_ ), .Z(_05554_ ) );
NOR4_X1 _26348_ ( .A1(_05554_ ), .A2(_04544_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04550_ ), .ZN(_05555_ ) );
NOR3_X1 _26349_ ( .A1(_05551_ ), .A2(_05553_ ), .A3(_05555_ ), .ZN(_05556_ ) );
OR3_X1 _26350_ ( .A1(_05202_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04820_ ), .ZN(_05557_ ) );
INV_X1 _26351_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05558_ ) );
NAND3_X1 _26352_ ( .A1(_04562_ ), .A2(_05558_ ), .A3(_04224_ ), .ZN(_05559_ ) );
NAND3_X1 _26353_ ( .A1(_05556_ ), .A2(_05557_ ), .A3(_05559_ ), .ZN(_05560_ ) );
AOI211_X1 _26354_ ( .A(_04566_ ), .B(_04567_ ), .C1(_04568_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05561_ ) );
OAI211_X1 _26355_ ( .A(_04481_ ), .B(_05509_ ), .C1(_05560_ ), .C2(_05561_ ), .ZN(_05562_ ) );
NAND2_X1 _26356_ ( .A1(_05508_ ), .A2(_05562_ ), .ZN(\idu.io_out_bits_rs1_data [8] ) );
NAND2_X1 _26357_ ( .A1(\exu.io_out_bits_rd_wdata [7] ), .A2(_04356_ ), .ZN(_05563_ ) );
OR3_X1 _26358_ ( .A1(_04904_ ), .A2(\lsu.io_in_bits_lbu ), .A3(\lsu.io_in_bits_lb ), .ZN(_05564_ ) );
AND2_X2 _26359_ ( .A1(_05564_ ), .A2(\lsu.io_in_bits_ren ), .ZN(_05565_ ) );
AND2_X1 _26360_ ( .A1(_03915_ ), .A2(_05565_ ), .ZN(_05566_ ) );
AND2_X1 _26361_ ( .A1(_03926_ ), .A2(\lsu.io_in_bits_rd_wdata [7] ), .ZN(_05567_ ) );
OAI21_X1 _26362_ ( .A(_04340_ ), .B1(_05566_ ), .B2(_05567_ ), .ZN(_05568_ ) );
OR3_X1 _26363_ ( .A1(_03989_ ), .A2(_13919_ ), .A3(_04236_ ), .ZN(_05569_ ) );
OAI21_X1 _26364_ ( .A(_05568_ ), .B1(_04340_ ), .B2(_05569_ ), .ZN(_05570_ ) );
NAND2_X1 _26365_ ( .A1(_05570_ ), .A2(_03856_ ), .ZN(_05571_ ) );
AOI21_X1 _26366_ ( .A(\idu.rs_reg ), .B1(_05563_ ), .B2(_05571_ ), .ZN(_05572_ ) );
INV_X1 _26367_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05573_ ) );
AND4_X1 _26368_ ( .A1(_05573_ ), .A2(_04385_ ), .A3(_04110_ ), .A4(_04598_ ), .ZN(_05574_ ) );
NOR2_X1 _26369_ ( .A1(_04054_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05575_ ) );
NOR3_X1 _26370_ ( .A1(_04263_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10767_ ), .ZN(_05576_ ) );
NOR4_X1 _26371_ ( .A1(_04123_ ), .A2(_04918_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_10766_ ), .ZN(_05577_ ) );
NOR3_X1 _26372_ ( .A1(_05575_ ), .A2(_05576_ ), .A3(_05577_ ), .ZN(_05578_ ) );
OR2_X1 _26373_ ( .A1(_04069_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05579_ ) );
INV_X1 _26374_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05580_ ) );
NAND4_X1 _26375_ ( .A1(_04073_ ), .A2(_04074_ ), .A3(_05580_ ), .A4(_04039_ ), .ZN(_05581_ ) );
AND3_X1 _26376_ ( .A1(_05578_ ), .A2(_05579_ ), .A3(_05581_ ), .ZN(_05582_ ) );
OR3_X1 _26377_ ( .A1(_05372_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03992_ ), .ZN(_05583_ ) );
OR4_X1 _26378_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04123_ ), .A3(_04180_ ), .A4(_10767_ ), .ZN(_05584_ ) );
NAND3_X1 _26379_ ( .A1(_05582_ ), .A2(_05583_ ), .A3(_05584_ ), .ZN(_05585_ ) );
NOR3_X1 _26380_ ( .A1(_04186_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03993_ ), .ZN(_05586_ ) );
INV_X1 _26381_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05587_ ) );
AND3_X1 _26382_ ( .A1(_04088_ ), .A2(_05587_ ), .A3(_04073_ ), .ZN(_05588_ ) );
OR3_X1 _26383_ ( .A1(_05585_ ), .A2(_05586_ ), .A3(_05588_ ), .ZN(_05589_ ) );
NOR3_X1 _26384_ ( .A1(_04095_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03994_ ), .ZN(_05590_ ) );
OAI21_X1 _26385_ ( .A(_04413_ ), .B1(_04101_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05591_ ) );
OR3_X1 _26386_ ( .A1(_05589_ ), .A2(_05590_ ), .A3(_05591_ ), .ZN(_05592_ ) );
NAND3_X1 _26387_ ( .A1(_04287_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04038_ ), .ZN(_05593_ ) );
AOI21_X1 _26388_ ( .A(_05574_ ), .B1(_05592_ ), .B2(_05593_ ), .ZN(_05594_ ) );
OR2_X1 _26389_ ( .A1(_05019_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05595_ ) );
INV_X1 _26390_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05596_ ) );
NAND4_X1 _26391_ ( .A1(_04146_ ), .A2(_04111_ ), .A3(_05596_ ), .A4(_04513_ ), .ZN(_05597_ ) );
NAND3_X1 _26392_ ( .A1(_05594_ ), .A2(_05595_ ), .A3(_05597_ ), .ZN(_05598_ ) );
NOR3_X1 _26393_ ( .A1(_04131_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04946_ ), .ZN(_05599_ ) );
NOR3_X1 _26394_ ( .A1(_04294_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04189_ ), .ZN(_05600_ ) );
NOR3_X1 _26395_ ( .A1(_05598_ ), .A2(_05599_ ), .A3(_05600_ ), .ZN(_05601_ ) );
INV_X1 _26396_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05602_ ) );
NAND4_X1 _26397_ ( .A1(_04170_ ), .A2(_04151_ ), .A3(_05602_ ), .A4(_04020_ ), .ZN(_05603_ ) );
OR4_X1 _26398_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04125_ ), .A3(_04946_ ), .A4(_04513_ ), .ZN(_05604_ ) );
NAND3_X1 _26399_ ( .A1(_05601_ ), .A2(_05603_ ), .A3(_05604_ ), .ZN(_05605_ ) );
NOR3_X1 _26400_ ( .A1(_04029_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04317_ ), .ZN(_05606_ ) );
INV_X1 _26401_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05607_ ) );
AND4_X1 _26402_ ( .A1(_05607_ ), .A2(_04936_ ), .A3(_04156_ ), .A4(_04159_ ), .ZN(_05608_ ) );
NOR3_X1 _26403_ ( .A1(_05605_ ), .A2(_05606_ ), .A3(_05608_ ), .ZN(_05609_ ) );
INV_X1 _26404_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05610_ ) );
NAND4_X1 _26405_ ( .A1(_04168_ ), .A2(_04171_ ), .A3(_05610_ ), .A4(_04313_ ), .ZN(_05611_ ) );
OR4_X1 _26406_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04178_ ), .A3(_04181_ ), .A4(_04437_ ), .ZN(_05612_ ) );
NAND3_X1 _26407_ ( .A1(_05609_ ), .A2(_05611_ ), .A3(_05612_ ), .ZN(_05613_ ) );
NOR3_X1 _26408_ ( .A1(_04187_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04320_ ), .ZN(_05614_ ) );
INV_X1 _26409_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05615_ ) );
AND4_X1 _26410_ ( .A1(_04000_ ), .A2(_04196_ ), .A3(_05615_ ), .A4(_10756_ ), .ZN(_05616_ ) );
NOR3_X1 _26411_ ( .A1(_05613_ ), .A2(_05614_ ), .A3(_05616_ ), .ZN(_05617_ ) );
INV_X1 _26412_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05618_ ) );
NAND4_X1 _26413_ ( .A1(_04333_ ), .A2(_04615_ ), .A3(_05618_ ), .A4(_04538_ ), .ZN(_05619_ ) );
OR4_X1 _26414_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_05554_ ), .A3(_04316_ ), .A4(_04318_ ), .ZN(_05620_ ) );
NAND3_X1 _26415_ ( .A1(_05617_ ), .A2(_05619_ ), .A3(_05620_ ), .ZN(_05621_ ) );
INV_X1 _26416_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05622_ ) );
AND4_X1 _26417_ ( .A1(_05622_ ), .A2(_04445_ ), .A3(_04451_ ), .A4(_04623_ ), .ZN(_05623_ ) );
INV_X1 _26418_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05624_ ) );
AND3_X1 _26419_ ( .A1(_04215_ ), .A2(_05624_ ), .A3(_04223_ ), .ZN(_05625_ ) );
NOR3_X1 _26420_ ( .A1(_05621_ ), .A2(_05623_ ), .A3(_05625_ ), .ZN(_05626_ ) );
INV_X1 _26421_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05627_ ) );
OAI211_X1 _26422_ ( .A(_04215_ ), .B(_10792_ ), .C1(_05627_ ), .C2(_04455_ ), .ZN(_05628_ ) );
AOI221_X4 _26423_ ( .A(_04240_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B2(_04250_ ), .C1(_05626_ ), .C2(_05628_ ), .ZN(_05629_ ) );
OR2_X1 _26424_ ( .A1(_05572_ ), .A2(_05629_ ), .ZN(\idu.io_out_bits_rs1_data [7] ) );
NOR2_X1 _26425_ ( .A1(_05566_ ), .A2(_05567_ ), .ZN(_05630_ ) );
INV_X1 _26426_ ( .A(_05630_ ), .ZN(\lsu.io_out_bits_rd_wdata [7] ) );
OAI21_X1 _26427_ ( .A(fanout_net_1 ), .B1(_08562_ ), .B2(\io_master_rdata [6] ), .ZN(_05631_ ) );
AND4_X1 _26428_ ( .A1(fanout_net_1 ), .A2(_04982_ ), .A3(_04983_ ), .A4(lsu_io_out_bits_rd_wdata_$_MUX__Y_9_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05632_ ) );
OAI21_X1 _26429_ ( .A(_05498_ ), .B1(_05631_ ), .B2(_05632_ ), .ZN(_05633_ ) );
NAND2_X1 _26430_ ( .A1(_04981_ ), .A2(_04984_ ), .ZN(_05634_ ) );
MUX2_X1 _26431_ ( .A(_05634_ ), .B(_04347_ ), .S(\io_master_awaddr [0] ), .Z(_05635_ ) );
AOI22_X1 _26432_ ( .A1(_05635_ ), .A2(\io_master_awaddr [1] ), .B1(_03906_ ), .B2(_04980_ ), .ZN(_05636_ ) );
OAI211_X1 _26433_ ( .A(_05565_ ), .B(_05633_ ), .C1(_05636_ ), .C2(_04462_ ), .ZN(_05637_ ) );
NAND2_X1 _26434_ ( .A1(_03927_ ), .A2(\lsu.io_in_bits_rd_wdata [6] ), .ZN(_05638_ ) );
AND3_X1 _26435_ ( .A1(_05637_ ), .A2(_03925_ ), .A3(_05638_ ), .ZN(_05639_ ) );
NAND4_X1 _26436_ ( .A1(_03990_ ), .A2(\wbu.io_in_bits_rd_wdata [6] ), .A3(_03997_ ), .A4(_04010_ ), .ZN(_05640_ ) );
AOI211_X1 _26437_ ( .A(_03859_ ), .B(_05639_ ), .C1(_03931_ ), .C2(_05640_ ), .ZN(_05641_ ) );
AOI21_X1 _26438_ ( .A(_05641_ ), .B1(\exu.io_out_bits_rd_wdata [6] ), .B2(_04459_ ), .ZN(_05642_ ) );
OR4_X1 _26439_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_05437_ ), .A3(_04124_ ), .A4(_03994_ ), .ZN(_05643_ ) );
INV_X1 _26440_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_05644_ ) );
NAND3_X1 _26441_ ( .A1(_04134_ ), .A2(_05644_ ), .A3(_11099_ ), .ZN(_05645_ ) );
MUX2_X1 _26442_ ( .A(_05645_ ), .B(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(_04053_ ), .Z(_05646_ ) );
INV_X1 _26443_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05647_ ) );
NAND4_X1 _26444_ ( .A1(_04144_ ), .A2(_04149_ ), .A3(_05647_ ), .A4(_11100_ ), .ZN(_05648_ ) );
OR2_X1 _26445_ ( .A1(_04497_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05649_ ) );
NAND3_X1 _26446_ ( .A1(_05646_ ), .A2(_05648_ ), .A3(_05649_ ), .ZN(_05650_ ) );
INV_X1 _26447_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05651_ ) );
AND4_X1 _26448_ ( .A1(_05651_ ), .A2(_04107_ ), .A3(_04154_ ), .A4(_04080_ ), .ZN(_05652_ ) );
CLKBUF_X2 _26449_ ( .A(_05372_ ), .Z(_05653_ ) );
NOR3_X1 _26450_ ( .A1(_05653_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04127_ ), .ZN(_05654_ ) );
NOR3_X1 _26451_ ( .A1(_05650_ ), .A2(_05652_ ), .A3(_05654_ ), .ZN(_05655_ ) );
INV_X1 _26452_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05656_ ) );
NAND4_X1 _26453_ ( .A1(_04145_ ), .A2(_04858_ ), .A3(_05656_ ), .A4(_11101_ ), .ZN(_05657_ ) );
NAND2_X1 _26454_ ( .A1(_05655_ ), .A2(_05657_ ), .ZN(_05658_ ) );
NOR3_X1 _26455_ ( .A1(_04592_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04128_ ), .ZN(_05659_ ) );
OAI22_X1 _26456_ ( .A1(_04093_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(_04095_ ), .B2(_04138_ ), .ZN(_05660_ ) );
NOR3_X1 _26457_ ( .A1(_05658_ ), .A2(_05659_ ), .A3(_05660_ ), .ZN(_05661_ ) );
AND3_X1 _26458_ ( .A1(_04048_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04283_ ), .ZN(_05662_ ) );
OAI21_X1 _26459_ ( .A(_05643_ ), .B1(_05661_ ), .B2(_05662_ ), .ZN(_05663_ ) );
NOR3_X1 _26460_ ( .A1(_05201_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04129_ ), .ZN(_05664_ ) );
INV_X1 _26461_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05665_ ) );
AND4_X1 _26462_ ( .A1(_05665_ ), .A2(_04385_ ), .A3(_04110_ ), .A4(_04113_ ), .ZN(_05666_ ) );
NOR3_X1 _26463_ ( .A1(_05663_ ), .A2(_05664_ ), .A3(_05666_ ), .ZN(_05667_ ) );
OR2_X1 _26464_ ( .A1(_05019_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05668_ ) );
INV_X1 _26465_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05669_ ) );
NAND4_X1 _26466_ ( .A1(_04147_ ), .A2(_04522_ ), .A3(_05669_ ), .A4(_04295_ ), .ZN(_05670_ ) );
AND3_X1 _26467_ ( .A1(_05667_ ), .A2(_05668_ ), .A3(_05670_ ), .ZN(_05671_ ) );
OR3_X1 _26468_ ( .A1(_04131_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04946_ ), .ZN(_05672_ ) );
OR3_X1 _26469_ ( .A1(_04294_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04295_ ), .ZN(_05673_ ) );
NAND3_X1 _26470_ ( .A1(_05671_ ), .A2(_05672_ ), .A3(_05673_ ), .ZN(_05674_ ) );
INV_X1 _26471_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05675_ ) );
AND4_X1 _26472_ ( .A1(_05675_ ), .A2(_04297_ ), .A3(_04151_ ), .A4(_04174_ ), .ZN(_05676_ ) );
OAI21_X1 _26473_ ( .A(_04428_ ), .B1(_04303_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05677_ ) );
NOR3_X1 _26474_ ( .A1(_05674_ ), .A2(_05676_ ), .A3(_05677_ ), .ZN(_05678_ ) );
AND3_X1 _26475_ ( .A1(_04444_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04309_ ), .ZN(_05679_ ) );
NOR2_X1 _26476_ ( .A1(_05678_ ), .A2(_05679_ ), .ZN(_05680_ ) );
INV_X1 _26477_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05681_ ) );
AND4_X1 _26478_ ( .A1(_05681_ ), .A2(_04217_ ), .A3(_04309_ ), .A4(_04175_ ), .ZN(_05682_ ) );
NOR3_X1 _26479_ ( .A1(_05653_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04549_ ), .ZN(_05683_ ) );
NOR3_X1 _26480_ ( .A1(_05680_ ), .A2(_05682_ ), .A3(_05683_ ), .ZN(_05684_ ) );
OR4_X1 _26481_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04179_ ), .A3(_04182_ ), .A4(_04184_ ), .ZN(_05685_ ) );
OR3_X1 _26482_ ( .A1(_04188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04549_ ), .ZN(_05686_ ) );
AND3_X1 _26483_ ( .A1(_05684_ ), .A2(_05685_ ), .A3(_05686_ ), .ZN(_05687_ ) );
INV_X1 _26484_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05688_ ) );
NAND4_X1 _26485_ ( .A1(_04552_ ), .A2(_04553_ ), .A3(_05688_ ), .A4(_04555_ ), .ZN(_05689_ ) );
OR3_X1 _26486_ ( .A1(_04326_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04819_ ), .ZN(_05690_ ) );
NAND3_X1 _26487_ ( .A1(_05687_ ), .A2(_05689_ ), .A3(_05690_ ), .ZN(_05691_ ) );
NOR4_X1 _26488_ ( .A1(_05554_ ), .A2(_04544_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04550_ ), .ZN(_05692_ ) );
NOR3_X1 _26489_ ( .A1(_05202_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04637_ ), .ZN(_05693_ ) );
NOR3_X1 _26490_ ( .A1(_05691_ ), .A2(_05692_ ), .A3(_05693_ ), .ZN(_05694_ ) );
INV_X1 _26491_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05695_ ) );
NAND3_X1 _26492_ ( .A1(_04562_ ), .A2(_05695_ ), .A3(_04224_ ), .ZN(_05696_ ) );
INV_X1 _26493_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05697_ ) );
OAI211_X1 _26494_ ( .A(_04221_ ), .B(_10792_ ), .C1(_05697_ ), .C2(_04555_ ), .ZN(_05698_ ) );
AND3_X1 _26495_ ( .A1(_05694_ ), .A2(_05696_ ), .A3(_05698_ ), .ZN(_05699_ ) );
AND3_X1 _26496_ ( .A1(_04221_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04242_ ), .ZN(_05700_ ) );
OR2_X1 _26497_ ( .A1(_04240_ ), .A2(_05700_ ), .ZN(_05701_ ) );
OAI22_X1 _26498_ ( .A1(_05642_ ), .A2(\idu.rs_reg ), .B1(_05699_ ), .B2(_05701_ ), .ZN(\idu.io_out_bits_rs1_data [6] ) );
AND2_X1 _26499_ ( .A1(_05637_ ), .A2(_05638_ ), .ZN(_05702_ ) );
INV_X1 _26500_ ( .A(_05702_ ), .ZN(\lsu.io_out_bits_rd_wdata [6] ) );
NAND3_X1 _26501_ ( .A1(_04571_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04243_ ), .ZN(_05703_ ) );
OR3_X1 _26502_ ( .A1(_04636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04637_ ), .ZN(_05704_ ) );
INV_X1 _26503_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05705_ ) );
AND4_X1 _26504_ ( .A1(_05705_ ), .A2(_04216_ ), .A3(_04151_ ), .A4(_04020_ ), .ZN(_05706_ ) );
INV_X1 _26505_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05707_ ) );
AND4_X1 _26506_ ( .A1(_05707_ ), .A2(_04109_ ), .A3(_04111_ ), .A4(_04513_ ), .ZN(_05708_ ) );
OR2_X1 _26507_ ( .A1(_05293_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05709_ ) );
OAI21_X1 _26508_ ( .A(_05709_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .B2(_04493_ ), .ZN(_05710_ ) );
INV_X1 _26509_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05711_ ) );
AOI21_X1 _26510_ ( .A(_05710_ ), .B1(_05711_ ), .B2(_04392_ ), .ZN(_05712_ ) );
OR2_X1 _26511_ ( .A1(_04070_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05713_ ) );
INV_X1 _26512_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05714_ ) );
NAND4_X1 _26513_ ( .A1(_04107_ ), .A2(_04154_ ), .A3(_05714_ ), .A4(_04080_ ), .ZN(_05715_ ) );
AND3_X1 _26514_ ( .A1(_05712_ ), .A2(_05713_ ), .A3(_05715_ ), .ZN(_05716_ ) );
OR3_X1 _26515_ ( .A1(_05372_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04127_ ), .ZN(_05717_ ) );
INV_X1 _26516_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05718_ ) );
NAND4_X1 _26517_ ( .A1(_04145_ ), .A2(_04858_ ), .A3(_05718_ ), .A4(_04282_ ), .ZN(_05719_ ) );
AND3_X1 _26518_ ( .A1(_05716_ ), .A2(_05717_ ), .A3(_05719_ ), .ZN(_05720_ ) );
OR3_X1 _26519_ ( .A1(_04592_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03994_ ), .ZN(_05721_ ) );
INV_X1 _26520_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05722_ ) );
NAND3_X1 _26521_ ( .A1(_04504_ ), .A2(_05722_ ), .A3(_04385_ ), .ZN(_05723_ ) );
NAND3_X1 _26522_ ( .A1(_05720_ ), .A2(_05721_ ), .A3(_05723_ ), .ZN(_05724_ ) );
INV_X1 _26523_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05725_ ) );
AND4_X1 _26524_ ( .A1(_05725_ ), .A2(_04331_ ), .A3(_04117_ ), .A4(_04598_ ), .ZN(_05726_ ) );
OAI21_X1 _26525_ ( .A(_04414_ ), .B1(_04102_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05727_ ) );
OR3_X1 _26526_ ( .A1(_05724_ ), .A2(_05726_ ), .A3(_05727_ ), .ZN(_05728_ ) );
NAND3_X1 _26527_ ( .A1(_04606_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04157_ ), .ZN(_05729_ ) );
AOI21_X1 _26528_ ( .A(_05708_ ), .B1(_05728_ ), .B2(_05729_ ), .ZN(_05730_ ) );
OR2_X1 _26529_ ( .A1(_05019_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05731_ ) );
NOR3_X1 _26530_ ( .A1(_04943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04254_ ), .ZN(_05732_ ) );
NOR2_X1 _26531_ ( .A1(_04292_ ), .A2(_05732_ ), .ZN(_05733_ ) );
NAND3_X1 _26532_ ( .A1(_05730_ ), .A2(_05731_ ), .A3(_05733_ ), .ZN(_05734_ ) );
NAND3_X1 _26533_ ( .A1(_04027_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04525_ ), .ZN(_05735_ ) );
AOI21_X1 _26534_ ( .A(_05706_ ), .B1(_05734_ ), .B2(_05735_ ), .ZN(_05736_ ) );
OR2_X1 _26535_ ( .A1(_04711_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05737_ ) );
INV_X1 _26536_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05738_ ) );
NAND4_X1 _26537_ ( .A1(_04241_ ), .A2(_04529_ ), .A3(_05738_ ), .A4(_04175_ ), .ZN(_05739_ ) );
NAND3_X1 _26538_ ( .A1(_05736_ ), .A2(_05737_ ), .A3(_05739_ ), .ZN(_05740_ ) );
NOR3_X1 _26539_ ( .A1(_04030_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04182_ ), .ZN(_05741_ ) );
INV_X1 _26540_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05742_ ) );
AND4_X1 _26541_ ( .A1(_05742_ ), .A2(_04216_ ), .A3(_04309_ ), .A4(_04310_ ), .ZN(_05743_ ) );
NOR3_X1 _26542_ ( .A1(_05740_ ), .A2(_05741_ ), .A3(_05743_ ), .ZN(_05744_ ) );
INV_X1 _26543_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05745_ ) );
NAND4_X1 _26544_ ( .A1(_04536_ ), .A2(_04615_ ), .A3(_05745_ ), .A4(_04538_ ), .ZN(_05746_ ) );
OR4_X1 _26545_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04316_ ), .A3(_04182_ ), .A4(_04184_ ), .ZN(_05747_ ) );
AND3_X1 _26546_ ( .A1(_05744_ ), .A2(_05746_ ), .A3(_05747_ ), .ZN(_05748_ ) );
OR3_X1 _26547_ ( .A1(_04548_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04327_ ), .ZN(_05749_ ) );
INV_X1 _26548_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05750_ ) );
NAND4_X1 _26549_ ( .A1(_04197_ ), .A2(_04194_ ), .A3(_05750_ ), .A4(_04199_ ), .ZN(_05751_ ) );
NAND3_X1 _26550_ ( .A1(_05748_ ), .A2(_05749_ ), .A3(_05751_ ), .ZN(_05752_ ) );
INV_X1 _26551_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05753_ ) );
AND4_X1 _26552_ ( .A1(_05753_ ), .A2(_04333_ ), .A3(_04615_ ), .A4(_04210_ ), .ZN(_05754_ ) );
OAI21_X1 _26553_ ( .A(_04447_ ), .B1(_04202_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05755_ ) );
NOR3_X1 _26554_ ( .A1(_05752_ ), .A2(_05754_ ), .A3(_05755_ ), .ZN(_05756_ ) );
AND3_X1 _26555_ ( .A1(_04444_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04633_ ), .ZN(_05757_ ) );
OAI21_X1 _26556_ ( .A(_05704_ ), .B1(_05756_ ), .B2(_05757_ ), .ZN(_05758_ ) );
AOI211_X1 _26557_ ( .A(_04015_ ), .B(_04023_ ), .C1(_04005_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05759_ ) );
OAI211_X1 _26558_ ( .A(_04247_ ), .B(_05703_ ), .C1(_05758_ ), .C2(_05759_ ), .ZN(_05760_ ) );
AOI21_X1 _26559_ ( .A(_03856_ ), .B1(_03105_ ), .B2(_03106_ ), .ZN(_05761_ ) );
NOR3_X1 _26560_ ( .A1(_03989_ ), .A2(_00484_ ), .A3(_04236_ ), .ZN(_05762_ ) );
OAI21_X1 _26561_ ( .A(fanout_net_1 ), .B1(_08562_ ), .B2(\io_master_rdata [5] ), .ZN(_05763_ ) );
AND4_X1 _26562_ ( .A1(fanout_net_1 ), .A2(_04982_ ), .A3(_04983_ ), .A4(lsu_io_out_bits_rd_wdata_$_MUX__Y_10_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05764_ ) );
OAI21_X1 _26563_ ( .A(_05498_ ), .B1(_05763_ ), .B2(_05764_ ), .ZN(_05765_ ) );
AOI22_X1 _26564_ ( .A1(_04368_ ), .A2(\io_master_awaddr [1] ), .B1(_03906_ ), .B2(_05059_ ), .ZN(_05766_ ) );
OAI211_X1 _26565_ ( .A(_05565_ ), .B(_05765_ ), .C1(_05766_ ), .C2(_04462_ ), .ZN(_05767_ ) );
NAND2_X1 _26566_ ( .A1(_03926_ ), .A2(\lsu.io_in_bits_rd_wdata [5] ), .ZN(_05768_ ) );
AND2_X1 _26567_ ( .A1(_05767_ ), .A2(_05768_ ), .ZN(_05769_ ) );
INV_X1 _26568_ ( .A(_05769_ ), .ZN(\lsu.io_out_bits_rd_wdata [5] ) );
MUX2_X1 _26569_ ( .A(_05762_ ), .B(\lsu.io_out_bits_rd_wdata [5] ), .S(_04340_ ), .Z(_05770_ ) );
AOI21_X1 _26570_ ( .A(_05761_ ), .B1(_04738_ ), .B2(_05770_ ), .ZN(_05771_ ) );
OAI21_X1 _26571_ ( .A(_05760_ ), .B1(_05771_ ), .B2(\idu.rs_reg ), .ZN(\idu.io_out_bits_rs1_data [5] ) );
AOI21_X1 _26572_ ( .A(_03856_ ), .B1(_03165_ ), .B2(_03166_ ), .ZN(_05772_ ) );
NOR3_X1 _26573_ ( .A1(_03989_ ), .A2(_00485_ ), .A3(_04236_ ), .ZN(_05773_ ) );
OAI21_X1 _26574_ ( .A(fanout_net_1 ), .B1(_08562_ ), .B2(\io_master_rdata [4] ), .ZN(_05774_ ) );
AND4_X1 _26575_ ( .A1(fanout_net_1 ), .A2(_04982_ ), .A3(_04983_ ), .A4(lsu_io_out_bits_rd_wdata_$_MUX__Y_11_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05775_ ) );
OAI21_X1 _26576_ ( .A(_05498_ ), .B1(_05774_ ), .B2(_05775_ ), .ZN(_05776_ ) );
AND3_X1 _26577_ ( .A1(_05136_ ), .A2(_03906_ ), .A3(_05137_ ), .ZN(_05777_ ) );
AOI21_X1 _26578_ ( .A(_05777_ ), .B1(_04473_ ), .B2(\io_master_awaddr [1] ), .ZN(_05778_ ) );
OAI211_X1 _26579_ ( .A(_05776_ ), .B(_05565_ ), .C1(_04462_ ), .C2(_05778_ ), .ZN(_05779_ ) );
NAND2_X1 _26580_ ( .A1(_03926_ ), .A2(\lsu.io_in_bits_rd_wdata [4] ), .ZN(_05780_ ) );
AND2_X1 _26581_ ( .A1(_05779_ ), .A2(_05780_ ), .ZN(_05781_ ) );
INV_X1 _26582_ ( .A(_05781_ ), .ZN(\lsu.io_out_bits_rd_wdata [4] ) );
MUX2_X1 _26583_ ( .A(_05773_ ), .B(\lsu.io_out_bits_rd_wdata [4] ), .S(_04340_ ), .Z(_05782_ ) );
AOI21_X1 _26584_ ( .A(_05772_ ), .B1(_04738_ ), .B2(_05782_ ), .ZN(_05783_ ) );
NAND3_X1 _26585_ ( .A1(_04207_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04211_ ), .ZN(_05784_ ) );
AOI211_X1 _26586_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_05325_ ), .C1(\idu.io_in_bits_inst [19] ), .C2(_11030_ ), .ZN(_05785_ ) );
OR3_X1 _26587_ ( .A1(_04263_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_03992_ ), .ZN(_05786_ ) );
OAI21_X1 _26588_ ( .A(_05786_ ), .B1(_05293_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05787_ ) );
NOR4_X1 _26589_ ( .A1(_04124_ ), .A2(_04918_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04016_ ), .ZN(_05788_ ) );
OR3_X1 _26590_ ( .A1(_05787_ ), .A2(_04068_ ), .A3(_05788_ ), .ZN(_05789_ ) );
NAND4_X1 _26591_ ( .A1(_04155_ ), .A2(_04037_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_11101_ ), .ZN(_05790_ ) );
AOI21_X1 _26592_ ( .A(_05785_ ), .B1(_05789_ ), .B2(_05790_ ), .ZN(_05791_ ) );
INV_X1 _26593_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05792_ ) );
NAND3_X1 _26594_ ( .A1(_04078_ ), .A2(_05792_ ), .A3(_04283_ ), .ZN(_05793_ ) );
INV_X1 _26595_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05794_ ) );
NAND4_X1 _26596_ ( .A1(_04145_ ), .A2(_04155_ ), .A3(_05794_ ), .A4(_04598_ ), .ZN(_05795_ ) );
NAND3_X1 _26597_ ( .A1(_05791_ ), .A2(_05793_ ), .A3(_05795_ ), .ZN(_05796_ ) );
NOR3_X1 _26598_ ( .A1(_04187_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04018_ ), .ZN(_05797_ ) );
NOR3_X1 _26599_ ( .A1(_05011_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04018_ ), .ZN(_05798_ ) );
NOR3_X1 _26600_ ( .A1(_05796_ ), .A2(_05797_ ), .A3(_05798_ ), .ZN(_05799_ ) );
OR3_X1 _26601_ ( .A1(_04095_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04163_ ), .ZN(_05800_ ) );
OR4_X1 _26602_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_05437_ ), .A3(_04125_ ), .A4(_04128_ ), .ZN(_05801_ ) );
NAND3_X1 _26603_ ( .A1(_05799_ ), .A2(_05800_ ), .A3(_05801_ ), .ZN(_05802_ ) );
INV_X1 _26604_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05803_ ) );
AND4_X1 _26605_ ( .A1(_05803_ ), .A2(_04036_ ), .A3(_04038_ ), .A4(_04513_ ), .ZN(_05804_ ) );
INV_X1 _26606_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05805_ ) );
AND4_X1 _26607_ ( .A1(_05805_ ), .A2(_04109_ ), .A3(_04036_ ), .A4(_04513_ ), .ZN(_05806_ ) );
NOR3_X1 _26608_ ( .A1(_05802_ ), .A2(_05804_ ), .A3(_05806_ ), .ZN(_05807_ ) );
OR2_X1 _26609_ ( .A1(_05019_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05808_ ) );
OR3_X1 _26610_ ( .A1(_04943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04173_ ), .ZN(_05809_ ) );
NAND3_X1 _26611_ ( .A1(_05807_ ), .A2(_05808_ ), .A3(_05809_ ), .ZN(_05810_ ) );
INV_X1 _26612_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05811_ ) );
AND4_X1 _26613_ ( .A1(_05811_ ), .A2(_04253_ ), .A3(_04157_ ), .A4(_04159_ ), .ZN(_05812_ ) );
NOR3_X1 _26614_ ( .A1(_04485_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04183_ ), .ZN(_05813_ ) );
NOR3_X1 _26615_ ( .A1(_05810_ ), .A2(_05812_ ), .A3(_05813_ ), .ZN(_05814_ ) );
OR2_X1 _26616_ ( .A1(_04711_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05815_ ) );
OR4_X1 _26617_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04178_ ), .A3(_04947_ ), .A4(_04437_ ), .ZN(_05816_ ) );
NAND3_X1 _26618_ ( .A1(_05814_ ), .A2(_05815_ ), .A3(_05816_ ), .ZN(_05817_ ) );
INV_X1 _26619_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05818_ ) );
AND4_X1 _26620_ ( .A1(_05818_ ), .A2(_04309_ ), .A3(_04158_ ), .A4(_04310_ ), .ZN(_05819_ ) );
NOR3_X1 _26621_ ( .A1(_05325_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04184_ ), .ZN(_05820_ ) );
NOR3_X1 _26622_ ( .A1(_05817_ ), .A2(_05819_ ), .A3(_05820_ ), .ZN(_05821_ ) );
OR3_X1 _26623_ ( .A1(_05653_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04191_ ), .ZN(_05822_ ) );
OR4_X1 _26624_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04316_ ), .A3(_04317_ ), .A4(_04318_ ), .ZN(_05823_ ) );
AND3_X1 _26625_ ( .A1(_05821_ ), .A2(_05822_ ), .A3(_05823_ ), .ZN(_05824_ ) );
OR3_X1 _26626_ ( .A1(_04188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04327_ ), .ZN(_05825_ ) );
INV_X1 _26627_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05826_ ) );
NAND4_X1 _26628_ ( .A1(_04197_ ), .A2(_04194_ ), .A3(_05826_ ), .A4(_04199_ ), .ZN(_05827_ ) );
NAND3_X1 _26629_ ( .A1(_05824_ ), .A2(_05825_ ), .A3(_05827_ ), .ZN(_05828_ ) );
OAI21_X1 _26630_ ( .A(_04558_ ), .B1(_04204_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05829_ ) );
OAI21_X1 _26631_ ( .A(_05784_ ), .B1(_05828_ ), .B2(_05829_ ), .ZN(_05830_ ) );
INV_X1 _26632_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05831_ ) );
NAND4_X1 _26633_ ( .A1(_04633_ ), .A2(_04621_ ), .A3(_05831_ ), .A4(_04212_ ), .ZN(_05832_ ) );
OR3_X1 _26634_ ( .A1(_04636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04637_ ), .ZN(_05833_ ) );
NAND4_X1 _26635_ ( .A1(_05830_ ), .A2(_05207_ ), .A3(_05832_ ), .A4(_05833_ ), .ZN(_05834_ ) );
NAND3_X1 _26636_ ( .A1(_04562_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04728_ ), .ZN(_05835_ ) );
AOI21_X1 _26637_ ( .A(_04250_ ), .B1(_05834_ ), .B2(_05835_ ), .ZN(_05836_ ) );
NAND3_X1 _26638_ ( .A1(_04571_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04243_ ), .ZN(_05837_ ) );
NAND2_X1 _26639_ ( .A1(_04247_ ), .A2(_05837_ ), .ZN(_05838_ ) );
OAI22_X1 _26640_ ( .A1(_05783_ ), .A2(\idu.rs_reg ), .B1(_05836_ ), .B2(_05838_ ), .ZN(\idu.io_out_bits_rs1_data [4] ) );
AOI21_X1 _26641_ ( .A(_03857_ ), .B1(_03225_ ), .B2(_03226_ ), .ZN(_05839_ ) );
OAI21_X1 _26642_ ( .A(\arbiter._io_axi_araddr_T ), .B1(_08562_ ), .B2(\io_master_rdata [3] ), .ZN(_05840_ ) );
AND4_X1 _26643_ ( .A1(\arbiter._io_axi_araddr_T ), .A2(_04982_ ), .A3(_04983_ ), .A4(lsu_io_out_bits_rd_wdata_$_MUX__Y_12_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05841_ ) );
OAI21_X1 _26644_ ( .A(_05498_ ), .B1(_05840_ ), .B2(_05841_ ), .ZN(_05842_ ) );
NOR2_X1 _26645_ ( .A1(_04650_ ), .A2(_03872_ ), .ZN(_05843_ ) );
AOI21_X1 _26646_ ( .A(_05843_ ), .B1(_03906_ ), .B2(_05280_ ), .ZN(_05844_ ) );
OAI211_X1 _26647_ ( .A(_05565_ ), .B(_05842_ ), .C1(_05844_ ), .C2(_04462_ ), .ZN(_05845_ ) );
NAND2_X1 _26648_ ( .A1(_03927_ ), .A2(\lsu.io_in_bits_rd_wdata [3] ), .ZN(_05846_ ) );
AND3_X1 _26649_ ( .A1(_05845_ ), .A2(_03925_ ), .A3(_05846_ ), .ZN(_05847_ ) );
NAND4_X1 _26650_ ( .A1(_03991_ ), .A2(\wbu.io_in_bits_rd_wdata [3] ), .A3(_03998_ ), .A4(_04011_ ), .ZN(_05848_ ) );
AOI211_X1 _26651_ ( .A(_03859_ ), .B(_05847_ ), .C1(_03932_ ), .C2(_05848_ ), .ZN(_05849_ ) );
OAI21_X1 _26652_ ( .A(_03850_ ), .B1(_05839_ ), .B2(_05849_ ), .ZN(_05850_ ) );
NAND3_X1 _26653_ ( .A1(_04207_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04211_ ), .ZN(_05851_ ) );
NOR3_X1 _26654_ ( .A1(_04485_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04190_ ), .ZN(_05852_ ) );
INV_X1 _26655_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_05853_ ) );
NAND3_X1 _26656_ ( .A1(_04134_ ), .A2(_05853_ ), .A3(_11099_ ), .ZN(_05854_ ) );
OAI21_X1 _26657_ ( .A(_05854_ ), .B1(_05293_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05855_ ) );
INV_X1 _26658_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05856_ ) );
AOI21_X1 _26659_ ( .A(_05855_ ), .B1(_05856_ ), .B2(_04392_ ), .ZN(_05857_ ) );
OR2_X1 _26660_ ( .A1(_04497_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05858_ ) );
INV_X1 _26661_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05859_ ) );
NAND4_X1 _26662_ ( .A1(_04107_ ), .A2(_04154_ ), .A3(_05859_ ), .A4(_11100_ ), .ZN(_05860_ ) );
AND3_X1 _26663_ ( .A1(_05857_ ), .A2(_05858_ ), .A3(_05860_ ), .ZN(_05861_ ) );
OR3_X1 _26664_ ( .A1(_05653_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04127_ ), .ZN(_05862_ ) );
INV_X1 _26665_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05863_ ) );
NAND4_X1 _26666_ ( .A1(_04145_ ), .A2(_04858_ ), .A3(_05863_ ), .A4(_11101_ ), .ZN(_05864_ ) );
NAND3_X1 _26667_ ( .A1(_05861_ ), .A2(_05862_ ), .A3(_05864_ ), .ZN(_05865_ ) );
NOR3_X1 _26668_ ( .A1(_04592_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04138_ ), .ZN(_05866_ ) );
INV_X1 _26669_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05867_ ) );
AND3_X1 _26670_ ( .A1(_04257_ ), .A2(_05867_ ), .A3(_04384_ ), .ZN(_05868_ ) );
NOR3_X1 _26671_ ( .A1(_05865_ ), .A2(_05866_ ), .A3(_05868_ ), .ZN(_05869_ ) );
INV_X1 _26672_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05870_ ) );
NAND4_X1 _26673_ ( .A1(_04509_ ), .A2(_04169_ ), .A3(_05870_ ), .A4(_04113_ ), .ZN(_05871_ ) );
OR4_X1 _26674_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_05437_ ), .A3(_04124_ ), .A4(_04017_ ), .ZN(_05872_ ) );
AND3_X1 _26675_ ( .A1(_05869_ ), .A2(_05871_ ), .A3(_05872_ ), .ZN(_05873_ ) );
OR3_X1 _26676_ ( .A1(_05201_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04163_ ), .ZN(_05874_ ) );
INV_X1 _26677_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05875_ ) );
NAND4_X1 _26678_ ( .A1(_04109_ ), .A2(_04111_ ), .A3(_05875_ ), .A4(_04114_ ), .ZN(_05876_ ) );
NAND3_X1 _26679_ ( .A1(_05873_ ), .A2(_05874_ ), .A3(_05876_ ), .ZN(_05877_ ) );
INV_X1 _26680_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05878_ ) );
AND4_X1 _26681_ ( .A1(_05878_ ), .A2(_04119_ ), .A3(_04111_ ), .A4(_04513_ ), .ZN(_05879_ ) );
INV_X1 _26682_ ( .A(_04292_ ), .ZN(_05880_ ) );
OAI21_X1 _26683_ ( .A(_05880_ ), .B1(_04707_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05881_ ) );
OR3_X1 _26684_ ( .A1(_05877_ ), .A2(_05879_ ), .A3(_05881_ ), .ZN(_05882_ ) );
NAND3_X1 _26685_ ( .A1(_04027_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04525_ ), .ZN(_05883_ ) );
AOI21_X1 _26686_ ( .A(_05852_ ), .B1(_05882_ ), .B2(_05883_ ), .ZN(_05884_ ) );
INV_X1 _26687_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05885_ ) );
NAND4_X1 _26688_ ( .A1(_04528_ ), .A2(_04529_ ), .A3(_05885_ ), .A4(_04209_ ), .ZN(_05886_ ) );
OR4_X1 _26689_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04178_ ), .A3(_04947_ ), .A4(_04183_ ), .ZN(_05887_ ) );
NAND3_X1 _26690_ ( .A1(_05884_ ), .A2(_05886_ ), .A3(_05887_ ), .ZN(_05888_ ) );
INV_X1 _26691_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05889_ ) );
AND4_X1 _26692_ ( .A1(_05889_ ), .A2(_04309_ ), .A3(_04158_ ), .A4(_04175_ ), .ZN(_05890_ ) );
INV_X1 _26693_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05891_ ) );
AND4_X1 _26694_ ( .A1(_05891_ ), .A2(_04217_ ), .A3(_04309_ ), .A4(_04313_ ), .ZN(_05892_ ) );
NOR3_X1 _26695_ ( .A1(_05888_ ), .A2(_05890_ ), .A3(_05892_ ), .ZN(_05893_ ) );
OR3_X1 _26696_ ( .A1(_05653_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04549_ ), .ZN(_05894_ ) );
OR4_X1 _26697_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04316_ ), .A3(_04182_ ), .A4(_04184_ ), .ZN(_05895_ ) );
AND3_X1 _26698_ ( .A1(_05893_ ), .A2(_05894_ ), .A3(_05895_ ), .ZN(_05896_ ) );
INV_X1 _26699_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05897_ ) );
NAND4_X1 _26700_ ( .A1(_04620_ ), .A2(_04621_ ), .A3(_05897_ ), .A4(_04211_ ), .ZN(_05898_ ) );
INV_X1 _26701_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05899_ ) );
NAND4_X1 _26702_ ( .A1(_04197_ ), .A2(_04194_ ), .A3(_05899_ ), .A4(_04455_ ), .ZN(_05900_ ) );
NAND3_X1 _26703_ ( .A1(_05896_ ), .A2(_05898_ ), .A3(_05900_ ), .ZN(_05901_ ) );
OAI21_X1 _26704_ ( .A(_04558_ ), .B1(_04204_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05902_ ) );
OAI21_X1 _26705_ ( .A(_05851_ ), .B1(_05901_ ), .B2(_05902_ ), .ZN(_05903_ ) );
INV_X1 _26706_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05904_ ) );
NAND4_X1 _26707_ ( .A1(_04633_ ), .A2(_04621_ ), .A3(_05904_ ), .A4(_04212_ ), .ZN(_05905_ ) );
OR3_X1 _26708_ ( .A1(_04636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04637_ ), .ZN(_05906_ ) );
NAND4_X1 _26709_ ( .A1(_05903_ ), .A2(_05207_ ), .A3(_05905_ ), .A4(_05906_ ), .ZN(_05907_ ) );
NAND3_X1 _26710_ ( .A1(_04222_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04728_ ), .ZN(_05908_ ) );
AOI21_X1 _26711_ ( .A(_04250_ ), .B1(_05907_ ), .B2(_05908_ ), .ZN(_05909_ ) );
NAND3_X1 _26712_ ( .A1(_04222_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04482_ ), .ZN(_05910_ ) );
NAND2_X1 _26713_ ( .A1(_04481_ ), .A2(_05910_ ), .ZN(_05911_ ) );
OAI21_X1 _26714_ ( .A(_05850_ ), .B1(_05909_ ), .B2(_05911_ ), .ZN(\idu.io_out_bits_rs1_data [3] ) );
AND2_X1 _26715_ ( .A1(_05845_ ), .A2(_05846_ ), .ZN(_05912_ ) );
INV_X1 _26716_ ( .A(_05912_ ), .ZN(\lsu.io_out_bits_rd_wdata [3] ) );
NOR3_X1 _26717_ ( .A1(_03284_ ), .A2(_03285_ ), .A3(_03856_ ), .ZN(_05913_ ) );
OAI21_X1 _26718_ ( .A(\arbiter._io_axi_araddr_T ), .B1(_08562_ ), .B2(\io_master_rdata [2] ), .ZN(_05914_ ) );
AND4_X1 _26719_ ( .A1(\arbiter._io_axi_araddr_T ), .A2(_04982_ ), .A3(_04983_ ), .A4(lsu_io_out_bits_rd_wdata_$_MUX__Y_13_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05915_ ) );
OAI21_X1 _26720_ ( .A(_05498_ ), .B1(_05914_ ), .B2(_05915_ ), .ZN(_05916_ ) );
AOI22_X1 _26721_ ( .A1(_04669_ ), .A2(\io_master_awaddr [1] ), .B1(_03906_ ), .B2(_05353_ ), .ZN(_05917_ ) );
OAI211_X1 _26722_ ( .A(_05916_ ), .B(_05565_ ), .C1(_05917_ ), .C2(_04462_ ), .ZN(_05918_ ) );
NAND2_X1 _26723_ ( .A1(_03927_ ), .A2(\lsu.io_in_bits_rd_wdata [2] ), .ZN(_05919_ ) );
AND3_X1 _26724_ ( .A1(_05918_ ), .A2(_03925_ ), .A3(_05919_ ), .ZN(_05920_ ) );
NAND4_X1 _26725_ ( .A1(_03991_ ), .A2(\wbu.io_in_bits_rd_wdata [2] ), .A3(_03998_ ), .A4(_04011_ ), .ZN(_05921_ ) );
AOI211_X1 _26726_ ( .A(_03859_ ), .B(_05920_ ), .C1(_03932_ ), .C2(_05921_ ), .ZN(_05922_ ) );
OAI21_X1 _26727_ ( .A(_03850_ ), .B1(_05913_ ), .B2(_05922_ ), .ZN(_05923_ ) );
NAND3_X1 _26728_ ( .A1(_04444_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04529_ ), .ZN(_05924_ ) );
INV_X1 _26729_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05925_ ) );
NAND3_X1 _26730_ ( .A1(_04504_ ), .A2(_05925_ ), .A3(_04038_ ), .ZN(_05926_ ) );
INV_X1 _26731_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05927_ ) );
AND4_X1 _26732_ ( .A1(_05927_ ), .A2(_04403_ ), .A3(_04116_ ), .A4(_04080_ ), .ZN(_05928_ ) );
OR2_X1 _26733_ ( .A1(_04083_ ), .A2(_05928_ ), .ZN(_05929_ ) );
NAND4_X1 _26734_ ( .A1(_04858_ ), .A2(_04026_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04041_ ), .ZN(_05930_ ) );
INV_X1 _26735_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05931_ ) );
NAND4_X1 _26736_ ( .A1(_04144_ ), .A2(_04149_ ), .A3(_05931_ ), .A4(_04080_ ), .ZN(_05932_ ) );
NOR3_X1 _26737_ ( .A1(_04294_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_03992_ ), .ZN(_05933_ ) );
NOR2_X1 _26738_ ( .A1(_04053_ ), .A2(_05933_ ), .ZN(_05934_ ) );
AND4_X1 _26739_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04116_ ), .A3(_04148_ ), .A4(_04399_ ), .ZN(_05935_ ) );
OAI21_X1 _26740_ ( .A(_05932_ ), .B1(_05934_ ), .B2(_05935_ ), .ZN(_05936_ ) );
OAI21_X1 _26741_ ( .A(_05930_ ), .B1(_05936_ ), .B2(_04068_ ), .ZN(_05937_ ) );
NAND2_X1 _26742_ ( .A1(_05937_ ), .A2(_04496_ ), .ZN(_05938_ ) );
NAND4_X1 _26743_ ( .A1(_04108_ ), .A2(_04155_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04042_ ), .ZN(_05939_ ) );
AOI21_X1 _26744_ ( .A(_05929_ ), .B1(_05938_ ), .B2(_05939_ ), .ZN(_05940_ ) );
AND3_X1 _26745_ ( .A1(_04082_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04042_ ), .ZN(_05941_ ) );
OAI21_X1 _26746_ ( .A(_05926_ ), .B1(_05940_ ), .B2(_05941_ ), .ZN(_05942_ ) );
NOR3_X1 _26747_ ( .A1(_05011_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04163_ ), .ZN(_05943_ ) );
INV_X1 _26748_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05944_ ) );
AND4_X1 _26749_ ( .A1(_05944_ ), .A2(_04331_ ), .A3(_04118_ ), .A4(_04598_ ), .ZN(_05945_ ) );
OR3_X1 _26750_ ( .A1(_05942_ ), .A2(_05943_ ), .A3(_05945_ ), .ZN(_05946_ ) );
INV_X1 _26751_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05947_ ) );
AND4_X1 _26752_ ( .A1(_05947_ ), .A2(_04509_ ), .A3(_04146_ ), .A4(_04114_ ), .ZN(_05948_ ) );
NOR3_X1 _26753_ ( .A1(_05201_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04254_ ), .ZN(_05949_ ) );
NOR3_X1 _26754_ ( .A1(_05946_ ), .A2(_05948_ ), .A3(_05949_ ), .ZN(_05950_ ) );
OR3_X1 _26755_ ( .A1(_04519_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04254_ ), .ZN(_05951_ ) );
INV_X1 _26756_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05952_ ) );
NAND4_X1 _26757_ ( .A1(_04297_ ), .A2(_04445_ ), .A3(_05952_ ), .A4(_04183_ ), .ZN(_05953_ ) );
NAND3_X1 _26758_ ( .A1(_05950_ ), .A2(_05951_ ), .A3(_05953_ ), .ZN(_05954_ ) );
OAI21_X1 _26759_ ( .A(_05880_ ), .B1(_04707_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05955_ ) );
OAI21_X1 _26760_ ( .A(_05924_ ), .B1(_05954_ ), .B2(_05955_ ), .ZN(_05956_ ) );
OR3_X1 _26761_ ( .A1(_04485_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04318_ ), .ZN(_05957_ ) );
INV_X1 _26762_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05958_ ) );
NAND4_X1 _26763_ ( .A1(_04528_ ), .A2(_04529_ ), .A3(_05958_ ), .A4(_04209_ ), .ZN(_05959_ ) );
NAND3_X1 _26764_ ( .A1(_05956_ ), .A2(_05957_ ), .A3(_05959_ ), .ZN(_05960_ ) );
INV_X1 _26765_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05961_ ) );
AND4_X1 _26766_ ( .A1(_05961_ ), .A2(_04241_ ), .A3(_04529_ ), .A4(_04175_ ), .ZN(_05962_ ) );
NOR3_X1 _26767_ ( .A1(_04030_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04534_ ), .ZN(_05963_ ) );
NOR3_X1 _26768_ ( .A1(_05960_ ), .A2(_05962_ ), .A3(_05963_ ), .ZN(_05964_ ) );
OR3_X1 _26769_ ( .A1(_05325_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04549_ ), .ZN(_05965_ ) );
INV_X1 _26770_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05966_ ) );
NAND4_X1 _26771_ ( .A1(_04536_ ), .A2(_04615_ ), .A3(_05966_ ), .A4(_04210_ ), .ZN(_05967_ ) );
NAND3_X1 _26772_ ( .A1(_05964_ ), .A2(_05965_ ), .A3(_05967_ ), .ZN(_05968_ ) );
NOR4_X1 _26773_ ( .A1(_04544_ ), .A2(_04534_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04327_ ), .ZN(_05969_ ) );
NOR3_X1 _26774_ ( .A1(_04548_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04550_ ), .ZN(_05970_ ) );
NOR3_X1 _26775_ ( .A1(_05968_ ), .A2(_05969_ ), .A3(_05970_ ), .ZN(_05971_ ) );
INV_X1 _26776_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05972_ ) );
NAND4_X1 _26777_ ( .A1(_04552_ ), .A2(_04553_ ), .A3(_05972_ ), .A4(_04555_ ), .ZN(_05973_ ) );
OR3_X1 _26778_ ( .A1(_04326_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04550_ ), .ZN(_05974_ ) );
AND3_X1 _26779_ ( .A1(_05971_ ), .A2(_05973_ ), .A3(_05974_ ), .ZN(_05975_ ) );
OR4_X1 _26780_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_05554_ ), .A3(_04544_ ), .A4(_04637_ ), .ZN(_05976_ ) );
INV_X1 _26781_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05977_ ) );
NAND4_X1 _26782_ ( .A1(_04633_ ), .A2(_04621_ ), .A3(_05977_ ), .A4(_04212_ ), .ZN(_05978_ ) );
NAND3_X1 _26783_ ( .A1(_05975_ ), .A2(_05976_ ), .A3(_05978_ ), .ZN(_05979_ ) );
INV_X1 _26784_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05980_ ) );
AND3_X1 _26785_ ( .A1(_04221_ ), .A2(_05980_ ), .A3(_04224_ ), .ZN(_05981_ ) );
AOI211_X1 _26786_ ( .A(_04015_ ), .B(_04023_ ), .C1(_04005_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05982_ ) );
NOR3_X1 _26787_ ( .A1(_05979_ ), .A2(_05981_ ), .A3(_05982_ ), .ZN(_05983_ ) );
NAND3_X1 _26788_ ( .A1(_04222_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04482_ ), .ZN(_05984_ ) );
NAND2_X1 _26789_ ( .A1(_04481_ ), .A2(_05984_ ), .ZN(_05985_ ) );
OAI21_X1 _26790_ ( .A(_05923_ ), .B1(_05983_ ), .B2(_05985_ ), .ZN(\idu.io_out_bits_rs1_data [2] ) );
AND2_X1 _26791_ ( .A1(_05918_ ), .A2(_05919_ ), .ZN(_05986_ ) );
INV_X1 _26792_ ( .A(_05986_ ), .ZN(\lsu.io_out_bits_rd_wdata [2] ) );
NAND2_X1 _26793_ ( .A1(_05213_ ), .A2(_05214_ ), .ZN(\lsu.io_out_bits_rd_wdata [29] ) );
NAND3_X1 _26794_ ( .A1(_05131_ ), .A2(\arbiter._io_axi_araddr_T ), .A3(\arbiter.io_lsu_arsize [1] ), .ZN(_05987_ ) );
OAI21_X1 _26795_ ( .A(_04642_ ), .B1(_03899_ ), .B2(_05987_ ), .ZN(_05988_ ) );
OAI21_X1 _26796_ ( .A(\lsu.io_in_bits_ren ), .B1(_05988_ ), .B2(_03916_ ), .ZN(_05989_ ) );
NAND2_X1 _26797_ ( .A1(_03926_ ), .A2(\lsu.io_in_bits_rd_wdata [28] ), .ZN(_05990_ ) );
NAND2_X1 _26798_ ( .A1(_05989_ ), .A2(_05990_ ), .ZN(\lsu.io_out_bits_rd_wdata [28] ) );
NAND2_X1 _26799_ ( .A1(\lsu.io_out_bits_rd_wdata [28] ), .A2(_04340_ ), .ZN(_05991_ ) );
OAI211_X1 _26800_ ( .A(\wbu.io_in_bits_rd_wdata [28] ), .B(_04656_ ), .C1(_08570_ ), .C2(_04658_ ), .ZN(_05992_ ) );
AOI21_X1 _26801_ ( .A(_04228_ ), .B1(_05991_ ), .B2(_05992_ ), .ZN(_05993_ ) );
AOI21_X1 _26802_ ( .A(_05993_ ), .B1(\exu.io_out_bits_rd_wdata [28] ), .B2(_04459_ ), .ZN(_05994_ ) );
NOR2_X1 _26803_ ( .A1(_05994_ ), .A2(\idu.rs_reg ), .ZN(_05995_ ) );
NOR3_X1 _26804_ ( .A1(_04028_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04946_ ), .ZN(_05996_ ) );
AND4_X1 _26805_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04057_ ), .A3(_04074_ ), .A4(_11098_ ), .ZN(_05997_ ) );
OR3_X1 _26806_ ( .A1(_04262_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10766_ ), .ZN(_05998_ ) );
MUX2_X1 _26807_ ( .A(_05998_ ), .B(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(_04053_ ), .Z(_05999_ ) );
MUX2_X1 _26808_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_05999_ ), .S(_04064_ ), .Z(_06000_ ) );
OR2_X1 _26809_ ( .A1(_04069_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06001_ ) );
AND2_X1 _26810_ ( .A1(_06000_ ), .A2(_06001_ ), .ZN(_06002_ ) );
AOI21_X1 _26811_ ( .A(_05997_ ), .B1(_06002_ ), .B2(_04496_ ), .ZN(_06003_ ) );
INV_X1 _26812_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06004_ ) );
AND4_X1 _26813_ ( .A1(_06004_ ), .A2(_04074_ ), .A3(_04116_ ), .A4(_04039_ ), .ZN(_06005_ ) );
OAI21_X1 _26814_ ( .A(_04090_ ), .B1(_04084_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06006_ ) );
NOR3_X1 _26815_ ( .A1(_06003_ ), .A2(_06005_ ), .A3(_06006_ ), .ZN(_06007_ ) );
AND3_X1 _26816_ ( .A1(_04088_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04026_ ), .ZN(_06008_ ) );
NOR2_X1 _26817_ ( .A1(_06007_ ), .A2(_06008_ ), .ZN(_06009_ ) );
NOR3_X1 _26818_ ( .A1(_05011_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04127_ ), .ZN(_06010_ ) );
NOR3_X1 _26819_ ( .A1(_04095_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03993_ ), .ZN(_06011_ ) );
NOR3_X1 _26820_ ( .A1(_06009_ ), .A2(_06010_ ), .A3(_06011_ ), .ZN(_06012_ ) );
OR4_X1 _26821_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_05437_ ), .A3(_04124_ ), .A4(_04016_ ), .ZN(_06013_ ) );
INV_X1 _26822_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06014_ ) );
NAND4_X1 _26823_ ( .A1(_04032_ ), .A2(_04037_ ), .A3(_06014_ ), .A4(_04282_ ), .ZN(_06015_ ) );
NAND3_X1 _26824_ ( .A1(_06012_ ), .A2(_06013_ ), .A3(_06015_ ), .ZN(_06016_ ) );
INV_X1 _26825_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06017_ ) );
AND4_X1 _26826_ ( .A1(_06017_ ), .A2(_04384_ ), .A3(_04032_ ), .A4(_04411_ ), .ZN(_06018_ ) );
OAI21_X1 _26827_ ( .A(_04707_ ), .B1(_04703_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06019_ ) );
OR3_X1 _26828_ ( .A1(_06016_ ), .A2(_06018_ ), .A3(_06019_ ), .ZN(_06020_ ) );
NAND3_X1 _26829_ ( .A1(_04606_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04146_ ), .ZN(_06021_ ) );
AOI21_X1 _26830_ ( .A(_05996_ ), .B1(_06020_ ), .B2(_06021_ ), .ZN(_06022_ ) );
OR3_X1 _26831_ ( .A1(_04294_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04043_ ), .ZN(_06023_ ) );
INV_X1 _26832_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06024_ ) );
NAND4_X1 _26833_ ( .A1(_04119_ ), .A2(_04253_ ), .A3(_06024_ ), .A4(_04173_ ), .ZN(_06025_ ) );
NAND3_X1 _26834_ ( .A1(_06022_ ), .A2(_06023_ ), .A3(_06025_ ), .ZN(_06026_ ) );
NOR4_X1 _26835_ ( .A1(_04126_ ), .A2(_04946_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04189_ ), .ZN(_06027_ ) );
NOR3_X1 _26836_ ( .A1(_04131_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04181_ ), .ZN(_06028_ ) );
NOR3_X1 _26837_ ( .A1(_06026_ ), .A2(_06027_ ), .A3(_06028_ ), .ZN(_06029_ ) );
INV_X1 _26838_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06030_ ) );
NAND4_X1 _26839_ ( .A1(_04216_ ), .A2(_04156_ ), .A3(_06030_ ), .A4(_04208_ ), .ZN(_06031_ ) );
INV_X1 _26840_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06032_ ) );
NAND4_X1 _26841_ ( .A1(_04167_ ), .A2(_04297_ ), .A3(_06032_ ), .A4(_04174_ ), .ZN(_06033_ ) );
NAND3_X1 _26842_ ( .A1(_06029_ ), .A2(_06031_ ), .A3(_06033_ ), .ZN(_06034_ ) );
NOR4_X1 _26843_ ( .A1(_04178_ ), .A2(_04317_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04183_ ), .ZN(_06035_ ) );
NOR3_X1 _26844_ ( .A1(_04187_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04190_ ), .ZN(_06036_ ) );
NOR3_X1 _26845_ ( .A1(_06034_ ), .A2(_06035_ ), .A3(_06036_ ), .ZN(_06037_ ) );
INV_X1 _26846_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06038_ ) );
NAND4_X1 _26847_ ( .A1(_04196_ ), .A2(_04000_ ), .A3(_06038_ ), .A4(_10756_ ), .ZN(_06039_ ) );
INV_X1 _26848_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06040_ ) );
AOI22_X1 _26849_ ( .A1(_04203_ ), .A2(_06040_ ), .B1(_04175_ ), .B2(_04207_ ), .ZN(_06041_ ) );
AND3_X1 _26850_ ( .A1(_06037_ ), .A2(_06039_ ), .A3(_06041_ ), .ZN(_06042_ ) );
AND3_X1 _26851_ ( .A1(_04207_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04842_ ), .ZN(_06043_ ) );
NOR2_X1 _26852_ ( .A1(_06042_ ), .A2(_06043_ ), .ZN(_06044_ ) );
INV_X1 _26853_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06045_ ) );
AND4_X1 _26854_ ( .A1(_06045_ ), .A2(_04445_ ), .A3(_04451_ ), .A4(_04623_ ), .ZN(_06046_ ) );
NOR3_X1 _26855_ ( .A1(_04519_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04327_ ), .ZN(_06047_ ) );
NOR3_X1 _26856_ ( .A1(_06044_ ), .A2(_06046_ ), .A3(_06047_ ), .ZN(_06048_ ) );
NOR4_X1 _26857_ ( .A1(_04022_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10595_ ), .A4(_04199_ ), .ZN(_06049_ ) );
NOR2_X1 _26858_ ( .A1(_06049_ ), .A2(_04249_ ), .ZN(_06050_ ) );
AOI221_X4 _26859_ ( .A(_04239_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B2(_04250_ ), .C1(_06048_ ), .C2(_06050_ ), .ZN(_06051_ ) );
OR2_X1 _26860_ ( .A1(_05995_ ), .A2(_06051_ ), .ZN(\idu.io_out_bits_rs1_data [28] ) );
NOR3_X1 _26861_ ( .A1(_03385_ ), .A2(_03386_ ), .A3(_04738_ ), .ZN(_06052_ ) );
OAI21_X1 _26862_ ( .A(\arbiter._io_axi_araddr_T ), .B1(_08562_ ), .B2(\io_master_rdata [1] ), .ZN(_06053_ ) );
AND4_X1 _26863_ ( .A1(\arbiter._io_axi_araddr_T ), .A2(_04982_ ), .A3(_04983_ ), .A4(lsu_io_out_bits_rd_wdata_$_MUX__Y_14_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06054_ ) );
OAI21_X1 _26864_ ( .A(_05498_ ), .B1(_06053_ ), .B2(_06054_ ), .ZN(_06055_ ) );
AOI22_X1 _26865_ ( .A1(_04759_ ), .A2(\io_master_awaddr [1] ), .B1(_03906_ ), .B2(_05427_ ), .ZN(_06056_ ) );
OAI211_X1 _26866_ ( .A(_05565_ ), .B(_06055_ ), .C1(_06056_ ), .C2(_04462_ ), .ZN(_06057_ ) );
NAND2_X1 _26867_ ( .A1(_03927_ ), .A2(\lsu.io_in_bits_rd_wdata [1] ), .ZN(_06058_ ) );
AND2_X1 _26868_ ( .A1(_06057_ ), .A2(_06058_ ), .ZN(_06059_ ) );
OR2_X1 _26869_ ( .A1(_06059_ ), .A2(_03931_ ), .ZN(_06060_ ) );
OAI211_X1 _26870_ ( .A(\wbu.io_in_bits_rd_wdata [1] ), .B(_04656_ ), .C1(_04657_ ), .C2(_04658_ ), .ZN(_06061_ ) );
AOI21_X1 _26871_ ( .A(_04459_ ), .B1(_06060_ ), .B2(_06061_ ), .ZN(_06062_ ) );
OAI21_X1 _26872_ ( .A(_03851_ ), .B1(_06052_ ), .B2(_06062_ ), .ZN(_06063_ ) );
NAND3_X1 _26873_ ( .A1(_04571_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04482_ ), .ZN(_06064_ ) );
NAND3_X1 _26874_ ( .A1(_04207_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04212_ ), .ZN(_06065_ ) );
NOR4_X1 _26875_ ( .A1(_04544_ ), .A2(_04534_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04545_ ), .ZN(_06066_ ) );
INV_X1 _26876_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06067_ ) );
NAND4_X1 _26877_ ( .A1(_04217_ ), .A2(_04529_ ), .A3(_06067_ ), .A4(_04313_ ), .ZN(_06068_ ) );
NAND3_X1 _26878_ ( .A1(_04606_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04147_ ), .ZN(_06069_ ) );
NOR4_X1 _26879_ ( .A1(_05554_ ), .A2(_04125_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04018_ ), .ZN(_06070_ ) );
INV_X1 _26880_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_06071_ ) );
NAND3_X1 _26881_ ( .A1(_04134_ ), .A2(_06071_ ), .A3(_04040_ ), .ZN(_06072_ ) );
OAI21_X1 _26882_ ( .A(_06072_ ), .B1(_05293_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06073_ ) );
NOR2_X1 _26883_ ( .A1(_04497_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06074_ ) );
INV_X1 _26884_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06075_ ) );
AND4_X1 _26885_ ( .A1(_06075_ ), .A2(_04098_ ), .A3(_04148_ ), .A4(_11099_ ), .ZN(_06076_ ) );
NOR3_X1 _26886_ ( .A1(_06073_ ), .A2(_06074_ ), .A3(_06076_ ), .ZN(_06077_ ) );
INV_X1 _26887_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06078_ ) );
NAND4_X1 _26888_ ( .A1(_04107_ ), .A2(_04154_ ), .A3(_06078_ ), .A4(_04041_ ), .ZN(_06079_ ) );
OR3_X1 _26889_ ( .A1(_05372_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04016_ ), .ZN(_06080_ ) );
AND3_X1 _26890_ ( .A1(_06077_ ), .A2(_06079_ ), .A3(_06080_ ), .ZN(_06081_ ) );
INV_X1 _26891_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06082_ ) );
NAND4_X1 _26892_ ( .A1(_04145_ ), .A2(_04155_ ), .A3(_06082_ ), .A4(_04042_ ), .ZN(_06083_ ) );
AND2_X1 _26893_ ( .A1(_06081_ ), .A2(_06083_ ), .ZN(_06084_ ) );
OR3_X1 _26894_ ( .A1(_04592_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04138_ ), .ZN(_06085_ ) );
INV_X1 _26895_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06086_ ) );
AOI22_X1 _26896_ ( .A1(_06086_ ), .A2(_04092_ ), .B1(_04048_ ), .B2(_04283_ ), .ZN(_06087_ ) );
NAND3_X1 _26897_ ( .A1(_06084_ ), .A2(_06085_ ), .A3(_06087_ ), .ZN(_06088_ ) );
NAND3_X1 _26898_ ( .A1(_04048_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04513_ ), .ZN(_06089_ ) );
AOI21_X1 _26899_ ( .A(_06070_ ), .B1(_06088_ ), .B2(_06089_ ), .ZN(_06090_ ) );
OR3_X1 _26900_ ( .A1(_05201_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04129_ ), .ZN(_06091_ ) );
INV_X1 _26901_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06092_ ) );
NAND4_X1 _26902_ ( .A1(_04936_ ), .A2(_04522_ ), .A3(_06092_ ), .A4(_04189_ ), .ZN(_06093_ ) );
NAND3_X1 _26903_ ( .A1(_06090_ ), .A2(_06091_ ), .A3(_06093_ ), .ZN(_06094_ ) );
OAI21_X1 _26904_ ( .A(_04707_ ), .B1(_05019_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06095_ ) );
OAI21_X1 _26905_ ( .A(_06069_ ), .B1(_06094_ ), .B2(_06095_ ), .ZN(_06096_ ) );
AND2_X1 _26906_ ( .A1(_06096_ ), .A2(_05880_ ), .ZN(_06097_ ) );
AND4_X1 _26907_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04525_ ), .A3(_04158_ ), .A4(_04208_ ), .ZN(_06098_ ) );
OAI21_X1 _26908_ ( .A(_06068_ ), .B1(_06097_ ), .B2(_06098_ ), .ZN(_06099_ ) );
NOR2_X1 _26909_ ( .A1(_04711_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06100_ ) );
NOR4_X1 _26910_ ( .A1(_04316_ ), .A2(_04947_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04318_ ), .ZN(_06101_ ) );
NOR3_X1 _26911_ ( .A1(_06099_ ), .A2(_06100_ ), .A3(_06101_ ), .ZN(_06102_ ) );
INV_X1 _26912_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06103_ ) );
NAND4_X1 _26913_ ( .A1(_04542_ ), .A2(_04451_ ), .A3(_06103_ ), .A4(_04538_ ), .ZN(_06104_ ) );
INV_X1 _26914_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06105_ ) );
NAND4_X1 _26915_ ( .A1(_04223_ ), .A2(_04542_ ), .A3(_06105_ ), .A4(_04623_ ), .ZN(_06106_ ) );
NAND4_X1 _26916_ ( .A1(_06102_ ), .A2(_04435_ ), .A3(_06104_ ), .A4(_06106_ ), .ZN(_06107_ ) );
NAND4_X1 _26917_ ( .A1(_04536_ ), .A2(_04615_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04210_ ), .ZN(_06108_ ) );
AOI21_X1 _26918_ ( .A(_06066_ ), .B1(_06107_ ), .B2(_06108_ ), .ZN(_06109_ ) );
INV_X1 _26919_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06110_ ) );
NAND4_X1 _26920_ ( .A1(_04620_ ), .A2(_04621_ ), .A3(_06110_ ), .A4(_04211_ ), .ZN(_06111_ ) );
INV_X1 _26921_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06112_ ) );
NAND4_X1 _26922_ ( .A1(_04552_ ), .A2(_04553_ ), .A3(_06112_ ), .A4(_04555_ ), .ZN(_06113_ ) );
NAND3_X1 _26923_ ( .A1(_06109_ ), .A2(_06111_ ), .A3(_06113_ ), .ZN(_06114_ ) );
OAI21_X1 _26924_ ( .A(_04558_ ), .B1(_04204_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06115_ ) );
OAI21_X1 _26925_ ( .A(_06065_ ), .B1(_06114_ ), .B2(_06115_ ), .ZN(_06116_ ) );
INV_X1 _26926_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06117_ ) );
NAND4_X1 _26927_ ( .A1(_04633_ ), .A2(_04621_ ), .A3(_06117_ ), .A4(_04212_ ), .ZN(_06118_ ) );
OR3_X1 _26928_ ( .A1(_04636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04820_ ), .ZN(_06119_ ) );
NAND3_X1 _26929_ ( .A1(_06116_ ), .A2(_06118_ ), .A3(_06119_ ), .ZN(_06120_ ) );
AOI211_X1 _26930_ ( .A(_04566_ ), .B(_04567_ ), .C1(_04568_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06121_ ) );
OAI211_X1 _26931_ ( .A(_04481_ ), .B(_06064_ ), .C1(_06120_ ), .C2(_06121_ ), .ZN(_06122_ ) );
NAND2_X1 _26932_ ( .A1(_06063_ ), .A2(_06122_ ), .ZN(\idu.io_out_bits_rs1_data [1] ) );
INV_X1 _26933_ ( .A(_06059_ ), .ZN(\lsu.io_out_bits_rd_wdata [1] ) );
AOI21_X1 _26934_ ( .A(_03857_ ), .B1(_03524_ ), .B2(_03525_ ), .ZN(_06123_ ) );
OAI21_X1 _26935_ ( .A(\arbiter._io_axi_araddr_T ), .B1(_08562_ ), .B2(\io_master_rdata [0] ), .ZN(_06124_ ) );
AND4_X1 _26936_ ( .A1(\arbiter._io_axi_araddr_T ), .A2(_04982_ ), .A3(_04983_ ), .A4(lsu_io_out_bits_rd_wdata_$_MUX__Y_15_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06125_ ) );
OAI21_X1 _26937_ ( .A(_05498_ ), .B1(_06124_ ), .B2(_06125_ ), .ZN(_06126_ ) );
AND3_X1 _26938_ ( .A1(_05496_ ), .A2(_03906_ ), .A3(_05495_ ), .ZN(_06127_ ) );
AOI21_X1 _26939_ ( .A(_06127_ ), .B1(_04833_ ), .B2(\io_master_awaddr [1] ), .ZN(_06128_ ) );
OAI211_X1 _26940_ ( .A(_05565_ ), .B(_06126_ ), .C1(_06128_ ), .C2(_04462_ ), .ZN(_06129_ ) );
NAND2_X1 _26941_ ( .A1(_03927_ ), .A2(\lsu.io_in_bits_rd_wdata [0] ), .ZN(_06130_ ) );
AND3_X1 _26942_ ( .A1(_06129_ ), .A2(_03925_ ), .A3(_06130_ ), .ZN(_06131_ ) );
NAND4_X1 _26943_ ( .A1(_03990_ ), .A2(\wbu.io_in_bits_rd_wdata [0] ), .A3(_03997_ ), .A4(_04010_ ), .ZN(_06132_ ) );
AOI211_X1 _26944_ ( .A(_03859_ ), .B(_06131_ ), .C1(_03931_ ), .C2(_06132_ ), .ZN(_06133_ ) );
OAI21_X1 _26945_ ( .A(_03850_ ), .B1(_06123_ ), .B2(_06133_ ), .ZN(_06134_ ) );
INV_X1 _26946_ ( .A(\wbu.rf_24 [0] ), .ZN(_06135_ ) );
NOR3_X1 _26947_ ( .A1(_04548_ ), .A2(_06135_ ), .A3(_04327_ ), .ZN(_06136_ ) );
AOI21_X1 _26948_ ( .A(_06136_ ), .B1(_04164_ ), .B2(\wbu.rf_21 [0] ), .ZN(_06137_ ) );
AND3_X1 _26949_ ( .A1(_04082_ ), .A2(\wbu.rf_7 [0] ), .A3(_04545_ ), .ZN(_06138_ ) );
AOI21_X1 _26950_ ( .A(_06138_ ), .B1(\wbu.rf_8 [0] ), .B2(_04089_ ), .ZN(_06139_ ) );
AOI22_X1 _26951_ ( .A1(\wbu._GEN_71 [0] ), .A2(_04059_ ), .B1(_04068_ ), .B2(\wbu.rf_4 [0] ), .ZN(_06140_ ) );
AOI22_X1 _26952_ ( .A1(\wbu.rf_22 [0] ), .A2(_04434_ ), .B1(_04305_ ), .B2(\wbu.rf_20 [0] ), .ZN(_06141_ ) );
AND4_X1 _26953_ ( .A1(_06137_ ), .A2(_06139_ ), .A3(_06140_ ), .A4(_06141_ ), .ZN(_06142_ ) );
NAND3_X1 _26954_ ( .A1(_04021_ ), .A2(\wbu.rf_31 [0] ), .A3(_04242_ ), .ZN(_06143_ ) );
NAND3_X1 _26955_ ( .A1(_04217_ ), .A2(\wbu.rf_25 [0] ), .A3(_04196_ ), .ZN(_06144_ ) );
NAND2_X1 _26956_ ( .A1(_06143_ ), .A2(_06144_ ), .ZN(_06145_ ) );
AOI221_X4 _26957_ ( .A(_06145_ ), .B1(\wbu.rf_30 [0] ), .B2(_05206_ ), .C1(\wbu.rf_29 [0] ), .C2(_04218_ ), .ZN(_06146_ ) );
AOI22_X1 _26958_ ( .A1(\wbu.rf_26 [0] ), .A2(_04203_ ), .B1(_04446_ ), .B2(\wbu.rf_28 [0] ), .ZN(_06147_ ) );
AOI22_X1 _26959_ ( .A1(\wbu.rf_27 [0] ), .A2(_04201_ ), .B1(_04100_ ), .B2(\wbu.rf_11 [0] ), .ZN(_06148_ ) );
NAND4_X1 _26960_ ( .A1(_06142_ ), .A2(_06146_ ), .A3(_06147_ ), .A4(_06148_ ), .ZN(_06149_ ) );
AOI22_X1 _26961_ ( .A1(\wbu.rf_23 [0] ), .A2(_05038_ ), .B1(_04139_ ), .B2(\wbu.rf_18 [0] ), .ZN(_06150_ ) );
AOI22_X1 _26962_ ( .A1(\wbu.rf_10 [0] ), .A2(_04845_ ), .B1(_04105_ ), .B2(\wbu.rf_12 [0] ), .ZN(_06151_ ) );
AOI22_X1 _26963_ ( .A1(\wbu.rf_13 [0] ), .A2(_04285_ ), .B1(_04292_ ), .B2(\wbu.rf_16 [0] ), .ZN(_06152_ ) );
AOI22_X1 _26964_ ( .A1(_04516_ ), .A2(\wbu.rf_14 [0] ), .B1(_04092_ ), .B2(\wbu.rf_9 [0] ), .ZN(_06153_ ) );
NAND4_X1 _26965_ ( .A1(_06150_ ), .A2(_06151_ ), .A3(_06152_ ), .A4(_06153_ ), .ZN(_06154_ ) );
AOI22_X1 _26966_ ( .A1(\wbu.rf_19 [0] ), .A2(_04301_ ), .B1(_04392_ ), .B2(\wbu.rf_3 [0] ), .ZN(_06155_ ) );
AOI22_X1 _26967_ ( .A1(\wbu.rf_5 [0] ), .A2(_04395_ ), .B1(_04578_ ), .B2(\wbu.rf_15 [0] ), .ZN(_06156_ ) );
AOI22_X1 _26968_ ( .A1(\wbu.rf_6 [0] ), .A2(_04271_ ), .B1(_04053_ ), .B2(\wbu.rf_2 [0] ), .ZN(_06157_ ) );
NAND3_X1 _26969_ ( .A1(_04134_ ), .A2(\wbu.rf_17 [0] ), .A3(_04212_ ), .ZN(_06158_ ) );
NAND4_X1 _26970_ ( .A1(_06155_ ), .A2(_06156_ ), .A3(_06157_ ), .A4(_06158_ ), .ZN(_06159_ ) );
NOR3_X1 _26971_ ( .A1(_06149_ ), .A2(_06154_ ), .A3(_06159_ ), .ZN(_06160_ ) );
OAI21_X1 _26972_ ( .A(_06134_ ), .B1(_04240_ ), .B2(_06160_ ), .ZN(\idu.io_out_bits_rs1_data [0] ) );
AND2_X1 _26973_ ( .A1(_06129_ ), .A2(_06130_ ), .ZN(_06161_ ) );
INV_X1 _26974_ ( .A(_06161_ ), .ZN(\lsu.io_out_bits_rd_wdata [0] ) );
NOR2_X1 _26975_ ( .A1(_03583_ ), .A2(_03857_ ), .ZN(_06162_ ) );
AND3_X1 _26976_ ( .A1(_05498_ ), .A2(\arbiter.io_lsu_arsize [1] ), .A3(_04649_ ), .ZN(_06163_ ) );
NOR3_X1 _26977_ ( .A1(_04461_ ), .A2(_03917_ ), .A3(_06163_ ), .ZN(_06164_ ) );
NOR2_X1 _26978_ ( .A1(\lsu.io_in_bits_ren ), .A2(\lsu.io_in_bits_rd_wdata [27] ), .ZN(_06165_ ) );
NOR2_X1 _26979_ ( .A1(_06164_ ), .A2(_06165_ ), .ZN(\lsu.io_out_bits_rd_wdata [27] ) );
NOR2_X1 _26980_ ( .A1(\lsu.io_out_bits_rd_wdata [27] ), .A2(_03931_ ), .ZN(_06166_ ) );
NAND4_X1 _26981_ ( .A1(_03991_ ), .A2(\wbu.io_in_bits_rd_wdata [27] ), .A3(_03998_ ), .A4(_04011_ ), .ZN(_06167_ ) );
AOI211_X1 _26982_ ( .A(_04459_ ), .B(_06166_ ), .C1(_03932_ ), .C2(_06167_ ), .ZN(_06168_ ) );
OAI21_X1 _26983_ ( .A(_03851_ ), .B1(_06162_ ), .B2(_06168_ ), .ZN(_06169_ ) );
NAND3_X1 _26984_ ( .A1(_04571_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04482_ ), .ZN(_06170_ ) );
NOR4_X1 _26985_ ( .A1(_04544_ ), .A2(_04534_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04545_ ), .ZN(_06171_ ) );
NOR3_X1 _26986_ ( .A1(_05325_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04549_ ), .ZN(_06172_ ) );
NOR2_X1 _26987_ ( .A1(_06172_ ), .A2(_04434_ ), .ZN(_06173_ ) );
AND3_X1 _26988_ ( .A1(_04162_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11101_ ), .ZN(_06174_ ) );
NAND4_X1 _26989_ ( .A1(_04155_ ), .A2(_04037_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_11101_ ), .ZN(_06175_ ) );
OR4_X1 _26990_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04123_ ), .A3(_04918_ ), .A4(_04016_ ), .ZN(_06176_ ) );
INV_X1 _26991_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_06177_ ) );
AOI22_X1 _26992_ ( .A1(_04059_ ), .A2(_06177_ ), .B1(_04411_ ), .B2(_04051_ ), .ZN(_06178_ ) );
AND4_X1 _26993_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04116_ ), .A3(_04149_ ), .A4(_11100_ ), .ZN(_06179_ ) );
OAI21_X1 _26994_ ( .A(_06176_ ), .B1(_06178_ ), .B2(_06179_ ), .ZN(_06180_ ) );
OAI21_X1 _26995_ ( .A(_06175_ ), .B1(_06180_ ), .B2(_04068_ ), .ZN(_06181_ ) );
AOI21_X1 _26996_ ( .A(_06174_ ), .B1(_06181_ ), .B2(_04496_ ), .ZN(_06182_ ) );
AOI211_X1 _26997_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_05653_ ), .C1(\idu.io_in_bits_inst [19] ), .C2(_04003_ ), .ZN(_06183_ ) );
NOR2_X1 _26998_ ( .A1(_06182_ ), .A2(_06183_ ), .ZN(_06184_ ) );
OR2_X1 _26999_ ( .A1(_04085_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06185_ ) );
OR3_X1 _27000_ ( .A1(_04187_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04018_ ), .ZN(_06186_ ) );
NAND3_X1 _27001_ ( .A1(_06184_ ), .A2(_06185_ ), .A3(_06186_ ), .ZN(_06187_ ) );
NOR3_X1 _27002_ ( .A1(_05011_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04019_ ), .ZN(_06188_ ) );
INV_X1 _27003_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06189_ ) );
AND4_X1 _27004_ ( .A1(_06189_ ), .A2(_04509_ ), .A3(_04169_ ), .A4(_04043_ ), .ZN(_06190_ ) );
NOR3_X1 _27005_ ( .A1(_06187_ ), .A2(_06188_ ), .A3(_06190_ ), .ZN(_06191_ ) );
INV_X1 _27006_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06192_ ) );
NAND4_X1 _27007_ ( .A1(_04332_ ), .A2(_04147_ ), .A3(_06192_ ), .A4(_04437_ ), .ZN(_06193_ ) );
OR3_X1 _27008_ ( .A1(_05201_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04173_ ), .ZN(_06194_ ) );
NAND3_X1 _27009_ ( .A1(_06191_ ), .A2(_06193_ ), .A3(_06194_ ), .ZN(_06195_ ) );
INV_X1 _27010_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06196_ ) );
AND4_X1 _27011_ ( .A1(_06196_ ), .A2(_04936_ ), .A3(_04522_ ), .A4(_04437_ ), .ZN(_06197_ ) );
INV_X1 _27012_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06198_ ) );
AND4_X1 _27013_ ( .A1(_06198_ ), .A2(_04170_ ), .A3(_04522_ ), .A4(_04295_ ), .ZN(_06199_ ) );
NOR3_X1 _27014_ ( .A1(_06195_ ), .A2(_06197_ ), .A3(_06199_ ), .ZN(_06200_ ) );
OR3_X1 _27015_ ( .A1(_04943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04174_ ), .ZN(_06201_ ) );
OR3_X1 _27016_ ( .A1(_04029_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04947_ ), .ZN(_06202_ ) );
NAND3_X1 _27017_ ( .A1(_06200_ ), .A2(_06201_ ), .A3(_06202_ ), .ZN(_06203_ ) );
NOR3_X1 _27018_ ( .A1(_04485_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04184_ ), .ZN(_06204_ ) );
OAI21_X1 _27019_ ( .A(_04303_ ), .B1(_04711_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06205_ ) );
NOR3_X1 _27020_ ( .A1(_06203_ ), .A2(_06204_ ), .A3(_06205_ ), .ZN(_06206_ ) );
AND3_X1 _27021_ ( .A1(_04062_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04842_ ), .ZN(_06207_ ) );
OAI221_X1 _27022_ ( .A(_06173_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04428_ ), .C1(_06206_ ), .C2(_06207_ ), .ZN(_06208_ ) );
NAND4_X1 _27023_ ( .A1(_04536_ ), .A2(_04615_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04210_ ), .ZN(_06209_ ) );
AOI21_X1 _27024_ ( .A(_06171_ ), .B1(_06208_ ), .B2(_06209_ ), .ZN(_06210_ ) );
OR3_X1 _27025_ ( .A1(_04548_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04819_ ), .ZN(_06211_ ) );
INV_X1 _27026_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06212_ ) );
NAND4_X1 _27027_ ( .A1(_04552_ ), .A2(_04553_ ), .A3(_06212_ ), .A4(_04455_ ), .ZN(_06213_ ) );
NAND3_X1 _27028_ ( .A1(_06210_ ), .A2(_06211_ ), .A3(_06213_ ), .ZN(_06214_ ) );
INV_X1 _27029_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06215_ ) );
AND4_X1 _27030_ ( .A1(_06215_ ), .A2(_04333_ ), .A3(_04728_ ), .A4(_04624_ ), .ZN(_06216_ ) );
NOR4_X1 _27031_ ( .A1(_05554_ ), .A2(_04544_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04550_ ), .ZN(_06217_ ) );
NOR3_X1 _27032_ ( .A1(_06214_ ), .A2(_06216_ ), .A3(_06217_ ), .ZN(_06218_ ) );
OR3_X1 _27033_ ( .A1(_05202_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04820_ ), .ZN(_06219_ ) );
INV_X1 _27034_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06220_ ) );
NAND3_X1 _27035_ ( .A1(_04562_ ), .A2(_06220_ ), .A3(_04224_ ), .ZN(_06221_ ) );
NAND3_X1 _27036_ ( .A1(_06218_ ), .A2(_06219_ ), .A3(_06221_ ), .ZN(_06222_ ) );
AOI211_X1 _27037_ ( .A(_04566_ ), .B(_04567_ ), .C1(_04568_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06223_ ) );
OAI211_X1 _27038_ ( .A(_04481_ ), .B(_06170_ ), .C1(_06222_ ), .C2(_06223_ ), .ZN(_06224_ ) );
NAND2_X1 _27039_ ( .A1(_06169_ ), .A2(_06224_ ), .ZN(\idu.io_out_bits_rs1_data [27] ) );
AOI21_X1 _27040_ ( .A(_04738_ ), .B1(_03628_ ), .B2(_03629_ ), .ZN(_06225_ ) );
NAND3_X1 _27041_ ( .A1(_05348_ ), .A2(\arbiter._io_axi_araddr_T ), .A3(\arbiter.io_lsu_arsize [1] ), .ZN(_06226_ ) );
OAI21_X1 _27042_ ( .A(_04642_ ), .B1(_03899_ ), .B2(_06226_ ), .ZN(_06227_ ) );
OAI21_X1 _27043_ ( .A(\lsu.io_in_bits_ren ), .B1(_06227_ ), .B2(_03917_ ), .ZN(_06228_ ) );
NAND2_X1 _27044_ ( .A1(_04351_ ), .A2(\lsu.io_in_bits_rd_wdata [26] ), .ZN(_06229_ ) );
NAND2_X1 _27045_ ( .A1(_06228_ ), .A2(_06229_ ), .ZN(\lsu.io_out_bits_rd_wdata [26] ) );
NAND2_X1 _27046_ ( .A1(\lsu.io_out_bits_rd_wdata [26] ), .A2(_04353_ ), .ZN(_06230_ ) );
OAI211_X1 _27047_ ( .A(\wbu.io_in_bits_rd_wdata [26] ), .B(_04656_ ), .C1(_04657_ ), .C2(_04658_ ), .ZN(_06231_ ) );
AOI21_X1 _27048_ ( .A(_04356_ ), .B1(_06230_ ), .B2(_06231_ ), .ZN(_06232_ ) );
OAI21_X1 _27049_ ( .A(_03851_ ), .B1(_06225_ ), .B2(_06232_ ), .ZN(_06233_ ) );
NAND3_X1 _27050_ ( .A1(_04571_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04243_ ), .ZN(_06234_ ) );
INV_X1 _27051_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_06235_ ) );
NAND3_X1 _27052_ ( .A1(_04134_ ), .A2(_06235_ ), .A3(_11100_ ), .ZN(_06236_ ) );
OAI21_X1 _27053_ ( .A(_06236_ ), .B1(_05293_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06237_ ) );
NOR2_X1 _27054_ ( .A1(_04497_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06238_ ) );
INV_X1 _27055_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06239_ ) );
AND4_X1 _27056_ ( .A1(_06239_ ), .A2(_04144_ ), .A3(_04149_ ), .A4(_04080_ ), .ZN(_06240_ ) );
NOR3_X1 _27057_ ( .A1(_06237_ ), .A2(_06238_ ), .A3(_06240_ ), .ZN(_06241_ ) );
INV_X1 _27058_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06242_ ) );
NAND4_X1 _27059_ ( .A1(_04108_ ), .A2(_04858_ ), .A3(_06242_ ), .A4(_11101_ ), .ZN(_06243_ ) );
OR3_X1 _27060_ ( .A1(_05653_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04017_ ), .ZN(_06244_ ) );
NAND3_X1 _27061_ ( .A1(_06241_ ), .A2(_06243_ ), .A3(_06244_ ), .ZN(_06245_ ) );
INV_X1 _27062_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06246_ ) );
AND4_X1 _27063_ ( .A1(_06246_ ), .A2(_04145_ ), .A3(_04858_ ), .A4(_04282_ ), .ZN(_06247_ ) );
NOR3_X1 _27064_ ( .A1(_04187_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04128_ ), .ZN(_06248_ ) );
NOR3_X1 _27065_ ( .A1(_06245_ ), .A2(_06247_ ), .A3(_06248_ ), .ZN(_06249_ ) );
INV_X1 _27066_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06250_ ) );
NAND3_X1 _27067_ ( .A1(_04504_ ), .A2(_06250_ ), .A3(_04385_ ), .ZN(_06251_ ) );
INV_X1 _27068_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06252_ ) );
NAND4_X1 _27069_ ( .A1(_04509_ ), .A2(_04169_ ), .A3(_06252_ ), .A4(_04113_ ), .ZN(_06253_ ) );
NAND3_X1 _27070_ ( .A1(_06249_ ), .A2(_06251_ ), .A3(_06253_ ), .ZN(_06254_ ) );
NOR4_X1 _27071_ ( .A1(_05554_ ), .A2(_04125_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04163_ ), .ZN(_06255_ ) );
NOR3_X1 _27072_ ( .A1(_05201_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04129_ ), .ZN(_06256_ ) );
NOR3_X1 _27073_ ( .A1(_06254_ ), .A2(_06255_ ), .A3(_06256_ ), .ZN(_06257_ ) );
INV_X1 _27074_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06258_ ) );
NAND4_X1 _27075_ ( .A1(_04936_ ), .A2(_04522_ ), .A3(_06258_ ), .A4(_04295_ ), .ZN(_06259_ ) );
INV_X1 _27076_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06260_ ) );
NAND4_X1 _27077_ ( .A1(_04170_ ), .A2(_04522_ ), .A3(_06260_ ), .A4(_04295_ ), .ZN(_06261_ ) );
NAND3_X1 _27078_ ( .A1(_06257_ ), .A2(_06259_ ), .A3(_06261_ ), .ZN(_06262_ ) );
NOR3_X1 _27079_ ( .A1(_04943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04159_ ), .ZN(_06263_ ) );
NOR3_X1 _27080_ ( .A1(_04029_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04947_ ), .ZN(_06264_ ) );
NOR3_X1 _27081_ ( .A1(_06262_ ), .A2(_06263_ ), .A3(_06264_ ), .ZN(_06265_ ) );
OR3_X1 _27082_ ( .A1(_04485_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04437_ ), .ZN(_06266_ ) );
INV_X1 _27083_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06267_ ) );
NAND4_X1 _27084_ ( .A1(_04297_ ), .A2(_04525_ ), .A3(_06267_ ), .A4(_04208_ ), .ZN(_06268_ ) );
NAND3_X1 _27085_ ( .A1(_06265_ ), .A2(_06266_ ), .A3(_06268_ ), .ZN(_06269_ ) );
NOR4_X1 _27086_ ( .A1(_04178_ ), .A2(_04947_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04190_ ), .ZN(_06270_ ) );
NOR3_X1 _27087_ ( .A1(_04029_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04317_ ), .ZN(_06271_ ) );
NOR3_X1 _27088_ ( .A1(_06269_ ), .A2(_06270_ ), .A3(_06271_ ), .ZN(_06272_ ) );
INV_X1 _27089_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06273_ ) );
NAND4_X1 _27090_ ( .A1(_04217_ ), .A2(_04168_ ), .A3(_06273_ ), .A4(_04842_ ), .ZN(_06274_ ) );
INV_X1 _27091_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06275_ ) );
NAND4_X1 _27092_ ( .A1(_04168_ ), .A2(_04528_ ), .A3(_06275_ ), .A4(_04842_ ), .ZN(_06276_ ) );
AND3_X1 _27093_ ( .A1(_06272_ ), .A2(_06274_ ), .A3(_06276_ ), .ZN(_06277_ ) );
OR4_X1 _27094_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04179_ ), .A3(_04182_ ), .A4(_04184_ ), .ZN(_06278_ ) );
OR3_X1 _27095_ ( .A1(_04188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04549_ ), .ZN(_06279_ ) );
NAND3_X1 _27096_ ( .A1(_06277_ ), .A2(_06278_ ), .A3(_06279_ ), .ZN(_06280_ ) );
INV_X1 _27097_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06281_ ) );
AND4_X1 _27098_ ( .A1(_04194_ ), .A2(_04197_ ), .A3(_06281_ ), .A4(_04199_ ), .ZN(_06282_ ) );
OAI21_X1 _27099_ ( .A(_04202_ ), .B1(_04204_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06283_ ) );
NOR3_X1 _27100_ ( .A1(_06280_ ), .A2(_06282_ ), .A3(_06283_ ), .ZN(_06284_ ) );
AND3_X1 _27101_ ( .A1(_04207_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04624_ ), .ZN(_06285_ ) );
OR2_X1 _27102_ ( .A1(_06284_ ), .A2(_06285_ ), .ZN(_06286_ ) );
OR3_X1 _27103_ ( .A1(_05202_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04820_ ), .ZN(_06287_ ) );
OR3_X1 _27104_ ( .A1(_04636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04820_ ), .ZN(_06288_ ) );
NAND3_X1 _27105_ ( .A1(_06286_ ), .A2(_06287_ ), .A3(_06288_ ), .ZN(_06289_ ) );
AOI211_X1 _27106_ ( .A(_04566_ ), .B(_04567_ ), .C1(_04568_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06290_ ) );
OAI211_X1 _27107_ ( .A(_04247_ ), .B(_06234_ ), .C1(_06289_ ), .C2(_06290_ ), .ZN(_06291_ ) );
NAND2_X1 _27108_ ( .A1(_06233_ ), .A2(_06291_ ), .ZN(\idu.io_out_bits_rs1_data [26] ) );
AOI21_X1 _27109_ ( .A(_04738_ ), .B1(_03676_ ), .B2(_03677_ ), .ZN(_06292_ ) );
AND3_X1 _27110_ ( .A1(_05498_ ), .A2(\arbiter.io_lsu_arsize [1] ), .A3(_04758_ ), .ZN(_06293_ ) );
OR2_X1 _27111_ ( .A1(_03898_ ), .A2(_06293_ ), .ZN(_06294_ ) );
OAI21_X1 _27112_ ( .A(\lsu.io_in_bits_ren ), .B1(_06294_ ), .B2(_03917_ ), .ZN(_06295_ ) );
NAND2_X1 _27113_ ( .A1(_04351_ ), .A2(\lsu.io_in_bits_rd_wdata [25] ), .ZN(_06296_ ) );
NAND2_X1 _27114_ ( .A1(_06295_ ), .A2(_06296_ ), .ZN(\lsu.io_out_bits_rd_wdata [25] ) );
NAND2_X1 _27115_ ( .A1(\lsu.io_out_bits_rd_wdata [25] ), .A2(_04353_ ), .ZN(_06297_ ) );
OAI211_X1 _27116_ ( .A(\wbu.io_in_bits_rd_wdata [25] ), .B(_04656_ ), .C1(_04657_ ), .C2(_04658_ ), .ZN(_06298_ ) );
AOI21_X1 _27117_ ( .A(_04356_ ), .B1(_06297_ ), .B2(_06298_ ), .ZN(_06299_ ) );
OAI21_X1 _27118_ ( .A(_03851_ ), .B1(_06292_ ), .B2(_06299_ ), .ZN(_06300_ ) );
NAND3_X1 _27119_ ( .A1(_04571_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04243_ ), .ZN(_06301_ ) );
NOR3_X1 _27120_ ( .A1(_04485_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04190_ ), .ZN(_06302_ ) );
NAND3_X1 _27121_ ( .A1(_04606_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04936_ ), .ZN(_06303_ ) );
NAND3_X1 _27122_ ( .A1(_04504_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04109_ ), .ZN(_06304_ ) );
INV_X1 _27123_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06305_ ) );
AND3_X1 _27124_ ( .A1(_04078_ ), .A2(_06305_ ), .A3(_04282_ ), .ZN(_06306_ ) );
INV_X1 _27125_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06307_ ) );
NAND3_X1 _27126_ ( .A1(_04051_ ), .A2(_06307_ ), .A3(_11100_ ), .ZN(_06308_ ) );
OAI21_X1 _27127_ ( .A(_06308_ ), .B1(_04493_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_06309_ ) );
NOR2_X1 _27128_ ( .A1(_04497_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06310_ ) );
INV_X1 _27129_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06311_ ) );
AND4_X1 _27130_ ( .A1(_06311_ ), .A2(_04144_ ), .A3(_04148_ ), .A4(_04040_ ), .ZN(_06312_ ) );
NOR3_X1 _27131_ ( .A1(_06309_ ), .A2(_06310_ ), .A3(_06312_ ), .ZN(_06313_ ) );
NAND2_X1 _27132_ ( .A1(_06313_ ), .A2(_04496_ ), .ZN(_06314_ ) );
NAND4_X1 _27133_ ( .A1(_04108_ ), .A2(_04155_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04042_ ), .ZN(_06315_ ) );
AOI21_X1 _27134_ ( .A(_06306_ ), .B1(_06314_ ), .B2(_06315_ ), .ZN(_06316_ ) );
OAI21_X1 _27135_ ( .A(_06316_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04085_ ), .ZN(_06317_ ) );
OAI21_X1 _27136_ ( .A(_04093_ ), .B1(_04090_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06318_ ) );
OAI21_X1 _27137_ ( .A(_06304_ ), .B1(_06317_ ), .B2(_06318_ ), .ZN(_06319_ ) );
INV_X1 _27138_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06320_ ) );
NAND4_X1 _27139_ ( .A1(_04332_ ), .A2(_04119_ ), .A3(_06320_ ), .A4(_04114_ ), .ZN(_06321_ ) );
INV_X1 _27140_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06322_ ) );
NAND4_X1 _27141_ ( .A1(_04332_ ), .A2(_04146_ ), .A3(_06322_ ), .A4(_04114_ ), .ZN(_06323_ ) );
NAND3_X1 _27142_ ( .A1(_06319_ ), .A2(_06321_ ), .A3(_06323_ ), .ZN(_06324_ ) );
OAI21_X1 _27143_ ( .A(_04704_ ), .B1(_04414_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06325_ ) );
OAI21_X1 _27144_ ( .A(_06303_ ), .B1(_06324_ ), .B2(_06325_ ), .ZN(_06326_ ) );
INV_X1 _27145_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06327_ ) );
NAND4_X1 _27146_ ( .A1(_04297_ ), .A2(_04445_ ), .A3(_06327_ ), .A4(_04183_ ), .ZN(_06328_ ) );
INV_X1 _27147_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06329_ ) );
NAND3_X1 _27148_ ( .A1(_04606_ ), .A2(_06329_ ), .A3(_04241_ ), .ZN(_06330_ ) );
NAND4_X1 _27149_ ( .A1(_06326_ ), .A2(_05880_ ), .A3(_06328_ ), .A4(_06330_ ), .ZN(_06331_ ) );
NAND4_X1 _27150_ ( .A1(_04525_ ), .A2(_04158_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04310_ ), .ZN(_06332_ ) );
AOI21_X1 _27151_ ( .A(_06302_ ), .B1(_06331_ ), .B2(_06332_ ), .ZN(_06333_ ) );
INV_X1 _27152_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06334_ ) );
NAND4_X1 _27153_ ( .A1(_04528_ ), .A2(_04529_ ), .A3(_06334_ ), .A4(_04209_ ), .ZN(_06335_ ) );
INV_X1 _27154_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06336_ ) );
NAND4_X1 _27155_ ( .A1(_04241_ ), .A2(_04529_ ), .A3(_06336_ ), .A4(_04175_ ), .ZN(_06337_ ) );
AND3_X1 _27156_ ( .A1(_06333_ ), .A2(_06335_ ), .A3(_06337_ ), .ZN(_06338_ ) );
OR3_X1 _27157_ ( .A1(_04030_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04182_ ), .ZN(_06339_ ) );
OR3_X1 _27158_ ( .A1(_05325_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04191_ ), .ZN(_06340_ ) );
NAND3_X1 _27159_ ( .A1(_06338_ ), .A2(_06339_ ), .A3(_06340_ ), .ZN(_06341_ ) );
INV_X1 _27160_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06342_ ) );
AND4_X1 _27161_ ( .A1(_06342_ ), .A2(_04542_ ), .A3(_04528_ ), .A4(_04623_ ), .ZN(_06343_ ) );
NOR4_X1 _27162_ ( .A1(_04179_ ), .A2(_04534_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04545_ ), .ZN(_06344_ ) );
NOR3_X1 _27163_ ( .A1(_06341_ ), .A2(_06343_ ), .A3(_06344_ ), .ZN(_06345_ ) );
OR3_X1 _27164_ ( .A1(_04548_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04819_ ), .ZN(_06346_ ) );
INV_X1 _27165_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06347_ ) );
NAND4_X1 _27166_ ( .A1(_04552_ ), .A2(_04553_ ), .A3(_06347_ ), .A4(_04455_ ), .ZN(_06348_ ) );
NAND3_X1 _27167_ ( .A1(_06345_ ), .A2(_06346_ ), .A3(_06348_ ), .ZN(_06349_ ) );
NOR3_X1 _27168_ ( .A1(_04326_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04637_ ), .ZN(_06350_ ) );
INV_X1 _27169_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06351_ ) );
AND4_X1 _27170_ ( .A1(_06351_ ), .A2(_04333_ ), .A3(_04242_ ), .A4(_04624_ ), .ZN(_06352_ ) );
NOR3_X1 _27171_ ( .A1(_06349_ ), .A2(_06350_ ), .A3(_06352_ ), .ZN(_06353_ ) );
OR3_X1 _27172_ ( .A1(_05202_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04820_ ), .ZN(_06354_ ) );
INV_X1 _27173_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06355_ ) );
NAND3_X1 _27174_ ( .A1(_04562_ ), .A2(_06355_ ), .A3(_04224_ ), .ZN(_06356_ ) );
NAND3_X1 _27175_ ( .A1(_06353_ ), .A2(_06354_ ), .A3(_06356_ ), .ZN(_06357_ ) );
AOI211_X1 _27176_ ( .A(_04566_ ), .B(_04567_ ), .C1(_04568_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06358_ ) );
OAI211_X1 _27177_ ( .A(_04247_ ), .B(_06301_ ), .C1(_06357_ ), .C2(_06358_ ), .ZN(_06359_ ) );
NAND2_X1 _27178_ ( .A1(_06300_ ), .A2(_06359_ ), .ZN(\idu.io_out_bits_rs1_data [25] ) );
AOI21_X1 _27179_ ( .A(_03857_ ), .B1(_03722_ ), .B2(_03723_ ), .ZN(_06360_ ) );
NOR3_X1 _27180_ ( .A1(_03899_ ), .A2(_03900_ ), .A3(_04829_ ), .ZN(_06361_ ) );
OR2_X1 _27181_ ( .A1(_03898_ ), .A2(_06361_ ), .ZN(_06362_ ) );
OAI21_X1 _27182_ ( .A(\lsu.io_in_bits_ren ), .B1(_06362_ ), .B2(_03917_ ), .ZN(_06363_ ) );
NAND2_X1 _27183_ ( .A1(_04351_ ), .A2(\lsu.io_in_bits_rd_wdata [24] ), .ZN(_06364_ ) );
AND3_X1 _27184_ ( .A1(_06363_ ), .A2(_03925_ ), .A3(_06364_ ), .ZN(_06365_ ) );
NAND4_X1 _27185_ ( .A1(_03991_ ), .A2(\wbu.io_in_bits_rd_wdata [24] ), .A3(_03998_ ), .A4(_04011_ ), .ZN(_06366_ ) );
AOI211_X1 _27186_ ( .A(_03859_ ), .B(_06365_ ), .C1(_03932_ ), .C2(_06366_ ), .ZN(_06367_ ) );
OAI21_X1 _27187_ ( .A(_03850_ ), .B1(_06360_ ), .B2(_06367_ ), .ZN(_06368_ ) );
NAND3_X1 _27188_ ( .A1(_04571_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04243_ ), .ZN(_06369_ ) );
OR4_X1 _27189_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04316_ ), .A3(_04317_ ), .A4(_04318_ ), .ZN(_06370_ ) );
INV_X1 _27190_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_06371_ ) );
NAND3_X1 _27191_ ( .A1(_04134_ ), .A2(_06371_ ), .A3(_04040_ ), .ZN(_06372_ ) );
OAI21_X1 _27192_ ( .A(_06372_ ), .B1(_05293_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06373_ ) );
INV_X1 _27193_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06374_ ) );
AOI21_X1 _27194_ ( .A(_06373_ ), .B1(_06374_ ), .B2(_04392_ ), .ZN(_06375_ ) );
OR2_X1 _27195_ ( .A1(_04497_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06376_ ) );
INV_X1 _27196_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06377_ ) );
NAND4_X1 _27197_ ( .A1(_04384_ ), .A2(_04858_ ), .A3(_06377_ ), .A4(_04411_ ), .ZN(_06378_ ) );
AND3_X1 _27198_ ( .A1(_06375_ ), .A2(_06376_ ), .A3(_06378_ ), .ZN(_06379_ ) );
OR3_X1 _27199_ ( .A1(_05653_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04017_ ), .ZN(_06380_ ) );
OR4_X1 _27200_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04124_ ), .A3(_04180_ ), .A4(_04127_ ), .ZN(_06381_ ) );
NAND3_X1 _27201_ ( .A1(_06379_ ), .A2(_06380_ ), .A3(_06381_ ), .ZN(_06382_ ) );
INV_X1 _27202_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06383_ ) );
AND3_X1 _27203_ ( .A1(_04504_ ), .A2(_06383_ ), .A3(_04037_ ), .ZN(_06384_ ) );
INV_X1 _27204_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06385_ ) );
AND3_X1 _27205_ ( .A1(_04504_ ), .A2(_06385_ ), .A3(_04108_ ), .ZN(_06386_ ) );
NOR3_X1 _27206_ ( .A1(_06382_ ), .A2(_06384_ ), .A3(_06386_ ), .ZN(_06387_ ) );
INV_X1 _27207_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06388_ ) );
NAND4_X1 _27208_ ( .A1(_04509_ ), .A2(_04169_ ), .A3(_06388_ ), .A4(_04043_ ), .ZN(_06389_ ) );
OR4_X1 _27209_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_05437_ ), .A3(_04125_ ), .A4(_04128_ ), .ZN(_06390_ ) );
NAND3_X1 _27210_ ( .A1(_06387_ ), .A2(_06389_ ), .A3(_06390_ ), .ZN(_06391_ ) );
INV_X1 _27211_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06392_ ) );
AND4_X1 _27212_ ( .A1(_06392_ ), .A2(_04036_ ), .A3(_04038_ ), .A4(_04043_ ), .ZN(_06393_ ) );
INV_X1 _27213_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06394_ ) );
AND4_X1 _27214_ ( .A1(_06394_ ), .A2(_04109_ ), .A3(_04036_ ), .A4(_04043_ ), .ZN(_06395_ ) );
NOR3_X1 _27215_ ( .A1(_06391_ ), .A2(_06393_ ), .A3(_06395_ ), .ZN(_06396_ ) );
OR2_X1 _27216_ ( .A1(_05019_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06397_ ) );
OR3_X1 _27217_ ( .A1(_04943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04019_ ), .ZN(_06398_ ) );
NAND3_X1 _27218_ ( .A1(_06396_ ), .A2(_06397_ ), .A3(_06398_ ), .ZN(_06399_ ) );
INV_X1 _27219_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06400_ ) );
AND4_X1 _27220_ ( .A1(_06400_ ), .A2(_04253_ ), .A3(_04157_ ), .A4(_04254_ ), .ZN(_06401_ ) );
INV_X1 _27221_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06402_ ) );
AND4_X1 _27222_ ( .A1(_06402_ ), .A2(_04936_ ), .A3(_04253_ ), .A4(_04254_ ), .ZN(_06403_ ) );
NOR3_X1 _27223_ ( .A1(_06399_ ), .A2(_06401_ ), .A3(_06403_ ), .ZN(_06404_ ) );
OR2_X1 _27224_ ( .A1(_04711_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06405_ ) );
OR4_X1 _27225_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04126_ ), .A3(_04947_ ), .A4(_04437_ ), .ZN(_06406_ ) );
NAND3_X1 _27226_ ( .A1(_06404_ ), .A2(_06405_ ), .A3(_06406_ ), .ZN(_06407_ ) );
INV_X1 _27227_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06408_ ) );
AND4_X1 _27228_ ( .A1(_06408_ ), .A2(_04167_ ), .A3(_04158_ ), .A4(_04208_ ), .ZN(_06409_ ) );
INV_X1 _27229_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06410_ ) );
AND4_X1 _27230_ ( .A1(_06410_ ), .A2(_04216_ ), .A3(_04167_ ), .A4(_04208_ ), .ZN(_06411_ ) );
NOR4_X1 _27231_ ( .A1(_06407_ ), .A2(_04434_ ), .A3(_06409_ ), .A4(_06411_ ), .ZN(_06412_ ) );
AND4_X1 _27232_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04168_ ), .A3(_04528_ ), .A4(_04209_ ), .ZN(_06413_ ) );
OAI21_X1 _27233_ ( .A(_06370_ ), .B1(_06412_ ), .B2(_06413_ ), .ZN(_06414_ ) );
INV_X1 _27234_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06415_ ) );
AND4_X1 _27235_ ( .A1(_06415_ ), .A2(_04332_ ), .A3(_04451_ ), .A4(_04623_ ), .ZN(_06416_ ) );
INV_X1 _27236_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06417_ ) );
AND4_X1 _27237_ ( .A1(_04000_ ), .A2(_04196_ ), .A3(_06417_ ), .A4(_10756_ ), .ZN(_06418_ ) );
NOR3_X1 _27238_ ( .A1(_06414_ ), .A2(_06416_ ), .A3(_06418_ ), .ZN(_06419_ ) );
INV_X1 _27239_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06420_ ) );
NAND4_X1 _27240_ ( .A1(_04620_ ), .A2(_04728_ ), .A3(_06420_ ), .A4(_04211_ ), .ZN(_06421_ ) );
OR4_X1 _27241_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_05554_ ), .A3(_04179_ ), .A4(_04545_ ), .ZN(_06422_ ) );
NAND3_X1 _27242_ ( .A1(_06419_ ), .A2(_06421_ ), .A3(_06422_ ), .ZN(_06423_ ) );
NOR3_X1 _27243_ ( .A1(_05202_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04637_ ), .ZN(_06424_ ) );
NOR3_X1 _27244_ ( .A1(_04636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04637_ ), .ZN(_06425_ ) );
OR3_X1 _27245_ ( .A1(_06423_ ), .A2(_06424_ ), .A3(_06425_ ), .ZN(_06426_ ) );
AOI211_X1 _27246_ ( .A(_04566_ ), .B(_04567_ ), .C1(_04568_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06427_ ) );
OAI211_X1 _27247_ ( .A(_04247_ ), .B(_06369_ ), .C1(_06426_ ), .C2(_06427_ ), .ZN(_06428_ ) );
NAND2_X1 _27248_ ( .A1(_06368_ ), .A2(_06428_ ), .ZN(\idu.io_out_bits_rs1_data [24] ) );
NAND2_X1 _27249_ ( .A1(_06363_ ), .A2(_06364_ ), .ZN(\lsu.io_out_bits_rd_wdata [24] ) );
NAND2_X1 _27250_ ( .A1(\exu.io_out_bits_rd_wdata [23] ), .A2(_04228_ ), .ZN(_06429_ ) );
OAI22_X1 _27251_ ( .A1(_03903_ ), .A2(_04370_ ), .B1(_03909_ ), .B2(_03892_ ), .ZN(_06430_ ) );
AOI22_X1 _27252_ ( .A1(_03897_ ), .A2(\lsu.io_in_bits_lh ), .B1(_06430_ ), .B2(\arbiter.io_lsu_arsize [1] ), .ZN(_06431_ ) );
AOI21_X1 _27253_ ( .A(_03927_ ), .B1(_04358_ ), .B2(_06431_ ), .ZN(_06432_ ) );
AND2_X1 _27254_ ( .A1(_03926_ ), .A2(\lsu.io_in_bits_rd_wdata [23] ), .ZN(_06433_ ) );
OR3_X1 _27255_ ( .A1(_06432_ ), .A2(_03930_ ), .A3(_06433_ ), .ZN(_06434_ ) );
NAND4_X1 _27256_ ( .A1(_03990_ ), .A2(\wbu.io_in_bits_rd_wdata [23] ), .A3(_03997_ ), .A4(_04010_ ), .ZN(_06435_ ) );
AOI21_X1 _27257_ ( .A(_03859_ ), .B1(_03931_ ), .B2(_06435_ ), .ZN(_06436_ ) );
NAND2_X1 _27258_ ( .A1(_06434_ ), .A2(_06436_ ), .ZN(_06437_ ) );
AOI21_X1 _27259_ ( .A(\idu.rs_reg ), .B1(_06429_ ), .B2(_06437_ ), .ZN(_06438_ ) );
NAND3_X1 _27260_ ( .A1(_04062_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04159_ ), .ZN(_06439_ ) );
NAND4_X1 _27261_ ( .A1(_04118_ ), .A2(_04110_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04598_ ), .ZN(_06440_ ) );
NAND4_X1 _27262_ ( .A1(_04073_ ), .A2(_04074_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04039_ ), .ZN(_06441_ ) );
INV_X1 _27263_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06442_ ) );
NAND4_X1 _27264_ ( .A1(_04046_ ), .A2(_04050_ ), .A3(_06442_ ), .A4(_11097_ ), .ZN(_06443_ ) );
OAI21_X1 _27265_ ( .A(_06443_ ), .B1(_04493_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_06444_ ) );
INV_X1 _27266_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06445_ ) );
AOI21_X1 _27267_ ( .A(_06444_ ), .B1(_06445_ ), .B2(_04392_ ), .ZN(_06446_ ) );
OR2_X1 _27268_ ( .A1(_04069_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06447_ ) );
NAND2_X1 _27269_ ( .A1(_06446_ ), .A2(_06447_ ), .ZN(_06448_ ) );
OAI21_X1 _27270_ ( .A(_06441_ ), .B1(_06448_ ), .B2(_04395_ ), .ZN(_06449_ ) );
INV_X1 _27271_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06450_ ) );
NAND3_X1 _27272_ ( .A1(_04077_ ), .A2(_06450_ ), .A3(_04399_ ), .ZN(_06451_ ) );
OR4_X1 _27273_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04123_ ), .A3(_04180_ ), .A4(_10766_ ), .ZN(_06452_ ) );
AND3_X1 _27274_ ( .A1(_06449_ ), .A2(_06451_ ), .A3(_06452_ ), .ZN(_06453_ ) );
OR3_X1 _27275_ ( .A1(_04186_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04016_ ), .ZN(_06454_ ) );
OR3_X1 _27276_ ( .A1(_05011_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03992_ ), .ZN(_06455_ ) );
NAND3_X1 _27277_ ( .A1(_06453_ ), .A2(_06454_ ), .A3(_06455_ ), .ZN(_06456_ ) );
NOR3_X1 _27278_ ( .A1(_04095_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04127_ ), .ZN(_06457_ ) );
NOR4_X1 _27279_ ( .A1(_05437_ ), .A2(_04124_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04016_ ), .ZN(_06458_ ) );
NOR3_X1 _27280_ ( .A1(_06456_ ), .A2(_06457_ ), .A3(_06458_ ), .ZN(_06459_ ) );
INV_X1 _27281_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06460_ ) );
NAND4_X1 _27282_ ( .A1(_04110_ ), .A2(_04037_ ), .A3(_06460_ ), .A4(_11101_ ), .ZN(_06461_ ) );
INV_X1 _27283_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06462_ ) );
NAND4_X1 _27284_ ( .A1(_04108_ ), .A2(_04032_ ), .A3(_06462_ ), .A4(_04282_ ), .ZN(_06463_ ) );
NAND3_X1 _27285_ ( .A1(_06459_ ), .A2(_06461_ ), .A3(_06463_ ), .ZN(_06464_ ) );
OAI21_X1 _27286_ ( .A(_06440_ ), .B1(_06464_ ), .B2(_04516_ ), .ZN(_06465_ ) );
INV_X1 _27287_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06466_ ) );
NAND4_X1 _27288_ ( .A1(_04146_ ), .A2(_04036_ ), .A3(_06466_ ), .A4(_04113_ ), .ZN(_06467_ ) );
OR3_X1 _27289_ ( .A1(_04028_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04918_ ), .ZN(_06468_ ) );
AND3_X1 _27290_ ( .A1(_06465_ ), .A2(_06467_ ), .A3(_06468_ ), .ZN(_06469_ ) );
OAI21_X1 _27291_ ( .A(_06469_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04136_ ), .ZN(_06470_ ) );
OAI21_X1 _27292_ ( .A(_04302_ ), .B1(_04140_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06471_ ) );
OAI21_X1 _27293_ ( .A(_06439_ ), .B1(_06470_ ), .B2(_06471_ ), .ZN(_06472_ ) );
OR3_X1 _27294_ ( .A1(_04131_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04181_ ), .ZN(_06473_ ) );
INV_X1 _27295_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06474_ ) );
NAND4_X1 _27296_ ( .A1(_04216_ ), .A2(_04156_ ), .A3(_06474_ ), .A4(_04174_ ), .ZN(_06475_ ) );
AND3_X1 _27297_ ( .A1(_06472_ ), .A2(_06473_ ), .A3(_06475_ ), .ZN(_06476_ ) );
OR3_X1 _27298_ ( .A1(_05653_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04190_ ), .ZN(_06477_ ) );
OR4_X1 _27299_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_04178_ ), .A3(_04181_ ), .A4(_04437_ ), .ZN(_06478_ ) );
NAND3_X1 _27300_ ( .A1(_06476_ ), .A2(_06477_ ), .A3(_06478_ ), .ZN(_06479_ ) );
NOR3_X1 _27301_ ( .A1(_04187_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04320_ ), .ZN(_06480_ ) );
INV_X1 _27302_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06481_ ) );
AND4_X1 _27303_ ( .A1(_04000_ ), .A2(_04196_ ), .A3(_06481_ ), .A4(_10756_ ), .ZN(_06482_ ) );
NOR3_X1 _27304_ ( .A1(_06479_ ), .A2(_06480_ ), .A3(_06482_ ), .ZN(_06483_ ) );
OR3_X1 _27305_ ( .A1(_04326_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04191_ ), .ZN(_06484_ ) );
OR4_X1 _27306_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_05554_ ), .A3(_04316_ ), .A4(_04318_ ), .ZN(_06485_ ) );
NAND3_X1 _27307_ ( .A1(_06483_ ), .A2(_06484_ ), .A3(_06485_ ), .ZN(_06486_ ) );
NOR3_X1 _27308_ ( .A1(_05202_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04819_ ), .ZN(_06487_ ) );
INV_X1 _27309_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06488_ ) );
AND3_X1 _27310_ ( .A1(_04215_ ), .A2(_06488_ ), .A3(_04223_ ), .ZN(_06489_ ) );
NOR3_X1 _27311_ ( .A1(_06486_ ), .A2(_06487_ ), .A3(_06489_ ), .ZN(_06490_ ) );
INV_X1 _27312_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06491_ ) );
OAI211_X1 _27313_ ( .A(_04215_ ), .B(_10792_ ), .C1(_06491_ ), .C2(_04455_ ), .ZN(_06492_ ) );
AOI221_X4 _27314_ ( .A(_04239_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B2(_04249_ ), .C1(_06490_ ), .C2(_06492_ ), .ZN(_06493_ ) );
OR2_X1 _27315_ ( .A1(_06438_ ), .A2(_06493_ ), .ZN(\idu.io_out_bits_rs1_data [23] ) );
OR2_X1 _27316_ ( .A1(_06432_ ), .A2(_06433_ ), .ZN(\lsu.io_out_bits_rd_wdata [23] ) );
AOI21_X1 _27317_ ( .A(_04738_ ), .B1(_03818_ ), .B2(_03819_ ), .ZN(_06494_ ) );
OAI22_X1 _27318_ ( .A1(_05635_ ), .A2(_04370_ ), .B1(_03909_ ), .B2(_05634_ ), .ZN(_06495_ ) );
AOI22_X1 _27319_ ( .A1(_03897_ ), .A2(\lsu.io_in_bits_lh ), .B1(_06495_ ), .B2(\arbiter.io_lsu_arsize [1] ), .ZN(_06496_ ) );
AOI21_X1 _27320_ ( .A(_04351_ ), .B1(_04358_ ), .B2(_06496_ ), .ZN(_06497_ ) );
AND2_X1 _27321_ ( .A1(_04351_ ), .A2(\lsu.io_in_bits_rd_wdata [22] ), .ZN(_06498_ ) );
OAI21_X1 _27322_ ( .A(_04353_ ), .B1(_06497_ ), .B2(_06498_ ), .ZN(_06499_ ) );
OAI211_X1 _27323_ ( .A(\wbu.io_in_bits_rd_wdata [22] ), .B(_04656_ ), .C1(_04657_ ), .C2(_04658_ ), .ZN(_06500_ ) );
AOI21_X1 _27324_ ( .A(_04356_ ), .B1(_06499_ ), .B2(_06500_ ), .ZN(_06501_ ) );
OAI21_X1 _27325_ ( .A(_03850_ ), .B1(_06494_ ), .B2(_06501_ ), .ZN(_06502_ ) );
NAND3_X1 _27326_ ( .A1(_04571_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_04243_ ), .ZN(_06503_ ) );
NAND3_X1 _27327_ ( .A1(_04444_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04542_ ), .ZN(_06504_ ) );
INV_X1 _27328_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_06505_ ) );
NAND3_X1 _27329_ ( .A1(_04134_ ), .A2(_06505_ ), .A3(_11099_ ), .ZN(_06506_ ) );
OAI21_X1 _27330_ ( .A(_06506_ ), .B1(_05293_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06507_ ) );
INV_X1 _27331_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06508_ ) );
AOI21_X1 _27332_ ( .A(_06507_ ), .B1(_06508_ ), .B2(_04392_ ), .ZN(_06509_ ) );
OR2_X1 _27333_ ( .A1(_04070_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06510_ ) );
INV_X1 _27334_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06511_ ) );
NAND4_X1 _27335_ ( .A1(_04107_ ), .A2(_04154_ ), .A3(_06511_ ), .A4(_11100_ ), .ZN(_06512_ ) );
AND3_X1 _27336_ ( .A1(_06509_ ), .A2(_06510_ ), .A3(_06512_ ), .ZN(_06513_ ) );
OR3_X1 _27337_ ( .A1(_05372_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04127_ ), .ZN(_06514_ ) );
INV_X1 _27338_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06515_ ) );
NAND4_X1 _27339_ ( .A1(_04145_ ), .A2(_04858_ ), .A3(_06515_ ), .A4(_04282_ ), .ZN(_06516_ ) );
NAND3_X1 _27340_ ( .A1(_06513_ ), .A2(_06514_ ), .A3(_06516_ ), .ZN(_06517_ ) );
NOR3_X1 _27341_ ( .A1(_04592_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04138_ ), .ZN(_06518_ ) );
INV_X1 _27342_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06519_ ) );
AND3_X1 _27343_ ( .A1(_04257_ ), .A2(_06519_ ), .A3(_04384_ ), .ZN(_06520_ ) );
NOR3_X1 _27344_ ( .A1(_06517_ ), .A2(_06518_ ), .A3(_06520_ ), .ZN(_06521_ ) );
INV_X1 _27345_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06522_ ) );
NAND3_X1 _27346_ ( .A1(_04048_ ), .A2(_06522_ ), .A3(_04113_ ), .ZN(_06523_ ) );
OR4_X1 _27347_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_05437_ ), .A3(_04124_ ), .A4(_04017_ ), .ZN(_06524_ ) );
AND3_X1 _27348_ ( .A1(_06521_ ), .A2(_06523_ ), .A3(_06524_ ), .ZN(_06525_ ) );
OR3_X1 _27349_ ( .A1(_05201_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04163_ ), .ZN(_06526_ ) );
INV_X1 _27350_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06527_ ) );
NAND4_X1 _27351_ ( .A1(_04109_ ), .A2(_04111_ ), .A3(_06527_ ), .A4(_04114_ ), .ZN(_06528_ ) );
NAND3_X1 _27352_ ( .A1(_06525_ ), .A2(_06526_ ), .A3(_06528_ ), .ZN(_06529_ ) );
INV_X1 _27353_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06530_ ) );
AND4_X1 _27354_ ( .A1(_06530_ ), .A2(_04169_ ), .A3(_04036_ ), .A4(_04513_ ), .ZN(_06531_ ) );
OAI21_X1 _27355_ ( .A(_05880_ ), .B1(_04707_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06532_ ) );
NOR3_X1 _27356_ ( .A1(_06529_ ), .A2(_06531_ ), .A3(_06532_ ), .ZN(_06533_ ) );
AND3_X1 _27357_ ( .A1(_04027_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04253_ ), .ZN(_06534_ ) );
OAI221_X1 _27358_ ( .A(_04711_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04136_ ), .C1(_06533_ ), .C2(_06534_ ), .ZN(_06535_ ) );
NAND4_X1 _27359_ ( .A1(_04171_ ), .A2(_04525_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04310_ ), .ZN(_06536_ ) );
AND2_X1 _27360_ ( .A1(_06535_ ), .A2(_06536_ ), .ZN(_06537_ ) );
OAI21_X1 _27361_ ( .A(_04428_ ), .B1(_04303_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06538_ ) );
OAI21_X1 _27362_ ( .A(_06504_ ), .B1(_06537_ ), .B2(_06538_ ), .ZN(_06539_ ) );
OR3_X1 _27363_ ( .A1(_05325_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04191_ ), .ZN(_06540_ ) );
OR3_X1 _27364_ ( .A1(_05653_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04191_ ), .ZN(_06541_ ) );
NAND3_X1 _27365_ ( .A1(_06539_ ), .A2(_06540_ ), .A3(_06541_ ), .ZN(_06542_ ) );
INV_X1 _27366_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06543_ ) );
AND4_X1 _27367_ ( .A1(_06543_ ), .A2(_04242_ ), .A3(_04542_ ), .A4(_04623_ ), .ZN(_06544_ ) );
NOR3_X1 _27368_ ( .A1(_04188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04327_ ), .ZN(_06545_ ) );
NOR3_X1 _27369_ ( .A1(_06542_ ), .A2(_06544_ ), .A3(_06545_ ), .ZN(_06546_ ) );
INV_X1 _27370_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06547_ ) );
NAND4_X1 _27371_ ( .A1(_04197_ ), .A2(_04194_ ), .A3(_06547_ ), .A4(_04455_ ), .ZN(_06548_ ) );
INV_X1 _27372_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06549_ ) );
NAND4_X1 _27373_ ( .A1(_04620_ ), .A2(_04728_ ), .A3(_06549_ ), .A4(_04211_ ), .ZN(_06550_ ) );
NAND3_X1 _27374_ ( .A1(_06546_ ), .A2(_06548_ ), .A3(_06550_ ), .ZN(_06551_ ) );
NOR4_X1 _27375_ ( .A1(_05554_ ), .A2(_04544_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_04550_ ), .ZN(_06552_ ) );
INV_X1 _27376_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06553_ ) );
AND4_X1 _27377_ ( .A1(_06553_ ), .A2(_04633_ ), .A3(_04621_ ), .A4(_04624_ ), .ZN(_06554_ ) );
NOR3_X1 _27378_ ( .A1(_06551_ ), .A2(_06552_ ), .A3(_06554_ ), .ZN(_06555_ ) );
OAI21_X1 _27379_ ( .A(_06555_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_04219_ ), .ZN(_06556_ ) );
AOI211_X1 _27380_ ( .A(_04015_ ), .B(_04023_ ), .C1(_04005_ ), .C2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06557_ ) );
OAI211_X1 _27381_ ( .A(_04247_ ), .B(_06503_ ), .C1(_06556_ ), .C2(_06557_ ), .ZN(_06558_ ) );
NAND2_X1 _27382_ ( .A1(_06502_ ), .A2(_06558_ ), .ZN(\idu.io_out_bits_rs1_data [22] ) );
OR2_X1 _27383_ ( .A1(_06497_ ), .A2(_06498_ ), .ZN(\lsu.io_out_bits_rd_wdata [22] ) );
NAND2_X1 _27384_ ( .A1(_03918_ ), .A2(_03928_ ), .ZN(\lsu.io_out_bits_rd_wdata [31] ) );
NOR4_X1 _27385_ ( .A1(_10811_ ), .A2(_10803_ ), .A3(_10813_ ), .A4(_03853_ ), .ZN(_06559_ ) );
AND2_X2 _27386_ ( .A1(_10817_ ), .A2(_06559_ ), .ZN(_06560_ ) );
OAI21_X1 _27387_ ( .A(_06560_ ), .B1(_01526_ ), .B2(_01527_ ), .ZN(_06561_ ) );
NAND3_X1 _27388_ ( .A1(_04003_ ), .A2(\idu.io_in_bits_inst [24] ), .A3(_08571_ ), .ZN(_06562_ ) );
OAI21_X1 _27389_ ( .A(\wbu.io_in_bits_rd [3] ), .B1(_11082_ ), .B2(_10614_ ), .ZN(_06563_ ) );
NOR3_X1 _27390_ ( .A1(_11082_ ), .A2(_10614_ ), .A3(\wbu.io_in_bits_rd [3] ), .ZN(_06564_ ) );
INV_X1 _27391_ ( .A(_06564_ ), .ZN(_06565_ ) );
NAND3_X1 _27392_ ( .A1(_04003_ ), .A2(\idu.io_in_bits_inst [22] ), .A3(_13006_ ), .ZN(_06566_ ) );
OAI21_X1 _27393_ ( .A(\wbu.io_in_bits_rd [2] ), .B1(_11082_ ), .B2(_10613_ ), .ZN(_06567_ ) );
AND4_X1 _27394_ ( .A1(_06563_ ), .A2(_06565_ ), .A3(_06566_ ), .A4(_06567_ ), .ZN(_06568_ ) );
OAI21_X1 _27395_ ( .A(fanout_net_36 ), .B1(_11082_ ), .B2(_10619_ ), .ZN(_06569_ ) );
OAI21_X1 _27396_ ( .A(\wbu.io_in_bits_rd [1] ), .B1(_11082_ ), .B2(_10617_ ), .ZN(_06570_ ) );
NAND3_X1 _27397_ ( .A1(_04003_ ), .A2(\idu.io_in_bits_inst [21] ), .A3(_08576_ ), .ZN(_06571_ ) );
NAND3_X1 _27398_ ( .A1(_04003_ ), .A2(\idu.io_in_bits_inst [20] ), .A3(_12972_ ), .ZN(_06572_ ) );
OAI21_X1 _27399_ ( .A(\wbu.io_in_bits_rd [0] ), .B1(_11082_ ), .B2(_10616_ ), .ZN(_06573_ ) );
AND4_X1 _27400_ ( .A1(_06570_ ), .A2(_06571_ ), .A3(_06572_ ), .A4(_06573_ ), .ZN(_06574_ ) );
AND4_X1 _27401_ ( .A1(_06562_ ), .A2(_06568_ ), .A3(_06569_ ), .A4(_06574_ ), .ZN(_06575_ ) );
AND4_X1 _27402_ ( .A1(_04235_ ), .A2(_06575_ ), .A3(_13180_ ), .A4(_13182_ ), .ZN(_06576_ ) );
NAND2_X1 _27403_ ( .A1(_03990_ ), .A2(_06576_ ), .ZN(_06577_ ) );
OAI21_X1 _27404_ ( .A(_10786_ ), .B1(_03920_ ), .B2(_03922_ ), .ZN(_06578_ ) );
AOI21_X1 _27405_ ( .A(_06578_ ), .B1(_08569_ ), .B2(_08567_ ), .ZN(_06579_ ) );
AOI211_X1 _27406_ ( .A(_12958_ ), .B(_06577_ ), .C1(_06579_ ), .C2(_10755_ ), .ZN(_06580_ ) );
AND2_X1 _27407_ ( .A1(_06579_ ), .A2(_10755_ ), .ZN(_06581_ ) );
AOI21_X1 _27408_ ( .A(_06580_ ), .B1(\lsu.io_out_bits_rd_wdata [31] ), .B2(_06581_ ), .ZN(_06582_ ) );
AOI21_X1 _27409_ ( .A(_06560_ ), .B1(_06579_ ), .B2(_10755_ ), .ZN(_06583_ ) );
NAND2_X1 _27410_ ( .A1(_06583_ ), .A2(_06577_ ), .ZN(_06584_ ) );
AND2_X1 _27411_ ( .A1(\idu.immI [1] ), .A2(\idu.io_in_bits_inst [20] ), .ZN(_06585_ ) );
CLKBUF_X3 _27412_ ( .A(_06585_ ), .Z(_06586_ ) );
CLKBUF_X2 _27413_ ( .A(_06586_ ), .Z(_06587_ ) );
AND2_X1 _27414_ ( .A1(\idu.immI [3] ), .A2(\idu.io_in_bits_inst [22] ), .ZN(_06588_ ) );
BUF_X2 _27415_ ( .A(_06588_ ), .Z(_06589_ ) );
AND2_X2 _27416_ ( .A1(_06587_ ), .A2(_06589_ ), .ZN(_06590_ ) );
BUF_X4 _27417_ ( .A(_06590_ ), .Z(_06591_ ) );
CLKBUF_X2 _27418_ ( .A(_11121_ ), .Z(_06592_ ) );
BUF_X2 _27419_ ( .A(_06592_ ), .Z(_06593_ ) );
BUF_X2 _27420_ ( .A(_06593_ ), .Z(_06594_ ) );
BUF_X2 _27421_ ( .A(_06594_ ), .Z(_06595_ ) );
BUF_X4 _27422_ ( .A(_06595_ ), .Z(_06596_ ) );
BUF_X4 _27423_ ( .A(_06596_ ), .Z(_06597_ ) );
AND2_X2 _27424_ ( .A1(_06591_ ), .A2(_06597_ ), .ZN(_06598_ ) );
INV_X1 _27425_ ( .A(_06598_ ), .ZN(_06599_ ) );
BUF_X2 _27426_ ( .A(_06599_ ), .Z(_06600_ ) );
AND2_X2 _27427_ ( .A1(\idu.immI [3] ), .A2(_10613_ ), .ZN(_06601_ ) );
AND2_X1 _27428_ ( .A1(_06601_ ), .A2(_10618_ ), .ZN(_06602_ ) );
BUF_X2 _27429_ ( .A(_06602_ ), .Z(_06603_ ) );
BUF_X2 _27430_ ( .A(_06603_ ), .Z(_06604_ ) );
BUF_X2 _27431_ ( .A(_11125_ ), .Z(_06605_ ) );
BUF_X4 _27432_ ( .A(_06605_ ), .Z(_06606_ ) );
BUF_X4 _27433_ ( .A(_06606_ ), .Z(_06607_ ) );
NAND3_X1 _27434_ ( .A1(_06604_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06607_ ), .ZN(_06608_ ) );
BUF_X4 _27435_ ( .A(_03832_ ), .Z(_06609_ ) );
BUF_X4 _27436_ ( .A(_06609_ ), .Z(_06610_ ) );
BUF_X2 _27437_ ( .A(_06610_ ), .Z(_06611_ ) );
BUF_X2 _27438_ ( .A(_06611_ ), .Z(_06612_ ) );
OR3_X1 _27439_ ( .A1(_11127_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06612_ ), .ZN(_06613_ ) );
AND2_X2 _27440_ ( .A1(_06586_ ), .A2(_06601_ ), .ZN(_06614_ ) );
NAND3_X1 _27441_ ( .A1(_06614_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06610_ ), .ZN(_06615_ ) );
NAND3_X1 _27442_ ( .A1(_10651_ ), .A2(_04056_ ), .A3(_10621_ ), .ZN(_06616_ ) );
MUX2_X1 _27443_ ( .A(_06616_ ), .B(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(_10687_ ), .Z(_06617_ ) );
AND2_X1 _27444_ ( .A1(_06585_ ), .A2(_10615_ ), .ZN(_06618_ ) );
AND2_X2 _27445_ ( .A1(_06618_ ), .A2(_10621_ ), .ZN(_06619_ ) );
INV_X1 _27446_ ( .A(_06619_ ), .ZN(_06620_ ) );
MUX2_X1 _27447_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_06617_ ), .S(_06620_ ), .Z(_06621_ ) );
AND2_X1 _27448_ ( .A1(\idu.immI [2] ), .A2(_10614_ ), .ZN(_06622_ ) );
AND2_X1 _27449_ ( .A1(_06622_ ), .A2(_10618_ ), .ZN(_06623_ ) );
INV_X1 _27450_ ( .A(_06623_ ), .ZN(_06624_ ) );
BUF_X2 _27451_ ( .A(_06624_ ), .Z(_06625_ ) );
OR3_X1 _27452_ ( .A1(_06625_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10783_ ), .ZN(_06626_ ) );
BUF_X2 _27453_ ( .A(_10650_ ), .Z(_06627_ ) );
BUF_X2 _27454_ ( .A(_06622_ ), .Z(_06628_ ) );
NAND4_X1 _27455_ ( .A1(_06627_ ), .A2(_06628_ ), .A3(_04072_ ), .A4(_11050_ ), .ZN(_06629_ ) );
NAND3_X1 _27456_ ( .A1(_06621_ ), .A2(_06626_ ), .A3(_06629_ ), .ZN(_06630_ ) );
AND2_X2 _27457_ ( .A1(_10685_ ), .A2(_06622_ ), .ZN(_06631_ ) );
AND2_X1 _27458_ ( .A1(_06631_ ), .A2(_11049_ ), .ZN(_06632_ ) );
INV_X1 _27459_ ( .A(_06632_ ), .ZN(_06633_ ) );
MUX2_X1 _27460_ ( .A(_04079_ ), .B(_06630_ ), .S(_06633_ ), .Z(_06634_ ) );
AND2_X1 _27461_ ( .A1(_06585_ ), .A2(_06622_ ), .ZN(_06635_ ) );
INV_X1 _27462_ ( .A(_06635_ ), .ZN(_06636_ ) );
BUF_X2 _27463_ ( .A(_06636_ ), .Z(_06637_ ) );
BUF_X2 _27464_ ( .A(_10812_ ), .Z(_06638_ ) );
NOR3_X1 _27465_ ( .A1(_06637_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06638_ ), .ZN(_06639_ ) );
INV_X1 _27466_ ( .A(_06602_ ), .ZN(_06640_ ) );
BUF_X4 _27467_ ( .A(_06640_ ), .Z(_06641_ ) );
NOR3_X1 _27468_ ( .A1(_06641_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06638_ ), .ZN(_06642_ ) );
NOR3_X1 _27469_ ( .A1(_06634_ ), .A2(_06639_ ), .A3(_06642_ ), .ZN(_06643_ ) );
AND2_X1 _27470_ ( .A1(_10650_ ), .A2(_06601_ ), .ZN(_06644_ ) );
AND2_X1 _27471_ ( .A1(_06644_ ), .A2(_11050_ ), .ZN(_06645_ ) );
INV_X1 _27472_ ( .A(_06645_ ), .ZN(_06646_ ) );
BUF_X2 _27473_ ( .A(_06646_ ), .Z(_06647_ ) );
OAI21_X1 _27474_ ( .A(_06643_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06647_ ), .ZN(_06648_ ) );
AND2_X1 _27475_ ( .A1(_06614_ ), .A2(_11051_ ), .ZN(_06649_ ) );
INV_X1 _27476_ ( .A(_06649_ ), .ZN(_06650_ ) );
BUF_X4 _27477_ ( .A(_06650_ ), .Z(_06651_ ) );
AND2_X1 _27478_ ( .A1(_10685_ ), .A2(_06601_ ), .ZN(_06652_ ) );
CLKBUF_X2 _27479_ ( .A(_11049_ ), .Z(_06653_ ) );
AND2_X1 _27480_ ( .A1(_06652_ ), .A2(_06653_ ), .ZN(_06654_ ) );
INV_X1 _27481_ ( .A(_06654_ ), .ZN(_06655_ ) );
OAI21_X1 _27482_ ( .A(_06651_ ), .B1(_06655_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06656_ ) );
OAI21_X1 _27483_ ( .A(_06615_ ), .B1(_06648_ ), .B2(_06656_ ), .ZN(_06657_ ) );
AND2_X2 _27484_ ( .A1(_06588_ ), .A2(_10618_ ), .ZN(_06658_ ) );
AND2_X1 _27485_ ( .A1(_06658_ ), .A2(_06653_ ), .ZN(_06659_ ) );
INV_X1 _27486_ ( .A(_06659_ ), .ZN(_06660_ ) );
BUF_X2 _27487_ ( .A(_06660_ ), .Z(_06661_ ) );
MUX2_X1 _27488_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_06657_ ), .S(_06661_ ), .Z(_06662_ ) );
BUF_X4 _27489_ ( .A(_06627_ ), .Z(_06663_ ) );
BUF_X4 _27490_ ( .A(_06663_ ), .Z(_06664_ ) );
BUF_X4 _27491_ ( .A(_06664_ ), .Z(_06665_ ) );
BUF_X2 _27492_ ( .A(_06589_ ), .Z(_06666_ ) );
NAND4_X1 _27493_ ( .A1(_06665_ ), .A2(_06666_ ), .A3(_04112_ ), .A4(_03835_ ), .ZN(_06667_ ) );
BUF_X2 _27494_ ( .A(_10685_ ), .Z(_06668_ ) );
BUF_X2 _27495_ ( .A(_06668_ ), .Z(_06669_ ) );
BUF_X2 _27496_ ( .A(_06669_ ), .Z(_06670_ ) );
NAND4_X1 _27497_ ( .A1(_06670_ ), .A2(_06666_ ), .A3(_04120_ ), .A4(_03835_ ), .ZN(_06671_ ) );
NAND3_X1 _27498_ ( .A1(_06662_ ), .A2(_06667_ ), .A3(_06671_ ), .ZN(_06672_ ) );
BUF_X2 _27499_ ( .A(_11050_ ), .Z(_06673_ ) );
BUF_X2 _27500_ ( .A(_06673_ ), .Z(_06674_ ) );
AND2_X1 _27501_ ( .A1(_06590_ ), .A2(_06674_ ), .ZN(_06675_ ) );
INV_X1 _27502_ ( .A(_06675_ ), .ZN(_06676_ ) );
BUF_X2 _27503_ ( .A(_06676_ ), .Z(_06677_ ) );
NOR2_X1 _27504_ ( .A1(_06677_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06678_ ) );
BUF_X2 _27505_ ( .A(_10651_ ), .Z(_06679_ ) );
AND2_X1 _27506_ ( .A1(_06679_ ), .A2(_11124_ ), .ZN(_06680_ ) );
INV_X1 _27507_ ( .A(_06680_ ), .ZN(_06681_ ) );
BUF_X2 _27508_ ( .A(_10615_ ), .Z(_06682_ ) );
CLKBUF_X2 _27509_ ( .A(_10618_ ), .Z(_06683_ ) );
AND2_X2 _27510_ ( .A1(_06682_ ), .A2(_06683_ ), .ZN(_06684_ ) );
AND2_X1 _27511_ ( .A1(_06684_ ), .A2(_06638_ ), .ZN(_06685_ ) );
INV_X1 _27512_ ( .A(_06685_ ), .ZN(_06686_ ) );
BUF_X2 _27513_ ( .A(_06686_ ), .Z(_06687_ ) );
OAI21_X1 _27514_ ( .A(_06681_ ), .B1(_06687_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06688_ ) );
NOR3_X1 _27515_ ( .A1(_06672_ ), .A2(_06678_ ), .A3(_06688_ ), .ZN(_06689_ ) );
CLKBUF_X2 _27516_ ( .A(_06593_ ), .Z(_06690_ ) );
BUF_X2 _27517_ ( .A(_06690_ ), .Z(_06691_ ) );
AND3_X1 _27518_ ( .A1(_06679_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06691_ ), .ZN(_06692_ ) );
OAI21_X1 _27519_ ( .A(_06613_ ), .B1(_06689_ ), .B2(_06692_ ), .ZN(_06693_ ) );
BUF_X2 _27520_ ( .A(_06618_ ), .Z(_06694_ ) );
AND3_X1 _27521_ ( .A1(_06694_ ), .A2(_04143_ ), .A3(_01099_ ), .ZN(_06695_ ) );
BUF_X2 _27522_ ( .A(_06628_ ), .Z(_06696_ ) );
BUF_X2 _27523_ ( .A(_06696_ ), .Z(_06697_ ) );
BUF_X2 _27524_ ( .A(_06697_ ), .Z(_06698_ ) );
BUF_X2 _27525_ ( .A(_06683_ ), .Z(_06699_ ) );
AND4_X1 _27526_ ( .A1(_04153_ ), .A2(_06698_ ), .A3(_06699_ ), .A4(_06691_ ), .ZN(_06700_ ) );
NOR3_X1 _27527_ ( .A1(_06693_ ), .A2(_06695_ ), .A3(_06700_ ), .ZN(_06701_ ) );
AND2_X1 _27528_ ( .A1(_10650_ ), .A2(_06622_ ), .ZN(_06702_ ) );
BUF_X2 _27529_ ( .A(_06702_ ), .Z(_06703_ ) );
AND2_X1 _27530_ ( .A1(_06703_ ), .A2(_06594_ ), .ZN(_06704_ ) );
INV_X1 _27531_ ( .A(_06704_ ), .ZN(_06705_ ) );
CLKBUF_X2 _27532_ ( .A(_06705_ ), .Z(_06706_ ) );
OR2_X1 _27533_ ( .A1(_06706_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06707_ ) );
BUF_X4 _27534_ ( .A(_06670_ ), .Z(_06708_ ) );
BUF_X4 _27535_ ( .A(_06708_ ), .Z(_06709_ ) );
BUF_X4 _27536_ ( .A(_06698_ ), .Z(_06710_ ) );
BUF_X4 _27537_ ( .A(_06710_ ), .Z(_06711_ ) );
NAND4_X1 _27538_ ( .A1(_06709_ ), .A2(_06711_ ), .A3(_04172_ ), .A4(_01100_ ), .ZN(_06712_ ) );
NAND3_X1 _27539_ ( .A1(_06701_ ), .A2(_06707_ ), .A3(_06712_ ), .ZN(_06713_ ) );
AND2_X1 _27540_ ( .A1(_06603_ ), .A2(_06595_ ), .ZN(_06714_ ) );
INV_X1 _27541_ ( .A(_06714_ ), .ZN(_06715_ ) );
AND2_X1 _27542_ ( .A1(_06635_ ), .A2(_06605_ ), .ZN(_06716_ ) );
INV_X1 _27543_ ( .A(_06716_ ), .ZN(_06717_ ) );
OAI21_X1 _27544_ ( .A(_06715_ ), .B1(_06717_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06718_ ) );
OAI21_X1 _27545_ ( .A(_06608_ ), .B1(_06713_ ), .B2(_06718_ ), .ZN(_06719_ ) );
BUF_X2 _27546_ ( .A(_06664_ ), .Z(_06720_ ) );
BUF_X4 _27547_ ( .A(_06720_ ), .Z(_06721_ ) );
BUF_X4 _27548_ ( .A(_06721_ ), .Z(_06722_ ) );
BUF_X2 _27549_ ( .A(_06601_ ), .Z(_06723_ ) );
BUF_X4 _27550_ ( .A(_06723_ ), .Z(_06724_ ) );
BUF_X4 _27551_ ( .A(_06724_ ), .Z(_06725_ ) );
BUF_X2 _27552_ ( .A(_06725_ ), .Z(_06726_ ) );
BUF_X4 _27553_ ( .A(_06726_ ), .Z(_06727_ ) );
BUF_X4 _27554_ ( .A(_06597_ ), .Z(_06728_ ) );
NAND4_X1 _27555_ ( .A1(_06722_ ), .A2(_06727_ ), .A3(_04198_ ), .A4(_06728_ ), .ZN(_06729_ ) );
CLKBUF_X2 _27556_ ( .A(_06652_ ), .Z(_06730_ ) );
AND2_X2 _27557_ ( .A1(_06730_ ), .A2(_06691_ ), .ZN(_06731_ ) );
INV_X1 _27558_ ( .A(_06731_ ), .ZN(_06732_ ) );
OR2_X1 _27559_ ( .A1(_06732_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06733_ ) );
NAND3_X1 _27560_ ( .A1(_06719_ ), .A2(_06729_ ), .A3(_06733_ ), .ZN(_06734_ ) );
BUF_X2 _27561_ ( .A(_06614_ ), .Z(_06735_ ) );
AND2_X1 _27562_ ( .A1(_06735_ ), .A2(_01099_ ), .ZN(_06736_ ) );
INV_X1 _27563_ ( .A(_06736_ ), .ZN(_06737_ ) );
BUF_X2 _27564_ ( .A(_06737_ ), .Z(_06738_ ) );
NOR2_X1 _27565_ ( .A1(_06738_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06739_ ) );
BUF_X2 _27566_ ( .A(_06658_ ), .Z(_06740_ ) );
BUF_X2 _27567_ ( .A(_11125_ ), .Z(_06741_ ) );
AND2_X1 _27568_ ( .A1(_06740_ ), .A2(_06741_ ), .ZN(_06742_ ) );
INV_X1 _27569_ ( .A(_06742_ ), .ZN(_06743_ ) );
NOR2_X1 _27570_ ( .A1(_06743_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06744_ ) );
AND2_X1 _27571_ ( .A1(_10685_ ), .A2(_06589_ ), .ZN(_06745_ ) );
AND2_X1 _27572_ ( .A1(_06745_ ), .A2(_06691_ ), .ZN(_06746_ ) );
BUF_X4 _27573_ ( .A(_06746_ ), .Z(_06747_ ) );
INV_X1 _27574_ ( .A(_06747_ ), .ZN(_06748_ ) );
AND2_X2 _27575_ ( .A1(_10650_ ), .A2(_06589_ ), .ZN(_06749_ ) );
BUF_X4 _27576_ ( .A(_06691_ ), .Z(_06750_ ) );
AND2_X1 _27577_ ( .A1(_06749_ ), .A2(_06750_ ), .ZN(_06751_ ) );
INV_X1 _27578_ ( .A(_06751_ ), .ZN(_06752_ ) );
OAI21_X1 _27579_ ( .A(_06748_ ), .B1(_06752_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06753_ ) );
NOR4_X1 _27580_ ( .A1(_06734_ ), .A2(_06739_ ), .A3(_06744_ ), .A4(_06753_ ), .ZN(_06754_ ) );
BUF_X4 _27581_ ( .A(_06708_ ), .Z(_06755_ ) );
BUF_X2 _27582_ ( .A(_06755_ ), .Z(_06756_ ) );
BUF_X2 _27583_ ( .A(_06666_ ), .Z(_06757_ ) );
BUF_X2 _27584_ ( .A(_06757_ ), .Z(_06758_ ) );
AND4_X1 _27585_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A2(_06756_ ), .A3(_06758_ ), .A4(_01102_ ), .ZN(_06759_ ) );
OAI21_X1 _27586_ ( .A(_06600_ ), .B1(_06754_ ), .B2(_06759_ ), .ZN(_06760_ ) );
BUF_X4 _27587_ ( .A(_06591_ ), .Z(_06761_ ) );
NAND3_X1 _27588_ ( .A1(_06761_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(\idu.immI [4] ), .ZN(_06762_ ) );
NAND2_X1 _27589_ ( .A1(_06760_ ), .A2(_06762_ ), .ZN(_06763_ ) );
OAI221_X1 _27590_ ( .A(_06561_ ), .B1(_06560_ ), .B2(_06582_ ), .C1(_06584_ ), .C2(_06763_ ), .ZN(\idu.io_out_bits_rs2_data [31] ) );
INV_X1 _27591_ ( .A(_03854_ ), .ZN(_06764_ ) );
NOR2_X1 _27592_ ( .A1(_06764_ ), .A2(_10814_ ), .ZN(_06765_ ) );
BUF_X4 _27593_ ( .A(_06765_ ), .Z(_06766_ ) );
BUF_X4 _27594_ ( .A(_06766_ ), .Z(_06767_ ) );
OAI21_X1 _27595_ ( .A(_06767_ ), .B1(_01717_ ), .B2(_01719_ ), .ZN(_06768_ ) );
OAI211_X1 _27596_ ( .A(_10786_ ), .B(_10755_ ), .C1(_03920_ ), .C2(_03922_ ), .ZN(_06769_ ) );
OR2_X1 _27597_ ( .A1(_08570_ ), .A2(_06769_ ), .ZN(_06770_ ) );
BUF_X2 _27598_ ( .A(_06770_ ), .Z(_06771_ ) );
INV_X1 _27599_ ( .A(_06765_ ), .ZN(_06772_ ) );
BUF_X4 _27600_ ( .A(_06772_ ), .Z(_06773_ ) );
AOI21_X1 _27601_ ( .A(_06564_ ), .B1(_11067_ ), .B2(\wbu.io_in_bits_rd [1] ), .ZN(_06774_ ) );
AND4_X1 _27602_ ( .A1(_04235_ ), .A2(_12964_ ), .A3(_06563_ ), .A4(_06774_ ), .ZN(_06775_ ) );
AND3_X1 _27603_ ( .A1(_06566_ ), .A2(_06562_ ), .A3(_06567_ ), .ZN(_06776_ ) );
AND4_X1 _27604_ ( .A1(_06573_ ), .A2(_06571_ ), .A3(_06572_ ), .A4(_06569_ ), .ZN(_06777_ ) );
NAND3_X1 _27605_ ( .A1(_06775_ ), .A2(_06776_ ), .A3(_06777_ ), .ZN(_06778_ ) );
NOR2_X1 _27606_ ( .A1(_03989_ ), .A2(_06778_ ), .ZN(_06779_ ) );
CLKBUF_X2 _27607_ ( .A(_06779_ ), .Z(_06780_ ) );
AND4_X1 _27608_ ( .A1(\wbu.io_in_bits_rd_wdata [30] ), .A2(_06771_ ), .A3(_06773_ ), .A4(_06780_ ), .ZN(_06781_ ) );
CLKBUF_X2 _27609_ ( .A(_06770_ ), .Z(_06782_ ) );
NOR2_X2 _27610_ ( .A1(_06782_ ), .A2(_06766_ ), .ZN(_06783_ ) );
BUF_X4 _27611_ ( .A(_06783_ ), .Z(_06784_ ) );
AOI21_X1 _27612_ ( .A(_06781_ ), .B1(\lsu.io_out_bits_rd_wdata [30] ), .B2(_06784_ ), .ZN(_06785_ ) );
OR2_X1 _27613_ ( .A1(_06732_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06786_ ) );
CLKBUF_X2 _27614_ ( .A(_06674_ ), .Z(_06787_ ) );
AND3_X1 _27615_ ( .A1(_06730_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06787_ ), .ZN(_06788_ ) );
OR3_X1 _27616_ ( .A1(_11126_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11121_ ), .ZN(_06789_ ) );
INV_X1 _27617_ ( .A(_10652_ ), .ZN(_06790_ ) );
BUF_X4 _27618_ ( .A(_06790_ ), .Z(_06791_ ) );
OAI21_X1 _27619_ ( .A(_06789_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .B2(_06791_ ), .ZN(_06792_ ) );
AOI21_X1 _27620_ ( .A(_06792_ ), .B1(_04260_ ), .B2(_06619_ ), .ZN(_06793_ ) );
BUF_X2 _27621_ ( .A(_06625_ ), .Z(_06794_ ) );
OR3_X1 _27622_ ( .A1(_06794_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11122_ ), .ZN(_06795_ ) );
CLKBUF_X2 _27623_ ( .A(_11051_ ), .Z(_06796_ ) );
NAND4_X1 _27624_ ( .A1(_06663_ ), .A2(_06696_ ), .A3(_04268_ ), .A4(_06796_ ), .ZN(_06797_ ) );
AND3_X1 _27625_ ( .A1(_06793_ ), .A2(_06795_ ), .A3(_06797_ ), .ZN(_06798_ ) );
CLKBUF_X2 _27626_ ( .A(_06633_ ), .Z(_06799_ ) );
OR2_X1 _27627_ ( .A1(_06799_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06800_ ) );
NAND2_X1 _27628_ ( .A1(_06798_ ), .A2(_06800_ ), .ZN(_06801_ ) );
BUF_X4 _27629_ ( .A(_06637_ ), .Z(_06802_ ) );
NOR3_X1 _27630_ ( .A1(_06802_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06593_ ), .ZN(_06803_ ) );
BUF_X4 _27631_ ( .A(_06641_ ), .Z(_06804_ ) );
AOI211_X1 _27632_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_06804_ ), .C1(\idu.io_in_bits_inst [24] ), .C2(_04003_ ), .ZN(_06805_ ) );
NOR3_X1 _27633_ ( .A1(_06801_ ), .A2(_06803_ ), .A3(_06805_ ), .ZN(_06806_ ) );
AOI22_X1 _27634_ ( .A1(_06645_ ), .A2(_04258_ ), .B1(_03834_ ), .B2(_06730_ ), .ZN(_06807_ ) );
AOI21_X1 _27635_ ( .A(_06788_ ), .B1(_06806_ ), .B2(_06807_ ), .ZN(_06808_ ) );
BUF_X4 _27636_ ( .A(_06651_ ), .Z(_06809_ ) );
NOR2_X1 _27637_ ( .A1(_06809_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06810_ ) );
BUF_X2 _27638_ ( .A(_03833_ ), .Z(_06811_ ) );
AND3_X1 _27639_ ( .A1(_06658_ ), .A2(_04281_ ), .A3(_06811_ ), .ZN(_06812_ ) );
NOR3_X1 _27640_ ( .A1(_06808_ ), .A2(_06810_ ), .A3(_06812_ ), .ZN(_06813_ ) );
BUF_X2 _27641_ ( .A(_06673_ ), .Z(_06814_ ) );
BUF_X2 _27642_ ( .A(_06814_ ), .Z(_06815_ ) );
BUF_X2 _27643_ ( .A(_06815_ ), .Z(_06816_ ) );
BUF_X4 _27644_ ( .A(_06816_ ), .Z(_06817_ ) );
NAND4_X1 _27645_ ( .A1(_06720_ ), .A2(_06666_ ), .A3(_04286_ ), .A4(_06817_ ), .ZN(_06818_ ) );
AND2_X1 _27646_ ( .A1(_06745_ ), .A2(_06609_ ), .ZN(_06819_ ) );
INV_X1 _27647_ ( .A(_06819_ ), .ZN(_06820_ ) );
OR2_X1 _27648_ ( .A1(_06820_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06821_ ) );
NAND3_X1 _27649_ ( .A1(_06813_ ), .A2(_06818_ ), .A3(_06821_ ), .ZN(_06822_ ) );
NOR2_X1 _27650_ ( .A1(_06677_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06823_ ) );
BUF_X4 _27651_ ( .A(_06687_ ), .Z(_06824_ ) );
NOR2_X1 _27652_ ( .A1(_06824_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06825_ ) );
NOR3_X1 _27653_ ( .A1(_06822_ ), .A2(_06823_ ), .A3(_06825_ ), .ZN(_06826_ ) );
INV_X1 _27654_ ( .A(_10651_ ), .ZN(_06827_ ) );
CLKBUF_X2 _27655_ ( .A(_06827_ ), .Z(_06828_ ) );
CLKBUF_X2 _27656_ ( .A(_06828_ ), .Z(_06829_ ) );
CLKBUF_X2 _27657_ ( .A(_06829_ ), .Z(_06830_ ) );
BUF_X2 _27658_ ( .A(_06611_ ), .Z(_06831_ ) );
OR3_X1 _27659_ ( .A1(_06830_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06831_ ), .ZN(_06832_ ) );
CLKBUF_X2 _27660_ ( .A(_06682_ ), .Z(_06833_ ) );
BUF_X2 _27661_ ( .A(_06833_ ), .Z(_06834_ ) );
BUF_X4 _27662_ ( .A(_06834_ ), .Z(_06835_ ) );
NAND4_X1 _27663_ ( .A1(_06708_ ), .A2(_06835_ ), .A3(_04298_ ), .A4(_06741_ ), .ZN(_06836_ ) );
NAND3_X1 _27664_ ( .A1(_06826_ ), .A2(_06832_ ), .A3(_06836_ ), .ZN(_06837_ ) );
AND2_X1 _27665_ ( .A1(_06694_ ), .A2(_11124_ ), .ZN(_06838_ ) );
INV_X1 _27666_ ( .A(_06838_ ), .ZN(_06839_ ) );
BUF_X2 _27667_ ( .A(_06839_ ), .Z(_06840_ ) );
BUF_X4 _27668_ ( .A(_06840_ ), .Z(_06841_ ) );
NOR2_X1 _27669_ ( .A1(_06841_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06842_ ) );
CLKBUF_X2 _27670_ ( .A(_06794_ ), .Z(_06843_ ) );
BUF_X2 _27671_ ( .A(_06843_ ), .Z(_06844_ ) );
BUF_X4 _27672_ ( .A(_06610_ ), .Z(_06845_ ) );
BUF_X2 _27673_ ( .A(_06845_ ), .Z(_06846_ ) );
BUF_X2 _27674_ ( .A(_06846_ ), .Z(_06847_ ) );
NOR3_X1 _27675_ ( .A1(_06844_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06847_ ), .ZN(_06848_ ) );
NOR3_X1 _27676_ ( .A1(_06837_ ), .A2(_06842_ ), .A3(_06848_ ), .ZN(_06849_ ) );
BUF_X4 _27677_ ( .A(_06721_ ), .Z(_06850_ ) );
NAND4_X1 _27678_ ( .A1(_06850_ ), .A2(_06711_ ), .A3(_04308_ ), .A4(_06597_ ), .ZN(_06851_ ) );
BUF_X2 _27679_ ( .A(_06741_ ), .Z(_06852_ ) );
NAND4_X1 _27680_ ( .A1(_06709_ ), .A2(_06711_ ), .A3(_04312_ ), .A4(_06852_ ), .ZN(_06853_ ) );
NAND3_X1 _27681_ ( .A1(_06849_ ), .A2(_06851_ ), .A3(_06853_ ), .ZN(_06854_ ) );
BUF_X4 _27682_ ( .A(_06802_ ), .Z(_06855_ ) );
BUF_X4 _27683_ ( .A(_06847_ ), .Z(_06856_ ) );
NOR3_X1 _27684_ ( .A1(_06855_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06856_ ), .ZN(_06857_ ) );
CLKBUF_X2 _27685_ ( .A(_06644_ ), .Z(_06858_ ) );
AND2_X1 _27686_ ( .A1(_06858_ ), .A2(_01099_ ), .ZN(_06859_ ) );
INV_X1 _27687_ ( .A(_06859_ ), .ZN(_06860_ ) );
OAI21_X1 _27688_ ( .A(_06860_ ), .B1(_06715_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06861_ ) );
NOR3_X1 _27689_ ( .A1(_06854_ ), .A2(_06857_ ), .A3(_06861_ ), .ZN(_06862_ ) );
AND3_X1 _27690_ ( .A1(_06858_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01101_ ), .ZN(_06863_ ) );
OAI21_X1 _27691_ ( .A(_06786_ ), .B1(_06862_ ), .B2(_06863_ ), .ZN(_06864_ ) );
BUF_X4 _27692_ ( .A(_06750_ ), .Z(_06865_ ) );
BUF_X2 _27693_ ( .A(_06865_ ), .Z(_06866_ ) );
AND3_X1 _27694_ ( .A1(_06735_ ), .A2(_04330_ ), .A3(_06866_ ), .ZN(_06867_ ) );
NOR2_X1 _27695_ ( .A1(_06743_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06868_ ) );
OR3_X1 _27696_ ( .A1(_06864_ ), .A2(_06867_ ), .A3(_06868_ ), .ZN(_06869_ ) );
BUF_X4 _27697_ ( .A(_06752_ ), .Z(_06870_ ) );
NOR2_X1 _27698_ ( .A1(_06870_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06871_ ) );
BUF_X4 _27699_ ( .A(_06748_ ), .Z(_06872_ ) );
OAI21_X1 _27700_ ( .A(_06600_ ), .B1(_06872_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06873_ ) );
NOR3_X1 _27701_ ( .A1(_06869_ ), .A2(_06871_ ), .A3(_06873_ ), .ZN(_06874_ ) );
AND2_X2 _27702_ ( .A1(_06770_ ), .A2(_06772_ ), .ZN(_06875_ ) );
INV_X1 _27703_ ( .A(_06779_ ), .ZN(_06876_ ) );
BUF_X4 _27704_ ( .A(_06876_ ), .Z(_06877_ ) );
OAI211_X1 _27705_ ( .A(_06875_ ), .B(_06877_ ), .C1(_04248_ ), .C2(_06600_ ), .ZN(_06878_ ) );
OAI211_X1 _27706_ ( .A(_06768_ ), .B(_06785_ ), .C1(_06874_ ), .C2(_06878_ ), .ZN(\idu.io_out_bits_rs2_data [30] ) );
BUF_X4 _27707_ ( .A(_06766_ ), .Z(_06879_ ) );
NAND2_X1 _27708_ ( .A1(\exu.io_out_bits_rd_wdata [21] ), .A2(_06879_ ), .ZN(_06880_ ) );
AND4_X1 _27709_ ( .A1(\wbu.io_in_bits_rd_wdata [21] ), .A2(_06771_ ), .A3(_06773_ ), .A4(_06780_ ), .ZN(_06881_ ) );
AOI21_X1 _27710_ ( .A(_06881_ ), .B1(\lsu.io_out_bits_rd_wdata [21] ), .B2(_06784_ ), .ZN(_06882_ ) );
BUF_X2 _27711_ ( .A(_06728_ ), .Z(_06883_ ) );
NAND3_X1 _27712_ ( .A1(_06740_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06883_ ), .ZN(_06884_ ) );
BUF_X2 _27713_ ( .A(_06597_ ), .Z(_06885_ ) );
NAND3_X1 _27714_ ( .A1(_06604_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06885_ ), .ZN(_06886_ ) );
NAND3_X1 _27715_ ( .A1(_06623_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06852_ ), .ZN(_06887_ ) );
NOR2_X1 _27716_ ( .A1(_06661_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06888_ ) );
OR3_X1 _27717_ ( .A1(_11127_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06592_ ), .ZN(_06889_ ) );
OAI21_X1 _27718_ ( .A(_06889_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .B2(_06791_ ), .ZN(_06890_ ) );
AND4_X1 _27719_ ( .A1(_04391_ ), .A2(_06587_ ), .A3(_06833_ ), .A4(_06814_ ), .ZN(_06891_ ) );
NOR3_X1 _27720_ ( .A1(_06794_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11123_ ), .ZN(_06892_ ) );
NOR3_X1 _27721_ ( .A1(_06890_ ), .A2(_06891_ ), .A3(_06892_ ), .ZN(_06893_ ) );
NAND4_X1 _27722_ ( .A1(_06664_ ), .A2(_06697_ ), .A3(_04396_ ), .A4(_06610_ ), .ZN(_06894_ ) );
OR2_X1 _27723_ ( .A1(_06799_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06895_ ) );
NAND3_X1 _27724_ ( .A1(_06893_ ), .A2(_06894_ ), .A3(_06895_ ), .ZN(_06896_ ) );
BUF_X2 _27725_ ( .A(_06587_ ), .Z(_06897_ ) );
BUF_X2 _27726_ ( .A(_06897_ ), .Z(_06898_ ) );
AND4_X1 _27727_ ( .A1(_04402_ ), .A2(_06898_ ), .A3(_06697_ ), .A4(_06815_ ), .ZN(_06899_ ) );
NOR3_X1 _27728_ ( .A1(_06804_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11124_ ), .ZN(_06900_ ) );
NOR3_X1 _27729_ ( .A1(_06896_ ), .A2(_06899_ ), .A3(_06900_ ), .ZN(_06901_ ) );
NAND4_X1 _27730_ ( .A1(_06665_ ), .A2(_06725_ ), .A3(_04407_ ), .A4(_06611_ ), .ZN(_06902_ ) );
AOI22_X1 _27731_ ( .A1(_06654_ ), .A2(_04410_ ), .B1(_06845_ ), .B2(_06614_ ), .ZN(_06903_ ) );
NAND3_X1 _27732_ ( .A1(_06901_ ), .A2(_06902_ ), .A3(_06903_ ), .ZN(_06904_ ) );
NAND3_X1 _27733_ ( .A1(_06614_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06817_ ), .ZN(_06905_ ) );
AOI21_X1 _27734_ ( .A(_06888_ ), .B1(_06904_ ), .B2(_06905_ ), .ZN(_06906_ ) );
BUF_X2 _27735_ ( .A(_06665_ ), .Z(_06907_ ) );
NAND4_X1 _27736_ ( .A1(_06907_ ), .A2(_06757_ ), .A3(_04386_ ), .A4(_06831_ ), .ZN(_06908_ ) );
BUF_X2 _27737_ ( .A(_06589_ ), .Z(_06909_ ) );
BUF_X2 _27738_ ( .A(_06909_ ), .Z(_06910_ ) );
NAND4_X1 _27739_ ( .A1(_06670_ ), .A2(_06910_ ), .A3(_04419_ ), .A4(_06612_ ), .ZN(_06911_ ) );
NAND3_X1 _27740_ ( .A1(_06906_ ), .A2(_06908_ ), .A3(_06911_ ), .ZN(_06912_ ) );
NOR2_X1 _27741_ ( .A1(_06677_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06913_ ) );
AND3_X1 _27742_ ( .A1(_06684_ ), .A2(_04423_ ), .A3(_06595_ ), .ZN(_06914_ ) );
NOR3_X1 _27743_ ( .A1(_06912_ ), .A2(_06913_ ), .A3(_06914_ ), .ZN(_06915_ ) );
BUF_X4 _27744_ ( .A(_06835_ ), .Z(_06916_ ) );
NAND4_X1 _27745_ ( .A1(_06721_ ), .A2(_06916_ ), .A3(_04425_ ), .A4(_06750_ ), .ZN(_06917_ ) );
CLKBUF_X2 _27746_ ( .A(_11127_ ), .Z(_06918_ ) );
CLKBUF_X2 _27747_ ( .A(_03835_ ), .Z(_06919_ ) );
OR3_X1 _27748_ ( .A1(_06918_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06919_ ), .ZN(_06920_ ) );
NAND3_X1 _27749_ ( .A1(_06915_ ), .A2(_06917_ ), .A3(_06920_ ), .ZN(_06921_ ) );
AND2_X1 _27750_ ( .A1(_06623_ ), .A2(_06594_ ), .ZN(_06922_ ) );
INV_X1 _27751_ ( .A(_06922_ ), .ZN(_06923_ ) );
OAI21_X1 _27752_ ( .A(_06923_ ), .B1(_06841_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06924_ ) );
OAI21_X1 _27753_ ( .A(_06887_ ), .B1(_06921_ ), .B2(_06924_ ), .ZN(_06925_ ) );
BUF_X4 _27754_ ( .A(_06710_ ), .Z(_06926_ ) );
NAND4_X1 _27755_ ( .A1(_06722_ ), .A2(_06926_ ), .A3(_04382_ ), .A4(_06607_ ), .ZN(_06927_ ) );
AND2_X1 _27756_ ( .A1(_06631_ ), .A2(_06690_ ), .ZN(_06928_ ) );
INV_X1 _27757_ ( .A(_06928_ ), .ZN(_06929_ ) );
CLKBUF_X2 _27758_ ( .A(_06929_ ), .Z(_06930_ ) );
OR2_X1 _27759_ ( .A1(_06930_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06931_ ) );
NAND3_X1 _27760_ ( .A1(_06925_ ), .A2(_06927_ ), .A3(_06931_ ), .ZN(_06932_ ) );
BUF_X4 _27761_ ( .A(_06715_ ), .Z(_06933_ ) );
OAI21_X1 _27762_ ( .A(_06933_ ), .B1(_06717_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06934_ ) );
OAI21_X1 _27763_ ( .A(_06886_ ), .B1(_06932_ ), .B2(_06934_ ), .ZN(_06935_ ) );
BUF_X2 _27764_ ( .A(_06722_ ), .Z(_06936_ ) );
BUF_X2 _27765_ ( .A(_06727_ ), .Z(_06937_ ) );
BUF_X2 _27766_ ( .A(_06607_ ), .Z(_06938_ ) );
NAND4_X1 _27767_ ( .A1(_06936_ ), .A2(_06937_ ), .A3(_04441_ ), .A4(_06938_ ), .ZN(_06939_ ) );
CLKBUF_X2 _27768_ ( .A(_06732_ ), .Z(_06940_ ) );
OR2_X1 _27769_ ( .A1(_06940_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06941_ ) );
NAND3_X1 _27770_ ( .A1(_06935_ ), .A2(_06939_ ), .A3(_06941_ ), .ZN(_06942_ ) );
BUF_X2 _27771_ ( .A(_06743_ ), .Z(_06943_ ) );
BUF_X2 _27772_ ( .A(_06738_ ), .Z(_06944_ ) );
OAI21_X1 _27773_ ( .A(_06943_ ), .B1(_06944_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06945_ ) );
OAI21_X1 _27774_ ( .A(_06884_ ), .B1(_06942_ ), .B2(_06945_ ), .ZN(_06946_ ) );
BUF_X4 _27775_ ( .A(_06850_ ), .Z(_06947_ ) );
BUF_X4 _27776_ ( .A(_06947_ ), .Z(_06948_ ) );
BUF_X4 _27777_ ( .A(_06758_ ), .Z(_06949_ ) );
BUF_X4 _27778_ ( .A(_01102_ ), .Z(_06950_ ) );
NAND4_X1 _27779_ ( .A1(_06948_ ), .A2(_06949_ ), .A3(_04380_ ), .A4(_06950_ ), .ZN(_06951_ ) );
BUF_X4 _27780_ ( .A(_01102_ ), .Z(_06952_ ) );
BUF_X4 _27781_ ( .A(_06591_ ), .Z(_06953_ ) );
AOI22_X1 _27782_ ( .A1(_06747_ ), .A2(_04454_ ), .B1(_06952_ ), .B2(_06953_ ), .ZN(_06954_ ) );
AND3_X1 _27783_ ( .A1(_06946_ ), .A2(_06951_ ), .A3(_06954_ ), .ZN(_06955_ ) );
BUF_X4 _27784_ ( .A(_06771_ ), .Z(_06956_ ) );
BUF_X4 _27785_ ( .A(_06773_ ), .Z(_06957_ ) );
NAND3_X1 _27786_ ( .A1(_06761_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(\idu.immI [4] ), .ZN(_06958_ ) );
NAND4_X1 _27787_ ( .A1(_06956_ ), .A2(_06957_ ), .A3(_06877_ ), .A4(_06958_ ), .ZN(_06959_ ) );
OAI211_X1 _27788_ ( .A(_06880_ ), .B(_06882_ ), .C1(_06955_ ), .C2(_06959_ ), .ZN(\idu.io_out_bits_rs2_data [21] ) );
NAND2_X1 _27789_ ( .A1(\exu.io_out_bits_rd_wdata [20] ), .A2(_06879_ ), .ZN(_06960_ ) );
AND4_X1 _27790_ ( .A1(\wbu.io_in_bits_rd_wdata [20] ), .A2(_06771_ ), .A3(_06773_ ), .A4(_06780_ ), .ZN(_06961_ ) );
AOI21_X1 _27791_ ( .A(_06961_ ), .B1(\lsu.io_out_bits_rd_wdata [20] ), .B2(_06784_ ), .ZN(_06962_ ) );
AND4_X1 _27792_ ( .A1(_04530_ ), .A2(_06670_ ), .A3(_06835_ ), .A4(_06595_ ), .ZN(_06963_ ) );
AND4_X1 _27793_ ( .A1(_04500_ ), .A2(_10685_ ), .A3(_06628_ ), .A4(_11051_ ), .ZN(_06964_ ) );
OR3_X1 _27794_ ( .A1(_06828_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10783_ ), .ZN(_06965_ ) );
BUF_X2 _27795_ ( .A(_10686_ ), .Z(_06966_ ) );
NAND3_X1 _27796_ ( .A1(_06966_ ), .A2(_04491_ ), .A3(_06653_ ), .ZN(_06967_ ) );
NAND4_X1 _27797_ ( .A1(_06586_ ), .A2(_06682_ ), .A3(_04490_ ), .A4(_11050_ ), .ZN(_06968_ ) );
AND3_X1 _27798_ ( .A1(_06965_ ), .A2(_06967_ ), .A3(_06968_ ), .ZN(_06969_ ) );
AND2_X1 _27799_ ( .A1(_06702_ ), .A2(_11049_ ), .ZN(_06970_ ) );
INV_X1 _27800_ ( .A(_06970_ ), .ZN(_06971_ ) );
BUF_X2 _27801_ ( .A(_06971_ ), .Z(_06972_ ) );
OR3_X1 _27802_ ( .A1(_06625_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11121_ ), .ZN(_06973_ ) );
NAND3_X1 _27803_ ( .A1(_06969_ ), .A2(_06972_ ), .A3(_06973_ ), .ZN(_06974_ ) );
NAND3_X1 _27804_ ( .A1(_06703_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11052_ ), .ZN(_06975_ ) );
AOI21_X1 _27805_ ( .A(_06964_ ), .B1(_06974_ ), .B2(_06975_ ), .ZN(_06976_ ) );
OR3_X1 _27806_ ( .A1(_06636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06592_ ), .ZN(_06977_ ) );
NAND4_X1 _27807_ ( .A1(_06723_ ), .A2(_06683_ ), .A3(_04505_ ), .A4(_06814_ ), .ZN(_06978_ ) );
NAND3_X1 _27808_ ( .A1(_06976_ ), .A2(_06977_ ), .A3(_06978_ ), .ZN(_06979_ ) );
NOR2_X1 _27809_ ( .A1(_06646_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06980_ ) );
AND4_X1 _27810_ ( .A1(_04510_ ), .A2(_06668_ ), .A3(_06723_ ), .A4(_06814_ ), .ZN(_06981_ ) );
NOR3_X1 _27811_ ( .A1(_06979_ ), .A2(_06980_ ), .A3(_06981_ ), .ZN(_06982_ ) );
NAND4_X1 _27812_ ( .A1(_06898_ ), .A2(_06724_ ), .A3(_04512_ ), .A4(_06610_ ), .ZN(_06983_ ) );
OR2_X1 _27813_ ( .A1(_06660_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06984_ ) );
NAND3_X1 _27814_ ( .A1(_06982_ ), .A2(_06983_ ), .A3(_06984_ ), .ZN(_06985_ ) );
AND2_X1 _27815_ ( .A1(_06749_ ), .A2(_06673_ ), .ZN(_06986_ ) );
INV_X1 _27816_ ( .A(_06986_ ), .ZN(_06987_ ) );
BUF_X2 _27817_ ( .A(_06987_ ), .Z(_06988_ ) );
NOR2_X1 _27818_ ( .A1(_06988_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06989_ ) );
INV_X1 _27819_ ( .A(_06745_ ), .ZN(_06990_ ) );
AOI211_X1 _27820_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_06990_ ), .C1(\idu.io_in_bits_inst [24] ), .C2(_04003_ ), .ZN(_06991_ ) );
OR3_X1 _27821_ ( .A1(_06985_ ), .A2(_06989_ ), .A3(_06991_ ), .ZN(_06992_ ) );
NOR2_X1 _27822_ ( .A1(_06677_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06993_ ) );
OAI21_X1 _27823_ ( .A(_06681_ ), .B1(_06687_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06994_ ) );
OR3_X1 _27824_ ( .A1(_06992_ ), .A2(_06993_ ), .A3(_06994_ ), .ZN(_06995_ ) );
NAND3_X1 _27825_ ( .A1(_06679_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06741_ ), .ZN(_06996_ ) );
AOI21_X1 _27826_ ( .A(_06963_ ), .B1(_06995_ ), .B2(_06996_ ), .ZN(_06997_ ) );
OR2_X1 _27827_ ( .A1(_06840_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06998_ ) );
OR3_X1 _27828_ ( .A1(_06844_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03836_ ), .ZN(_06999_ ) );
AND3_X1 _27829_ ( .A1(_06997_ ), .A2(_06998_ ), .A3(_06999_ ), .ZN(_07000_ ) );
BUF_X4 _27830_ ( .A(_06606_ ), .Z(_07001_ ) );
NAND4_X1 _27831_ ( .A1(_06722_ ), .A2(_06926_ ), .A3(_04537_ ), .A4(_07001_ ), .ZN(_07002_ ) );
NAND4_X1 _27832_ ( .A1(_06755_ ), .A2(_06926_ ), .A3(_04541_ ), .A4(_07001_ ), .ZN(_07003_ ) );
NAND3_X1 _27833_ ( .A1(_07000_ ), .A2(_07002_ ), .A3(_07003_ ), .ZN(_07004_ ) );
NOR3_X1 _27834_ ( .A1(_06855_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03838_ ), .ZN(_07005_ ) );
BUF_X4 _27835_ ( .A(_06804_ ), .Z(_07006_ ) );
BUF_X4 _27836_ ( .A(_03837_ ), .Z(_07007_ ) );
NOR3_X1 _27837_ ( .A1(_07006_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07007_ ), .ZN(_07008_ ) );
NOR3_X1 _27838_ ( .A1(_07004_ ), .A2(_07005_ ), .A3(_07008_ ), .ZN(_07009_ ) );
BUF_X4 _27839_ ( .A(_06727_ ), .Z(_07010_ ) );
BUF_X4 _27840_ ( .A(_06607_ ), .Z(_07011_ ) );
NAND4_X1 _27841_ ( .A1(_06947_ ), .A2(_07010_ ), .A3(_04554_ ), .A4(_07011_ ), .ZN(_07012_ ) );
OR2_X1 _27842_ ( .A1(_06940_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07013_ ) );
AND3_X1 _27843_ ( .A1(_07009_ ), .A2(_07012_ ), .A3(_07013_ ), .ZN(_07014_ ) );
OR2_X1 _27844_ ( .A1(_06944_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07015_ ) );
OR2_X1 _27845_ ( .A1(_06943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07016_ ) );
NAND3_X1 _27846_ ( .A1(_07014_ ), .A2(_07015_ ), .A3(_07016_ ), .ZN(_07017_ ) );
BUF_X2 _27847_ ( .A(_06885_ ), .Z(_07018_ ) );
AND4_X1 _27848_ ( .A1(_04563_ ), .A2(_06936_ ), .A3(_06758_ ), .A4(_07018_ ), .ZN(_07019_ ) );
OAI21_X1 _27849_ ( .A(_06600_ ), .B1(_06872_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07020_ ) );
NOR3_X1 _27850_ ( .A1(_07017_ ), .A2(_07019_ ), .A3(_07020_ ), .ZN(_07021_ ) );
NAND3_X1 _27851_ ( .A1(_06761_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(\idu.immI [4] ), .ZN(_07022_ ) );
NAND4_X1 _27852_ ( .A1(_06956_ ), .A2(_06957_ ), .A3(_06877_ ), .A4(_07022_ ), .ZN(_07023_ ) );
OAI211_X1 _27853_ ( .A(_06960_ ), .B(_06962_ ), .C1(_07021_ ), .C2(_07023_ ), .ZN(\idu.io_out_bits_rs2_data [20] ) );
OAI21_X1 _27854_ ( .A(_06767_ ), .B1(_02100_ ), .B2(_02101_ ), .ZN(_07024_ ) );
AND4_X1 _27855_ ( .A1(\wbu.io_in_bits_rd_wdata [19] ), .A2(_06771_ ), .A3(_06773_ ), .A4(_06780_ ), .ZN(_07025_ ) );
AOI21_X1 _27856_ ( .A(_07025_ ), .B1(\lsu.io_out_bits_rd_wdata [19] ), .B2(_06784_ ), .ZN(_07026_ ) );
NAND4_X1 _27857_ ( .A1(_06708_ ), .A2(_06835_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_01099_ ), .ZN(_07027_ ) );
OR3_X1 _27858_ ( .A1(_06990_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06593_ ), .ZN(_07028_ ) );
OR3_X1 _27859_ ( .A1(_06640_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10812_ ), .ZN(_07029_ ) );
OR3_X1 _27860_ ( .A1(_11126_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10620_ ), .ZN(_07030_ ) );
OAI21_X1 _27861_ ( .A(_07030_ ), .B1(_06790_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_07031_ ) );
NOR2_X1 _27862_ ( .A1(_06620_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07032_ ) );
AND4_X1 _27863_ ( .A1(_04584_ ), .A2(_06622_ ), .A3(_10618_ ), .A4(_11049_ ), .ZN(_07033_ ) );
OR3_X1 _27864_ ( .A1(_07031_ ), .A2(_07032_ ), .A3(_07033_ ), .ZN(_07034_ ) );
NOR2_X1 _27865_ ( .A1(_06971_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07035_ ) );
AND2_X1 _27866_ ( .A1(_06635_ ), .A2(_11049_ ), .ZN(_07036_ ) );
INV_X1 _27867_ ( .A(_07036_ ), .ZN(_07037_ ) );
OAI21_X1 _27868_ ( .A(_07037_ ), .B1(_06633_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07038_ ) );
NOR3_X1 _27869_ ( .A1(_07034_ ), .A2(_07035_ ), .A3(_07038_ ), .ZN(_07039_ ) );
AND3_X1 _27870_ ( .A1(_06635_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11051_ ), .ZN(_07040_ ) );
OAI21_X1 _27871_ ( .A(_07029_ ), .B1(_07039_ ), .B2(_07040_ ), .ZN(_07041_ ) );
AND3_X1 _27872_ ( .A1(_06644_ ), .A2(_04595_ ), .A3(_06673_ ), .ZN(_07042_ ) );
AND4_X1 _27873_ ( .A1(_04597_ ), .A2(_10685_ ), .A3(_06601_ ), .A4(_06673_ ), .ZN(_07043_ ) );
OR3_X1 _27874_ ( .A1(_07041_ ), .A2(_07042_ ), .A3(_07043_ ), .ZN(_07044_ ) );
NOR2_X1 _27875_ ( .A1(_06650_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07045_ ) );
OAI21_X1 _27876_ ( .A(_06987_ ), .B1(_06660_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07046_ ) );
NOR3_X1 _27877_ ( .A1(_07044_ ), .A2(_07045_ ), .A3(_07046_ ), .ZN(_07047_ ) );
AND3_X1 _27878_ ( .A1(_06749_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06815_ ), .ZN(_07048_ ) );
OAI21_X1 _27879_ ( .A(_07028_ ), .B1(_07047_ ), .B2(_07048_ ), .ZN(_07049_ ) );
AND3_X1 _27880_ ( .A1(_06590_ ), .A2(_04579_ ), .A3(_06787_ ), .ZN(_07050_ ) );
NOR2_X1 _27881_ ( .A1(_06686_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07051_ ) );
OR3_X1 _27882_ ( .A1(_07049_ ), .A2(_07050_ ), .A3(_07051_ ), .ZN(_07052_ ) );
NOR3_X1 _27883_ ( .A1(_06829_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06846_ ), .ZN(_07053_ ) );
OR2_X1 _27884_ ( .A1(_07052_ ), .A2(_07053_ ), .ZN(_07054_ ) );
AND2_X2 _27885_ ( .A1(_06966_ ), .A2(_06594_ ), .ZN(_07055_ ) );
OAI21_X1 _27886_ ( .A(_07027_ ), .B1(_07054_ ), .B2(_07055_ ), .ZN(_07056_ ) );
BUF_X2 _27887_ ( .A(_06898_ ), .Z(_07057_ ) );
BUF_X2 _27888_ ( .A(_07057_ ), .Z(_07058_ ) );
NAND4_X1 _27889_ ( .A1(_07058_ ), .A2(_06916_ ), .A3(_04574_ ), .A4(_06750_ ), .ZN(_07059_ ) );
OR3_X1 _27890_ ( .A1(_06843_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03836_ ), .ZN(_07060_ ) );
AND3_X1 _27891_ ( .A1(_07056_ ), .A2(_07059_ ), .A3(_07060_ ), .ZN(_07061_ ) );
OR2_X1 _27892_ ( .A1(_06706_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07062_ ) );
NAND4_X1 _27893_ ( .A1(_06755_ ), .A2(_06926_ ), .A3(_04616_ ), .A4(_07001_ ), .ZN(_07063_ ) );
NAND3_X1 _27894_ ( .A1(_07061_ ), .A2(_07062_ ), .A3(_07063_ ), .ZN(_07064_ ) );
NOR3_X1 _27895_ ( .A1(_06855_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03838_ ), .ZN(_07065_ ) );
BUF_X2 _27896_ ( .A(_06699_ ), .Z(_07066_ ) );
CLKBUF_X2 _27897_ ( .A(_07066_ ), .Z(_07067_ ) );
AND4_X1 _27898_ ( .A1(_04622_ ), .A2(_06727_ ), .A3(_07067_ ), .A4(_06597_ ), .ZN(_07068_ ) );
NOR3_X1 _27899_ ( .A1(_07064_ ), .A2(_07065_ ), .A3(_07068_ ), .ZN(_07069_ ) );
NAND4_X1 _27900_ ( .A1(_06947_ ), .A2(_07010_ ), .A3(_04626_ ), .A4(_07011_ ), .ZN(_07070_ ) );
BUF_X4 _27901_ ( .A(_06727_ ), .Z(_07071_ ) );
NAND4_X1 _27902_ ( .A1(_06756_ ), .A2(_07071_ ), .A3(_04629_ ), .A4(_07011_ ), .ZN(_07072_ ) );
AND3_X1 _27903_ ( .A1(_07069_ ), .A2(_07070_ ), .A3(_07072_ ), .ZN(_07073_ ) );
OR2_X1 _27904_ ( .A1(_06944_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07074_ ) );
NAND4_X1 _27905_ ( .A1(_06949_ ), .A2(_07067_ ), .A3(_04634_ ), .A4(_07018_ ), .ZN(_07075_ ) );
NAND3_X1 _27906_ ( .A1(_07073_ ), .A2(_07074_ ), .A3(_07075_ ), .ZN(_07076_ ) );
NOR2_X1 _27907_ ( .A1(_06870_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07077_ ) );
OAI21_X1 _27908_ ( .A(_06600_ ), .B1(_06872_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07078_ ) );
NOR3_X1 _27909_ ( .A1(_07076_ ), .A2(_07077_ ), .A3(_07078_ ), .ZN(_07079_ ) );
BUF_X4 _27910_ ( .A(_01102_ ), .Z(_07080_ ) );
NAND3_X1 _27911_ ( .A1(_06761_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_07080_ ), .ZN(_07081_ ) );
NAND4_X1 _27912_ ( .A1(_06956_ ), .A2(_06957_ ), .A3(_06877_ ), .A4(_07081_ ), .ZN(_07082_ ) );
OAI211_X1 _27913_ ( .A(_07024_ ), .B(_07026_ ), .C1(_07079_ ), .C2(_07082_ ), .ZN(\idu.io_out_bits_rs2_data [19] ) );
OAI21_X1 _27914_ ( .A(_06560_ ), .B1(_02179_ ), .B2(_02180_ ), .ZN(_07083_ ) );
INV_X1 _27915_ ( .A(_06581_ ), .ZN(_07084_ ) );
AND4_X1 _27916_ ( .A1(\wbu.io_in_bits_rd_wdata [18] ), .A2(_07084_ ), .A3(_03990_ ), .A4(_06576_ ), .ZN(_07085_ ) );
AOI21_X1 _27917_ ( .A(_07085_ ), .B1(\lsu.io_out_bits_rd_wdata [18] ), .B2(_06581_ ), .ZN(_07086_ ) );
NAND3_X1 _27918_ ( .A1(_06761_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(\idu.immI [4] ), .ZN(_07087_ ) );
NAND3_X1 _27919_ ( .A1(_06858_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06728_ ), .ZN(_07088_ ) );
OR2_X1 _27920_ ( .A1(_06840_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07089_ ) );
NAND4_X1 _27921_ ( .A1(_06669_ ), .A2(_06724_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_06787_ ), .ZN(_07090_ ) );
OR2_X1 _27922_ ( .A1(_06646_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07091_ ) );
OR3_X1 _27923_ ( .A1(_06828_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10783_ ), .ZN(_07092_ ) );
OAI21_X1 _27924_ ( .A(_07092_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_10688_ ), .ZN(_07093_ ) );
BUF_X4 _27925_ ( .A(_06620_ ), .Z(_07094_ ) );
MUX2_X1 _27926_ ( .A(_04688_ ), .B(_07093_ ), .S(_07094_ ), .Z(_07095_ ) );
NOR3_X1 _27927_ ( .A1(_06794_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11122_ ), .ZN(_07096_ ) );
NOR2_X1 _27928_ ( .A1(_06972_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07097_ ) );
NOR3_X1 _27929_ ( .A1(_07095_ ), .A2(_07096_ ), .A3(_07097_ ), .ZN(_07098_ ) );
NAND4_X1 _27930_ ( .A1(_06668_ ), .A2(_06696_ ), .A3(_04692_ ), .A4(_06796_ ), .ZN(_07099_ ) );
AOI22_X1 _27931_ ( .A1(_07036_ ), .A2(_04694_ ), .B1(_06796_ ), .B2(_06603_ ), .ZN(_07100_ ) );
AND3_X1 _27932_ ( .A1(_07098_ ), .A2(_07099_ ), .A3(_07100_ ), .ZN(_07101_ ) );
AND3_X1 _27933_ ( .A1(_06603_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06609_ ), .ZN(_07102_ ) );
OAI21_X1 _27934_ ( .A(_07091_ ), .B1(_07101_ ), .B2(_07102_ ), .ZN(_07103_ ) );
OAI21_X1 _27935_ ( .A(_07090_ ), .B1(_07103_ ), .B2(_06654_ ), .ZN(_07104_ ) );
NAND4_X1 _27936_ ( .A1(_06898_ ), .A2(_06724_ ), .A3(_04683_ ), .A4(_06816_ ), .ZN(_07105_ ) );
BUF_X2 _27937_ ( .A(_06660_ ), .Z(_07106_ ) );
OR2_X1 _27938_ ( .A1(_07106_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07107_ ) );
NAND3_X1 _27939_ ( .A1(_07104_ ), .A2(_07105_ ), .A3(_07107_ ), .ZN(_07108_ ) );
NOR2_X1 _27940_ ( .A1(_06988_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07109_ ) );
BUF_X2 _27941_ ( .A(_06990_ ), .Z(_07110_ ) );
NOR3_X1 _27942_ ( .A1(_07110_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06594_ ), .ZN(_07111_ ) );
NOR3_X1 _27943_ ( .A1(_07108_ ), .A2(_07109_ ), .A3(_07111_ ), .ZN(_07112_ ) );
OR2_X1 _27944_ ( .A1(_06676_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07113_ ) );
OR2_X1 _27945_ ( .A1(_06687_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07114_ ) );
NAND3_X1 _27946_ ( .A1(_07112_ ), .A2(_07113_ ), .A3(_07114_ ), .ZN(_07115_ ) );
NOR3_X1 _27947_ ( .A1(_06829_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06612_ ), .ZN(_07116_ ) );
NOR3_X1 _27948_ ( .A1(_07115_ ), .A2(_07055_ ), .A3(_07116_ ), .ZN(_07117_ ) );
AND3_X1 _27949_ ( .A1(_06966_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06605_ ), .ZN(_07118_ ) );
OAI21_X1 _27950_ ( .A(_07089_ ), .B1(_07117_ ), .B2(_07118_ ), .ZN(_07119_ ) );
AND3_X1 _27951_ ( .A1(_06623_ ), .A2(_04715_ ), .A3(_06596_ ), .ZN(_07120_ ) );
AND4_X1 _27952_ ( .A1(_04717_ ), .A2(_06721_ ), .A3(_06698_ ), .A4(_01099_ ), .ZN(_07121_ ) );
NOR3_X1 _27953_ ( .A1(_07119_ ), .A2(_07120_ ), .A3(_07121_ ), .ZN(_07122_ ) );
OR2_X1 _27954_ ( .A1(_06930_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07123_ ) );
NAND4_X1 _27955_ ( .A1(_07058_ ), .A2(_06711_ ), .A3(_04721_ ), .A4(_06597_ ), .ZN(_07124_ ) );
NAND3_X1 _27956_ ( .A1(_07122_ ), .A2(_07123_ ), .A3(_07124_ ), .ZN(_07125_ ) );
OAI21_X1 _27957_ ( .A(_06860_ ), .B1(_06933_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07126_ ) );
OAI21_X1 _27958_ ( .A(_07088_ ), .B1(_07125_ ), .B2(_07126_ ), .ZN(_07127_ ) );
NAND4_X1 _27959_ ( .A1(_06756_ ), .A2(_07071_ ), .A3(_04727_ ), .A4(_06866_ ), .ZN(_07128_ ) );
OR2_X1 _27960_ ( .A1(_06737_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07129_ ) );
AND3_X1 _27961_ ( .A1(_07127_ ), .A2(_07128_ ), .A3(_07129_ ), .ZN(_07130_ ) );
OR2_X1 _27962_ ( .A1(_06743_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07131_ ) );
NAND4_X1 _27963_ ( .A1(_06948_ ), .A2(_06758_ ), .A3(_04733_ ), .A4(_06883_ ), .ZN(_07132_ ) );
NAND3_X1 _27964_ ( .A1(_07130_ ), .A2(_07131_ ), .A3(_07132_ ), .ZN(_07133_ ) );
BUF_X4 _27965_ ( .A(_06599_ ), .Z(_07134_ ) );
OAI21_X1 _27966_ ( .A(_07134_ ), .B1(_06872_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07135_ ) );
OAI21_X1 _27967_ ( .A(_07087_ ), .B1(_07133_ ), .B2(_07135_ ), .ZN(_07136_ ) );
OAI221_X1 _27968_ ( .A(_07083_ ), .B1(_06560_ ), .B2(_07086_ ), .C1(_06584_ ), .C2(_07136_ ), .ZN(\idu.io_out_bits_rs2_data [18] ) );
OAI21_X1 _27969_ ( .A(_06767_ ), .B1(_02252_ ), .B2(_02253_ ), .ZN(_07137_ ) );
CLKBUF_X2 _27970_ ( .A(_06772_ ), .Z(_07138_ ) );
AND4_X1 _27971_ ( .A1(\wbu.io_in_bits_rd_wdata [17] ), .A2(_06771_ ), .A3(_07138_ ), .A4(_06780_ ), .ZN(_07139_ ) );
AOI21_X1 _27972_ ( .A(_07139_ ), .B1(\lsu.io_out_bits_rd_wdata [17] ), .B2(_06784_ ), .ZN(_07140_ ) );
OR2_X1 _27973_ ( .A1(_06752_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07141_ ) );
OR2_X1 _27974_ ( .A1(_06840_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07142_ ) );
NAND3_X1 _27975_ ( .A1(_06603_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06609_ ), .ZN(_07143_ ) );
NOR3_X1 _27976_ ( .A1(_06828_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_11121_ ), .ZN(_07144_ ) );
AOI21_X1 _27977_ ( .A(_07144_ ), .B1(_04772_ ), .B2(_10687_ ), .ZN(_07145_ ) );
NAND4_X1 _27978_ ( .A1(_06586_ ), .A2(_06682_ ), .A3(_04774_ ), .A4(_11051_ ), .ZN(_07146_ ) );
OR3_X1 _27979_ ( .A1(_06625_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11121_ ), .ZN(_07147_ ) );
AND3_X1 _27980_ ( .A1(_07145_ ), .A2(_07146_ ), .A3(_07147_ ), .ZN(_07148_ ) );
OR2_X1 _27981_ ( .A1(_06972_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07149_ ) );
NAND4_X1 _27982_ ( .A1(_06668_ ), .A2(_06696_ ), .A3(_04778_ ), .A4(_11052_ ), .ZN(_07150_ ) );
NAND3_X1 _27983_ ( .A1(_07148_ ), .A2(_07149_ ), .A3(_07150_ ), .ZN(_07151_ ) );
AND2_X1 _27984_ ( .A1(_06603_ ), .A2(_11051_ ), .ZN(_07152_ ) );
INV_X1 _27985_ ( .A(_07152_ ), .ZN(_07153_ ) );
OAI21_X1 _27986_ ( .A(_07153_ ), .B1(_07037_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07154_ ) );
OAI21_X1 _27987_ ( .A(_07143_ ), .B1(_07151_ ), .B2(_07154_ ), .ZN(_07155_ ) );
BUF_X2 _27988_ ( .A(_06601_ ), .Z(_07156_ ) );
NAND4_X1 _27989_ ( .A1(_06663_ ), .A2(_07156_ ), .A3(_04783_ ), .A4(_03833_ ), .ZN(_07157_ ) );
OR2_X1 _27990_ ( .A1(_06655_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07158_ ) );
NAND3_X1 _27991_ ( .A1(_07155_ ), .A2(_07157_ ), .A3(_07158_ ), .ZN(_07159_ ) );
NOR2_X1 _27992_ ( .A1(_06651_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07160_ ) );
NOR3_X1 _27993_ ( .A1(_07159_ ), .A2(_06659_ ), .A3(_07160_ ), .ZN(_07161_ ) );
AND3_X1 _27994_ ( .A1(_06658_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06787_ ), .ZN(_07162_ ) );
NOR2_X1 _27995_ ( .A1(_07161_ ), .A2(_07162_ ), .ZN(_07163_ ) );
NOR2_X1 _27996_ ( .A1(_06988_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07164_ ) );
NOR3_X1 _27997_ ( .A1(_07110_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06594_ ), .ZN(_07165_ ) );
NOR3_X1 _27998_ ( .A1(_07163_ ), .A2(_07164_ ), .A3(_07165_ ), .ZN(_07166_ ) );
NAND4_X1 _27999_ ( .A1(_07057_ ), .A2(_06666_ ), .A3(_04793_ ), .A4(_06817_ ), .ZN(_07167_ ) );
OR2_X1 _28000_ ( .A1(_06686_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07168_ ) );
NAND3_X1 _28001_ ( .A1(_07166_ ), .A2(_07167_ ), .A3(_07168_ ), .ZN(_07169_ ) );
NOR3_X1 _28002_ ( .A1(_06829_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06846_ ), .ZN(_07170_ ) );
NOR3_X1 _28003_ ( .A1(_07169_ ), .A2(_07055_ ), .A3(_07170_ ), .ZN(_07171_ ) );
AND3_X1 _28004_ ( .A1(_06966_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06691_ ), .ZN(_07172_ ) );
OAI21_X1 _28005_ ( .A(_07142_ ), .B1(_07171_ ), .B2(_07172_ ), .ZN(_07173_ ) );
AND3_X1 _28006_ ( .A1(_06623_ ), .A2(_04801_ ), .A3(_06741_ ), .ZN(_07174_ ) );
AND4_X1 _28007_ ( .A1(_04804_ ), .A2(_06907_ ), .A3(_06698_ ), .A4(_06605_ ), .ZN(_07175_ ) );
NOR3_X1 _28008_ ( .A1(_07173_ ), .A2(_07174_ ), .A3(_07175_ ), .ZN(_07176_ ) );
OR2_X1 _28009_ ( .A1(_06930_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07177_ ) );
NAND4_X1 _28010_ ( .A1(_07058_ ), .A2(_06711_ ), .A3(_04808_ ), .A4(_06852_ ), .ZN(_07178_ ) );
NAND3_X1 _28011_ ( .A1(_07176_ ), .A2(_07177_ ), .A3(_07178_ ), .ZN(_07179_ ) );
NOR3_X1 _28012_ ( .A1(_07006_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06856_ ), .ZN(_07180_ ) );
AND4_X1 _28013_ ( .A1(_04812_ ), .A2(_06721_ ), .A3(_06726_ ), .A4(_01100_ ), .ZN(_07181_ ) );
OR3_X1 _28014_ ( .A1(_07179_ ), .A2(_07180_ ), .A3(_07181_ ), .ZN(_07182_ ) );
NOR2_X1 _28015_ ( .A1(_06940_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07183_ ) );
OAI21_X1 _28016_ ( .A(_06743_ ), .B1(_06738_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07184_ ) );
NOR3_X1 _28017_ ( .A1(_07182_ ), .A2(_07183_ ), .A3(_07184_ ), .ZN(_07185_ ) );
AND3_X1 _28018_ ( .A1(_06740_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01102_ ), .ZN(_07186_ ) );
OAI21_X1 _28019_ ( .A(_07141_ ), .B1(_07185_ ), .B2(_07186_ ), .ZN(_07187_ ) );
BUF_X2 _28020_ ( .A(_07110_ ), .Z(_07188_ ) );
NOR3_X1 _28021_ ( .A1(_07188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03838_ ), .ZN(_07189_ ) );
NOR3_X1 _28022_ ( .A1(_07187_ ), .A2(_06598_ ), .A3(_07189_ ), .ZN(_07190_ ) );
OAI211_X1 _28023_ ( .A(_06875_ ), .B(_06877_ ), .C1(_04824_ ), .C2(_06600_ ), .ZN(_07191_ ) );
OAI211_X1 _28024_ ( .A(_07137_ ), .B(_07140_ ), .C1(_07190_ ), .C2(_07191_ ), .ZN(\idu.io_out_bits_rs2_data [17] ) );
AND3_X1 _28025_ ( .A1(_02326_ ), .A2(_02327_ ), .A3(_06767_ ), .ZN(_07192_ ) );
INV_X1 _28026_ ( .A(_06783_ ), .ZN(_07193_ ) );
INV_X1 _28027_ ( .A(_06875_ ), .ZN(_07194_ ) );
BUF_X4 _28028_ ( .A(_03989_ ), .Z(_07195_ ) );
BUF_X4 _28029_ ( .A(_06778_ ), .Z(_07196_ ) );
NOR3_X1 _28030_ ( .A1(_07195_ ), .A2(_13518_ ), .A3(_07196_ ), .ZN(_07197_ ) );
OAI22_X1 _28031_ ( .A1(\lsu.io_out_bits_rd_wdata [16] ), .A2(_07193_ ), .B1(_07194_ ), .B2(_07197_ ), .ZN(_07198_ ) );
CLKBUF_X2 _28032_ ( .A(_06611_ ), .Z(_07199_ ) );
OR3_X1 _28033_ ( .A1(_06918_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07199_ ), .ZN(_07200_ ) );
AND4_X1 _28034_ ( .A1(_04870_ ), .A2(_06669_ ), .A3(_06909_ ), .A4(_06816_ ), .ZN(_07201_ ) );
NAND3_X1 _28035_ ( .A1(_06966_ ), .A2(_04850_ ), .A3(_06653_ ), .ZN(_07202_ ) );
OAI21_X1 _28036_ ( .A(_07202_ ), .B1(_06791_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_07203_ ) );
AOI211_X1 _28037_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_06625_ ), .C1(\idu.io_in_bits_inst [24] ), .C2(_10646_ ), .ZN(_07204_ ) );
NOR2_X1 _28038_ ( .A1(_07094_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07205_ ) );
NOR3_X1 _28039_ ( .A1(_07203_ ), .A2(_07204_ ), .A3(_07205_ ), .ZN(_07206_ ) );
OR2_X1 _28040_ ( .A1(_06971_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07207_ ) );
NAND3_X1 _28041_ ( .A1(_06631_ ), .A2(_04856_ ), .A3(_03832_ ), .ZN(_07208_ ) );
AND3_X1 _28042_ ( .A1(_07206_ ), .A2(_07207_ ), .A3(_07208_ ), .ZN(_07209_ ) );
BUF_X2 _28043_ ( .A(_06628_ ), .Z(_07210_ ) );
NAND4_X1 _28044_ ( .A1(_06897_ ), .A2(_07210_ ), .A3(_04859_ ), .A4(_06674_ ), .ZN(_07211_ ) );
OR3_X1 _28045_ ( .A1(_06640_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06592_ ), .ZN(_07212_ ) );
AND3_X1 _28046_ ( .A1(_07209_ ), .A2(_07211_ ), .A3(_07212_ ), .ZN(_07213_ ) );
OR2_X1 _28047_ ( .A1(_06647_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07214_ ) );
BUF_X2 _28048_ ( .A(_06668_ ), .Z(_07215_ ) );
NAND4_X1 _28049_ ( .A1(_07215_ ), .A2(_07156_ ), .A3(_04846_ ), .A4(_06815_ ), .ZN(_07216_ ) );
NAND3_X1 _28050_ ( .A1(_07213_ ), .A2(_07214_ ), .A3(_07216_ ), .ZN(_07217_ ) );
NOR2_X1 _28051_ ( .A1(_06651_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07218_ ) );
OAI21_X1 _28052_ ( .A(_06988_ ), .B1(_07106_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07219_ ) );
OR3_X1 _28053_ ( .A1(_07217_ ), .A2(_07218_ ), .A3(_07219_ ), .ZN(_07220_ ) );
NAND3_X1 _28054_ ( .A1(_06749_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06817_ ), .ZN(_07221_ ) );
AOI21_X1 _28055_ ( .A(_07201_ ), .B1(_07220_ ), .B2(_07221_ ), .ZN(_07222_ ) );
OR2_X1 _28056_ ( .A1(_06677_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07223_ ) );
NOR2_X1 _28057_ ( .A1(_06687_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07224_ ) );
NOR2_X1 _28058_ ( .A1(_07224_ ), .A2(_06680_ ), .ZN(_07225_ ) );
AND3_X1 _28059_ ( .A1(_07222_ ), .A2(_07223_ ), .A3(_07225_ ), .ZN(_07226_ ) );
AND3_X1 _28060_ ( .A1(_06679_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06605_ ), .ZN(_07227_ ) );
OAI21_X1 _28061_ ( .A(_07200_ ), .B1(_07226_ ), .B2(_07227_ ), .ZN(_07228_ ) );
NOR2_X1 _28062_ ( .A1(_06841_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07229_ ) );
AND4_X1 _28063_ ( .A1(_04879_ ), .A2(_06698_ ), .A3(_06699_ ), .A4(_06741_ ), .ZN(_07230_ ) );
NOR3_X1 _28064_ ( .A1(_07228_ ), .A2(_07229_ ), .A3(_07230_ ), .ZN(_07231_ ) );
BUF_X4 _28065_ ( .A(_06710_ ), .Z(_07232_ ) );
NAND4_X1 _28066_ ( .A1(_06850_ ), .A2(_07232_ ), .A3(_04881_ ), .A4(_06865_ ), .ZN(_07233_ ) );
OR2_X1 _28067_ ( .A1(_06930_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07234_ ) );
NAND3_X1 _28068_ ( .A1(_07231_ ), .A2(_07233_ ), .A3(_07234_ ), .ZN(_07235_ ) );
NOR3_X1 _28069_ ( .A1(_06855_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06856_ ), .ZN(_07236_ ) );
AND4_X1 _28070_ ( .A1(_04887_ ), .A2(_06726_ ), .A3(_07066_ ), .A4(_06852_ ), .ZN(_07237_ ) );
NOR3_X1 _28071_ ( .A1(_07235_ ), .A2(_07236_ ), .A3(_07237_ ), .ZN(_07238_ ) );
NAND4_X1 _28072_ ( .A1(_06947_ ), .A2(_07071_ ), .A3(_04889_ ), .A4(_06866_ ), .ZN(_07239_ ) );
OR2_X1 _28073_ ( .A1(_06940_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07240_ ) );
AND3_X1 _28074_ ( .A1(_07238_ ), .A2(_07239_ ), .A3(_07240_ ), .ZN(_07241_ ) );
NAND4_X1 _28075_ ( .A1(_07058_ ), .A2(_06937_ ), .A3(_04893_ ), .A4(_07018_ ), .ZN(_07242_ ) );
OR2_X1 _28076_ ( .A1(_06743_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07243_ ) );
NAND3_X1 _28077_ ( .A1(_07241_ ), .A2(_07242_ ), .A3(_07243_ ), .ZN(_07244_ ) );
NOR2_X1 _28078_ ( .A1(_06870_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07245_ ) );
OAI21_X1 _28079_ ( .A(_07134_ ), .B1(_06748_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07246_ ) );
NOR3_X1 _28080_ ( .A1(_07244_ ), .A2(_07245_ ), .A3(_07246_ ), .ZN(_07247_ ) );
BUF_X4 _28081_ ( .A(_06771_ ), .Z(_07248_ ) );
BUF_X4 _28082_ ( .A(_06773_ ), .Z(_07249_ ) );
BUF_X4 _28083_ ( .A(_06876_ ), .Z(_07250_ ) );
BUF_X4 _28084_ ( .A(_06591_ ), .Z(_07251_ ) );
NAND3_X1 _28085_ ( .A1(_07251_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_06950_ ), .ZN(_07252_ ) );
NAND4_X1 _28086_ ( .A1(_07248_ ), .A2(_07249_ ), .A3(_07250_ ), .A4(_07252_ ), .ZN(_07253_ ) );
OAI22_X1 _28087_ ( .A1(_07192_ ), .A2(_07198_ ), .B1(_07247_ ), .B2(_07253_ ), .ZN(\idu.io_out_bits_rs2_data [16] ) );
NAND2_X1 _28088_ ( .A1(\exu.io_out_bits_rd_wdata [15] ), .A2(_06879_ ), .ZN(_07254_ ) );
AND4_X1 _28089_ ( .A1(\wbu.io_in_bits_rd_wdata [15] ), .A2(_06771_ ), .A3(_07138_ ), .A4(_06780_ ), .ZN(_07255_ ) );
AOI21_X1 _28090_ ( .A(_07255_ ), .B1(\lsu.io_out_bits_rd_wdata [15] ), .B2(_06784_ ), .ZN(_07256_ ) );
NOR2_X1 _28091_ ( .A1(_06824_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07257_ ) );
CLKBUF_X2 _28092_ ( .A(_11052_ ), .Z(_07258_ ) );
AND3_X1 _28093_ ( .A1(_06603_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07258_ ), .ZN(_07259_ ) );
OR3_X1 _28094_ ( .A1(_06827_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10620_ ), .ZN(_07260_ ) );
MUX2_X1 _28095_ ( .A(_07260_ ), .B(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(_10687_ ), .Z(_07261_ ) );
MUX2_X1 _28096_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_07261_ ), .S(_07094_ ), .Z(_07262_ ) );
AND2_X1 _28097_ ( .A1(_06623_ ), .A2(_11049_ ), .ZN(_07263_ ) );
INV_X1 _28098_ ( .A(_07263_ ), .ZN(_07264_ ) );
MUX2_X1 _28099_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_07262_ ), .S(_07264_ ), .Z(_07265_ ) );
NAND4_X1 _28100_ ( .A1(_06663_ ), .A2(_07210_ ), .A3(_04922_ ), .A4(_06609_ ), .ZN(_07266_ ) );
OR2_X1 _28101_ ( .A1(_06799_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07267_ ) );
AND3_X1 _28102_ ( .A1(_07265_ ), .A2(_07266_ ), .A3(_07267_ ), .ZN(_07268_ ) );
NOR3_X1 _28103_ ( .A1(_06637_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06593_ ), .ZN(_07269_ ) );
NOR2_X1 _28104_ ( .A1(_07269_ ), .A2(_07152_ ), .ZN(_07270_ ) );
AOI21_X1 _28105_ ( .A(_07259_ ), .B1(_07268_ ), .B2(_07270_ ), .ZN(_07271_ ) );
NOR2_X1 _28106_ ( .A1(_06647_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07272_ ) );
AND3_X1 _28107_ ( .A1(_06730_ ), .A2(_04930_ ), .A3(_06787_ ), .ZN(_07273_ ) );
NOR3_X1 _28108_ ( .A1(_07271_ ), .A2(_07272_ ), .A3(_07273_ ), .ZN(_07274_ ) );
NAND4_X1 _28109_ ( .A1(_06898_ ), .A2(_06725_ ), .A3(_04932_ ), .A4(_06611_ ), .ZN(_07275_ ) );
OR2_X1 _28110_ ( .A1(_06661_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07276_ ) );
AND3_X1 _28111_ ( .A1(_07274_ ), .A2(_07275_ ), .A3(_07276_ ), .ZN(_07277_ ) );
NAND4_X1 _28112_ ( .A1(_06907_ ), .A2(_06757_ ), .A3(_04937_ ), .A4(_06831_ ), .ZN(_07278_ ) );
AOI22_X1 _28113_ ( .A1(_06819_ ), .A2(_04940_ ), .B1(_06612_ ), .B2(_06590_ ), .ZN(_07279_ ) );
NAND3_X1 _28114_ ( .A1(_07277_ ), .A2(_07278_ ), .A3(_07279_ ), .ZN(_07280_ ) );
NAND3_X1 _28115_ ( .A1(_06591_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03836_ ), .ZN(_07281_ ) );
AOI21_X1 _28116_ ( .A(_07257_ ), .B1(_07280_ ), .B2(_07281_ ), .ZN(_07282_ ) );
OR3_X1 _28117_ ( .A1(_06830_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06919_ ), .ZN(_07283_ ) );
OR3_X1 _28118_ ( .A1(_06918_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07199_ ), .ZN(_07284_ ) );
NAND3_X1 _28119_ ( .A1(_07282_ ), .A2(_07283_ ), .A3(_07284_ ), .ZN(_07285_ ) );
NOR2_X1 _28120_ ( .A1(_06841_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07286_ ) );
NOR3_X1 _28121_ ( .A1(_06844_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03837_ ), .ZN(_07287_ ) );
NOR3_X1 _28122_ ( .A1(_07285_ ), .A2(_07286_ ), .A3(_07287_ ), .ZN(_07288_ ) );
NAND4_X1 _28123_ ( .A1(_06850_ ), .A2(_06926_ ), .A3(_04954_ ), .A4(_07001_ ), .ZN(_07289_ ) );
NAND4_X1 _28124_ ( .A1(_06755_ ), .A2(_07232_ ), .A3(_04956_ ), .A4(_07001_ ), .ZN(_07290_ ) );
NAND3_X1 _28125_ ( .A1(_07288_ ), .A2(_07289_ ), .A3(_07290_ ), .ZN(_07291_ ) );
NOR3_X1 _28126_ ( .A1(_06855_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07007_ ), .ZN(_07292_ ) );
NOR3_X1 _28127_ ( .A1(_07006_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07007_ ), .ZN(_07293_ ) );
NOR3_X1 _28128_ ( .A1(_07291_ ), .A2(_07292_ ), .A3(_07293_ ), .ZN(_07294_ ) );
NAND4_X1 _28129_ ( .A1(_06936_ ), .A2(_06937_ ), .A3(_04962_ ), .A4(_06938_ ), .ZN(_07295_ ) );
NAND4_X1 _28130_ ( .A1(_06756_ ), .A2(_07010_ ), .A3(_04964_ ), .A4(_07011_ ), .ZN(_07296_ ) );
NAND3_X1 _28131_ ( .A1(_07294_ ), .A2(_07295_ ), .A3(_07296_ ), .ZN(_07297_ ) );
NOR2_X1 _28132_ ( .A1(_06944_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07298_ ) );
NOR2_X1 _28133_ ( .A1(_06943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07299_ ) );
NOR3_X1 _28134_ ( .A1(_07297_ ), .A2(_07298_ ), .A3(_07299_ ), .ZN(_07300_ ) );
NAND4_X1 _28135_ ( .A1(_06948_ ), .A2(_06949_ ), .A3(_04969_ ), .A4(_06952_ ), .ZN(_07301_ ) );
AOI22_X1 _28136_ ( .A1(_06747_ ), .A2(_04971_ ), .B1(_06952_ ), .B2(_06953_ ), .ZN(_07302_ ) );
AND3_X1 _28137_ ( .A1(_07300_ ), .A2(_07301_ ), .A3(_07302_ ), .ZN(_07303_ ) );
NAND3_X1 _28138_ ( .A1(_06761_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_07080_ ), .ZN(_07304_ ) );
NAND4_X1 _28139_ ( .A1(_06956_ ), .A2(_06957_ ), .A3(_06877_ ), .A4(_07304_ ), .ZN(_07305_ ) );
OAI211_X1 _28140_ ( .A(_07254_ ), .B(_07256_ ), .C1(_07303_ ), .C2(_07305_ ), .ZN(\idu.io_out_bits_rs2_data [15] ) );
NAND2_X1 _28141_ ( .A1(\exu.io_out_bits_rd_wdata [14] ), .A2(_06560_ ), .ZN(_07306_ ) );
AOI211_X1 _28142_ ( .A(_13592_ ), .B(_06577_ ), .C1(_06579_ ), .C2(_10755_ ), .ZN(_07307_ ) );
AOI21_X1 _28143_ ( .A(_07307_ ), .B1(\lsu.io_out_bits_rd_wdata [14] ), .B2(_06581_ ), .ZN(_07308_ ) );
NAND3_X1 _28144_ ( .A1(_06761_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(\idu.immI [4] ), .ZN(_07309_ ) );
NAND4_X1 _28145_ ( .A1(_06721_ ), .A2(_06710_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_06606_ ), .ZN(_07310_ ) );
OR3_X1 _28146_ ( .A1(_06843_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07199_ ), .ZN(_07311_ ) );
OR3_X1 _28147_ ( .A1(_06990_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11124_ ), .ZN(_07312_ ) );
NAND4_X1 _28148_ ( .A1(_07215_ ), .A2(_07156_ ), .A3(_05014_ ), .A4(_06815_ ), .ZN(_07313_ ) );
NAND3_X1 _28149_ ( .A1(_06618_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06653_ ), .ZN(_07314_ ) );
OR3_X1 _28150_ ( .A1(_06828_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10620_ ), .ZN(_07315_ ) );
OAI21_X1 _28151_ ( .A(_07315_ ), .B1(_10688_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07316_ ) );
OAI21_X1 _28152_ ( .A(_07314_ ), .B1(_07316_ ), .B2(_06619_ ), .ZN(_07317_ ) );
OAI21_X1 _28153_ ( .A(_07317_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_07264_ ), .ZN(_07318_ ) );
AND4_X1 _28154_ ( .A1(_04997_ ), .A2(_06627_ ), .A3(_06628_ ), .A4(_06653_ ), .ZN(_07319_ ) );
NOR2_X1 _28155_ ( .A1(_06633_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07320_ ) );
OR3_X1 _28156_ ( .A1(_07318_ ), .A2(_07319_ ), .A3(_07320_ ), .ZN(_07321_ ) );
AOI211_X1 _28157_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_06637_ ), .C1(\idu.io_in_bits_inst [24] ), .C2(_11030_ ), .ZN(_07322_ ) );
AND4_X1 _28158_ ( .A1(_05008_ ), .A2(_06601_ ), .A3(_06683_ ), .A4(_11051_ ), .ZN(_07323_ ) );
OR2_X1 _28159_ ( .A1(_06645_ ), .A2(_07323_ ), .ZN(_07324_ ) );
NOR3_X1 _28160_ ( .A1(_07321_ ), .A2(_07322_ ), .A3(_07324_ ), .ZN(_07325_ ) );
AND3_X1 _28161_ ( .A1(_06858_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03833_ ), .ZN(_07326_ ) );
OAI21_X1 _28162_ ( .A(_07313_ ), .B1(_07325_ ), .B2(_07326_ ), .ZN(_07327_ ) );
NOR2_X1 _28163_ ( .A1(_06651_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07328_ ) );
OAI21_X1 _28164_ ( .A(_06988_ ), .B1(_07106_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07329_ ) );
NOR3_X1 _28165_ ( .A1(_07327_ ), .A2(_07328_ ), .A3(_07329_ ), .ZN(_07330_ ) );
AND3_X1 _28166_ ( .A1(_06749_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06811_ ), .ZN(_07331_ ) );
OAI21_X1 _28167_ ( .A(_07312_ ), .B1(_07330_ ), .B2(_07331_ ), .ZN(_07332_ ) );
AND4_X1 _28168_ ( .A1(_05024_ ), .A2(_06898_ ), .A3(_06909_ ), .A4(_06816_ ), .ZN(_07333_ ) );
NOR2_X1 _28169_ ( .A1(_06687_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07334_ ) );
NOR3_X1 _28170_ ( .A1(_07332_ ), .A2(_07333_ ), .A3(_07334_ ), .ZN(_07335_ ) );
NAND4_X1 _28171_ ( .A1(_06720_ ), .A2(_06834_ ), .A3(_05028_ ), .A4(_06595_ ), .ZN(_07336_ ) );
AOI22_X1 _28172_ ( .A1(_07055_ ), .A2(_05030_ ), .B1(_11125_ ), .B2(_06694_ ), .ZN(_07337_ ) );
AND3_X1 _28173_ ( .A1(_07335_ ), .A2(_07336_ ), .A3(_07337_ ), .ZN(_07338_ ) );
AND3_X1 _28174_ ( .A1(_06694_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06605_ ), .ZN(_07339_ ) );
OAI21_X1 _28175_ ( .A(_07311_ ), .B1(_07338_ ), .B2(_07339_ ), .ZN(_07340_ ) );
OAI21_X1 _28176_ ( .A(_07310_ ), .B1(_07340_ ), .B2(_06704_ ), .ZN(_07341_ ) );
NAND4_X1 _28177_ ( .A1(_06709_ ), .A2(_07232_ ), .A3(_05036_ ), .A4(_06865_ ), .ZN(_07342_ ) );
OR3_X1 _28178_ ( .A1(_06802_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06847_ ), .ZN(_07343_ ) );
NAND3_X1 _28179_ ( .A1(_07341_ ), .A2(_07342_ ), .A3(_07343_ ), .ZN(_07344_ ) );
NOR3_X1 _28180_ ( .A1(_07006_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06856_ ), .ZN(_07345_ ) );
AND4_X1 _28181_ ( .A1(_05043_ ), .A2(_06850_ ), .A3(_06726_ ), .A4(_06852_ ), .ZN(_07346_ ) );
NOR3_X1 _28182_ ( .A1(_07344_ ), .A2(_07345_ ), .A3(_07346_ ), .ZN(_07347_ ) );
NAND4_X1 _28183_ ( .A1(_06755_ ), .A2(_07071_ ), .A3(_05046_ ), .A4(_06866_ ), .ZN(_07348_ ) );
OR2_X1 _28184_ ( .A1(_06737_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07349_ ) );
AND3_X1 _28185_ ( .A1(_07347_ ), .A2(_07348_ ), .A3(_07349_ ), .ZN(_07350_ ) );
OR2_X1 _28186_ ( .A1(_06743_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07351_ ) );
NAND4_X1 _28187_ ( .A1(_06948_ ), .A2(_06758_ ), .A3(_05051_ ), .A4(_06883_ ), .ZN(_07352_ ) );
NAND3_X1 _28188_ ( .A1(_07350_ ), .A2(_07351_ ), .A3(_07352_ ), .ZN(_07353_ ) );
OAI21_X1 _28189_ ( .A(_07134_ ), .B1(_06872_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07354_ ) );
OAI21_X1 _28190_ ( .A(_07309_ ), .B1(_07353_ ), .B2(_07354_ ), .ZN(_07355_ ) );
OAI221_X1 _28191_ ( .A(_07306_ ), .B1(_06560_ ), .B2(_07308_ ), .C1(_06584_ ), .C2(_07355_ ), .ZN(\idu.io_out_bits_rs2_data [14] ) );
NAND2_X1 _28192_ ( .A1(\exu.io_out_bits_rd_wdata [13] ), .A2(_06879_ ), .ZN(_07356_ ) );
AND4_X1 _28193_ ( .A1(\wbu.io_in_bits_rd_wdata [13] ), .A2(_06771_ ), .A3(_07138_ ), .A4(_06780_ ), .ZN(_07357_ ) );
AOI21_X1 _28194_ ( .A(_07357_ ), .B1(\lsu.io_out_bits_rd_wdata [13] ), .B2(_06784_ ), .ZN(_07358_ ) );
AND4_X1 _28195_ ( .A1(_05105_ ), .A2(_06710_ ), .A3(_07066_ ), .A4(_06596_ ), .ZN(_07359_ ) );
NAND3_X1 _28196_ ( .A1(_06740_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06817_ ), .ZN(_07360_ ) );
NAND3_X1 _28197_ ( .A1(_06603_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06811_ ), .ZN(_07361_ ) );
NAND3_X1 _28198_ ( .A1(_06966_ ), .A2(_05071_ ), .A3(_06674_ ), .ZN(_07362_ ) );
OAI21_X1 _28199_ ( .A(_07362_ ), .B1(_06791_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_07363_ ) );
AND4_X1 _28200_ ( .A1(_05075_ ), .A2(_06897_ ), .A3(_06833_ ), .A4(_06814_ ), .ZN(_07364_ ) );
NOR3_X1 _28201_ ( .A1(_06843_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11123_ ), .ZN(_07365_ ) );
NOR3_X1 _28202_ ( .A1(_07363_ ), .A2(_07364_ ), .A3(_07365_ ), .ZN(_07366_ ) );
OR2_X1 _28203_ ( .A1(_06972_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07367_ ) );
NAND4_X1 _28204_ ( .A1(_07215_ ), .A2(_06697_ ), .A3(_05069_ ), .A4(_06610_ ), .ZN(_07368_ ) );
NAND3_X1 _28205_ ( .A1(_07366_ ), .A2(_07367_ ), .A3(_07368_ ), .ZN(_07369_ ) );
OAI21_X1 _28206_ ( .A(_07153_ ), .B1(_07037_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07370_ ) );
OAI21_X1 _28207_ ( .A(_07361_ ), .B1(_07369_ ), .B2(_07370_ ), .ZN(_07371_ ) );
NAND4_X1 _28208_ ( .A1(_06665_ ), .A2(_06725_ ), .A3(_05083_ ), .A4(_06611_ ), .ZN(_07372_ ) );
OR2_X1 _28209_ ( .A1(_06655_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07373_ ) );
NAND3_X1 _28210_ ( .A1(_07371_ ), .A2(_07372_ ), .A3(_07373_ ), .ZN(_07374_ ) );
OAI21_X1 _28211_ ( .A(_06661_ ), .B1(_06809_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07375_ ) );
OAI21_X1 _28212_ ( .A(_07360_ ), .B1(_07374_ ), .B2(_07375_ ), .ZN(_07376_ ) );
NAND4_X1 _28213_ ( .A1(_06907_ ), .A2(_06757_ ), .A3(_05091_ ), .A4(_06831_ ), .ZN(_07377_ ) );
OR3_X1 _28214_ ( .A1(_07188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11125_ ), .ZN(_07378_ ) );
NAND3_X1 _28215_ ( .A1(_07376_ ), .A2(_07377_ ), .A3(_07378_ ), .ZN(_07379_ ) );
AND4_X1 _28216_ ( .A1(_05095_ ), .A2(_07057_ ), .A3(_06910_ ), .A4(_06846_ ), .ZN(_07380_ ) );
NOR2_X1 _28217_ ( .A1(_06824_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07381_ ) );
NOR3_X1 _28218_ ( .A1(_07379_ ), .A2(_07380_ ), .A3(_07381_ ), .ZN(_07382_ ) );
NAND4_X1 _28219_ ( .A1(_06721_ ), .A2(_06916_ ), .A3(_05099_ ), .A4(_06750_ ), .ZN(_07383_ ) );
AOI22_X1 _28220_ ( .A1(_07055_ ), .A2(_05101_ ), .B1(_06596_ ), .B2(_06694_ ), .ZN(_07384_ ) );
NAND3_X1 _28221_ ( .A1(_07382_ ), .A2(_07383_ ), .A3(_07384_ ), .ZN(_07385_ ) );
NAND3_X1 _28222_ ( .A1(_06694_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06852_ ), .ZN(_07386_ ) );
AOI21_X1 _28223_ ( .A(_07359_ ), .B1(_07385_ ), .B2(_07386_ ), .ZN(_07387_ ) );
OR2_X1 _28224_ ( .A1(_06706_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07388_ ) );
NAND4_X1 _28225_ ( .A1(_06755_ ), .A2(_06926_ ), .A3(_05109_ ), .A4(_07001_ ), .ZN(_07389_ ) );
NAND3_X1 _28226_ ( .A1(_07387_ ), .A2(_07388_ ), .A3(_07389_ ), .ZN(_07390_ ) );
NOR3_X1 _28227_ ( .A1(_06855_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03838_ ), .ZN(_07391_ ) );
AND4_X1 _28228_ ( .A1(_05113_ ), .A2(_06726_ ), .A3(_07066_ ), .A4(_06597_ ), .ZN(_07392_ ) );
NOR3_X1 _28229_ ( .A1(_07390_ ), .A2(_07391_ ), .A3(_07392_ ), .ZN(_07393_ ) );
NAND4_X1 _28230_ ( .A1(_06947_ ), .A2(_07010_ ), .A3(_05116_ ), .A4(_07011_ ), .ZN(_07394_ ) );
NAND4_X1 _28231_ ( .A1(_06756_ ), .A2(_07071_ ), .A3(_05118_ ), .A4(_07011_ ), .ZN(_07395_ ) );
AND3_X1 _28232_ ( .A1(_07393_ ), .A2(_07394_ ), .A3(_07395_ ), .ZN(_07396_ ) );
OR2_X1 _28233_ ( .A1(_06944_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07397_ ) );
NAND4_X1 _28234_ ( .A1(_06949_ ), .A2(_07067_ ), .A3(_05123_ ), .A4(_07018_ ), .ZN(_07398_ ) );
NAND3_X1 _28235_ ( .A1(_07396_ ), .A2(_07397_ ), .A3(_07398_ ), .ZN(_07399_ ) );
NOR2_X1 _28236_ ( .A1(_06870_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07400_ ) );
OAI21_X1 _28237_ ( .A(_06600_ ), .B1(_06872_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07401_ ) );
NOR3_X1 _28238_ ( .A1(_07399_ ), .A2(_07400_ ), .A3(_07401_ ), .ZN(_07402_ ) );
NAND3_X1 _28239_ ( .A1(_07251_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_07080_ ), .ZN(_07403_ ) );
NAND4_X1 _28240_ ( .A1(_06956_ ), .A2(_06957_ ), .A3(_06877_ ), .A4(_07403_ ), .ZN(_07404_ ) );
OAI211_X1 _28241_ ( .A(_07356_ ), .B(_07358_ ), .C1(_07402_ ), .C2(_07404_ ), .ZN(\idu.io_out_bits_rs2_data [13] ) );
NAND2_X1 _28242_ ( .A1(\exu.io_out_bits_rd_wdata [12] ), .A2(_06879_ ), .ZN(_07405_ ) );
AND4_X1 _28243_ ( .A1(\wbu.io_in_bits_rd_wdata [12] ), .A2(_06782_ ), .A3(_07138_ ), .A4(_06780_ ), .ZN(_07406_ ) );
AOI21_X1 _28244_ ( .A(_07406_ ), .B1(\lsu.io_out_bits_rd_wdata [12] ), .B2(_06784_ ), .ZN(_07407_ ) );
AND3_X1 _28245_ ( .A1(_06730_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06607_ ), .ZN(_07408_ ) );
OR3_X1 _28246_ ( .A1(_06990_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11124_ ), .ZN(_07409_ ) );
NAND3_X1 _28247_ ( .A1(_06679_ ), .A2(_05147_ ), .A3(_11051_ ), .ZN(_07410_ ) );
OAI21_X1 _28248_ ( .A(_07410_ ), .B1(_10688_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07411_ ) );
AND4_X1 _28249_ ( .A1(_05150_ ), .A2(_06586_ ), .A3(_06682_ ), .A4(_06653_ ), .ZN(_07412_ ) );
NOR3_X1 _28250_ ( .A1(_06794_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11122_ ), .ZN(_07413_ ) );
NOR3_X1 _28251_ ( .A1(_07411_ ), .A2(_07412_ ), .A3(_07413_ ), .ZN(_07414_ ) );
NAND4_X1 _28252_ ( .A1(_06627_ ), .A2(_06696_ ), .A3(_05153_ ), .A4(_06796_ ), .ZN(_07415_ ) );
OR2_X1 _28253_ ( .A1(_06633_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07416_ ) );
NAND3_X1 _28254_ ( .A1(_07414_ ), .A2(_07415_ ), .A3(_07416_ ), .ZN(_07417_ ) );
AND4_X1 _28255_ ( .A1(_05158_ ), .A2(_06587_ ), .A3(_06696_ ), .A4(_11052_ ), .ZN(_07418_ ) );
NOR3_X1 _28256_ ( .A1(_06641_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06638_ ), .ZN(_07419_ ) );
NOR3_X1 _28257_ ( .A1(_07417_ ), .A2(_07418_ ), .A3(_07419_ ), .ZN(_07420_ ) );
NAND4_X1 _28258_ ( .A1(_06663_ ), .A2(_07156_ ), .A3(_05162_ ), .A4(_07258_ ), .ZN(_07421_ ) );
NAND4_X1 _28259_ ( .A1(_07215_ ), .A2(_07156_ ), .A3(_05164_ ), .A4(_07258_ ), .ZN(_07422_ ) );
NAND3_X1 _28260_ ( .A1(_07420_ ), .A2(_07421_ ), .A3(_07422_ ), .ZN(_07423_ ) );
NOR2_X1 _28261_ ( .A1(_06651_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07424_ ) );
OAI21_X1 _28262_ ( .A(_06987_ ), .B1(_07106_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07425_ ) );
NOR3_X1 _28263_ ( .A1(_07423_ ), .A2(_07424_ ), .A3(_07425_ ), .ZN(_07426_ ) );
AND3_X1 _28264_ ( .A1(_06749_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03834_ ), .ZN(_07427_ ) );
OAI21_X1 _28265_ ( .A(_07409_ ), .B1(_07426_ ), .B2(_07427_ ), .ZN(_07428_ ) );
AND3_X1 _28266_ ( .A1(_06590_ ), .A2(_05173_ ), .A3(_06845_ ), .ZN(_07429_ ) );
AND4_X1 _28267_ ( .A1(_05175_ ), .A2(_06833_ ), .A3(_06683_ ), .A4(_06594_ ), .ZN(_07430_ ) );
NOR3_X1 _28268_ ( .A1(_07428_ ), .A2(_07429_ ), .A3(_07430_ ), .ZN(_07431_ ) );
OR3_X1 _28269_ ( .A1(_06829_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06611_ ), .ZN(_07432_ ) );
NAND4_X1 _28270_ ( .A1(_06670_ ), .A2(_06834_ ), .A3(_05179_ ), .A4(_11125_ ), .ZN(_07433_ ) );
AND3_X1 _28271_ ( .A1(_07431_ ), .A2(_07432_ ), .A3(_07433_ ), .ZN(_07434_ ) );
NAND4_X1 _28272_ ( .A1(_07057_ ), .A2(_06835_ ), .A3(_05182_ ), .A4(_06741_ ), .ZN(_07435_ ) );
OR3_X1 _28273_ ( .A1(_06843_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06831_ ), .ZN(_07436_ ) );
AND3_X1 _28274_ ( .A1(_07434_ ), .A2(_07435_ ), .A3(_07436_ ), .ZN(_07437_ ) );
OR2_X1 _28275_ ( .A1(_06706_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07438_ ) );
NAND4_X1 _28276_ ( .A1(_06709_ ), .A2(_06710_ ), .A3(_05187_ ), .A4(_01100_ ), .ZN(_07439_ ) );
NAND3_X1 _28277_ ( .A1(_07437_ ), .A2(_07438_ ), .A3(_07439_ ), .ZN(_07440_ ) );
NOR3_X1 _28278_ ( .A1(_06802_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06856_ ), .ZN(_07441_ ) );
AND4_X1 _28279_ ( .A1(_05191_ ), .A2(_06726_ ), .A3(_07066_ ), .A4(_06606_ ), .ZN(_07442_ ) );
NOR3_X1 _28280_ ( .A1(_07440_ ), .A2(_07441_ ), .A3(_07442_ ), .ZN(_07443_ ) );
AOI22_X1 _28281_ ( .A1(_06859_ ), .A2(_05194_ ), .B1(_01101_ ), .B2(_06730_ ), .ZN(_07444_ ) );
AOI21_X1 _28282_ ( .A(_07408_ ), .B1(_07443_ ), .B2(_07444_ ), .ZN(_07445_ ) );
NOR2_X1 _28283_ ( .A1(_06738_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07446_ ) );
NOR3_X1 _28284_ ( .A1(_07445_ ), .A2(_06742_ ), .A3(_07446_ ), .ZN(_07447_ ) );
AND4_X1 _28285_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_06758_ ), .A3(_07067_ ), .A4(_06938_ ), .ZN(_07448_ ) );
OAI221_X1 _28286_ ( .A(_06872_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06870_ ), .C1(_07447_ ), .C2(_07448_ ), .ZN(_07449_ ) );
NAND4_X1 _28287_ ( .A1(_06756_ ), .A2(_06949_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A4(\idu.immI [4] ), .ZN(_07450_ ) );
AOI21_X1 _28288_ ( .A(_06598_ ), .B1(_07449_ ), .B2(_07450_ ), .ZN(_07451_ ) );
NAND3_X1 _28289_ ( .A1(_07251_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_07080_ ), .ZN(_07452_ ) );
NAND4_X1 _28290_ ( .A1(_06956_ ), .A2(_06957_ ), .A3(_06877_ ), .A4(_07452_ ), .ZN(_07453_ ) );
OAI211_X1 _28291_ ( .A(_07405_ ), .B(_07407_ ), .C1(_07451_ ), .C2(_07453_ ), .ZN(\idu.io_out_bits_rs2_data [12] ) );
OAI21_X1 _28292_ ( .A(_06767_ ), .B1(_02658_ ), .B2(_02659_ ), .ZN(_07454_ ) );
AND4_X1 _28293_ ( .A1(\wbu.io_in_bits_rd_wdata [29] ), .A2(_06782_ ), .A3(_07138_ ), .A4(_06780_ ), .ZN(_07455_ ) );
AOI21_X1 _28294_ ( .A(_07455_ ), .B1(\lsu.io_out_bits_rd_wdata [29] ), .B2(_06784_ ), .ZN(_07456_ ) );
OR2_X1 _28295_ ( .A1(_06943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07457_ ) );
NAND3_X1 _28296_ ( .A1(_06604_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06607_ ), .ZN(_07458_ ) );
NOR3_X1 _28297_ ( .A1(_06844_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06847_ ), .ZN(_07459_ ) );
AND4_X1 _28298_ ( .A1(_05235_ ), .A2(_07215_ ), .A3(_07156_ ), .A4(_07258_ ), .ZN(_07460_ ) );
NAND3_X1 _28299_ ( .A1(_06703_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11052_ ), .ZN(_07461_ ) );
AND4_X1 _28300_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_06586_ ), .A3(_06682_ ), .A4(_06653_ ), .ZN(_07462_ ) );
OR3_X1 _28301_ ( .A1(_06828_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_11121_ ), .ZN(_07463_ ) );
OR3_X1 _28302_ ( .A1(_11126_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11121_ ), .ZN(_07464_ ) );
AND2_X1 _28303_ ( .A1(_07463_ ), .A2(_07464_ ), .ZN(_07465_ ) );
AOI21_X1 _28304_ ( .A(_07462_ ), .B1(_07465_ ), .B2(_07094_ ), .ZN(_07466_ ) );
OAI21_X1 _28305_ ( .A(_06972_ ), .B1(_07264_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07467_ ) );
OAI21_X1 _28306_ ( .A(_07461_ ), .B1(_07466_ ), .B2(_07467_ ), .ZN(_07468_ ) );
NAND4_X1 _28307_ ( .A1(_06668_ ), .A2(_07210_ ), .A3(_05229_ ), .A4(_06674_ ), .ZN(_07469_ ) );
OR3_X1 _28308_ ( .A1(_06636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06592_ ), .ZN(_07470_ ) );
AND3_X1 _28309_ ( .A1(_07468_ ), .A2(_07469_ ), .A3(_07470_ ), .ZN(_07471_ ) );
OR3_X1 _28310_ ( .A1(_06641_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11123_ ), .ZN(_07472_ ) );
NAND3_X1 _28311_ ( .A1(_07471_ ), .A2(_06647_ ), .A3(_07472_ ), .ZN(_07473_ ) );
NAND3_X1 _28312_ ( .A1(_06858_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03834_ ), .ZN(_07474_ ) );
AOI21_X1 _28313_ ( .A(_07460_ ), .B1(_07473_ ), .B2(_07474_ ), .ZN(_07475_ ) );
NAND4_X1 _28314_ ( .A1(_06898_ ), .A2(_06725_ ), .A3(_05238_ ), .A4(_06816_ ), .ZN(_07476_ ) );
OR2_X1 _28315_ ( .A1(_06661_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07477_ ) );
AND3_X1 _28316_ ( .A1(_07475_ ), .A2(_07476_ ), .A3(_07477_ ), .ZN(_07478_ ) );
NAND4_X1 _28317_ ( .A1(_06720_ ), .A2(_06666_ ), .A3(_05241_ ), .A4(_06817_ ), .ZN(_07479_ ) );
NAND4_X1 _28318_ ( .A1(_06670_ ), .A2(_06666_ ), .A3(_05243_ ), .A4(_06817_ ), .ZN(_07480_ ) );
NAND3_X1 _28319_ ( .A1(_07478_ ), .A2(_07479_ ), .A3(_07480_ ), .ZN(_07481_ ) );
NOR2_X1 _28320_ ( .A1(_06677_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07482_ ) );
NOR2_X1 _28321_ ( .A1(_06824_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07483_ ) );
NOR3_X1 _28322_ ( .A1(_07481_ ), .A2(_07482_ ), .A3(_07483_ ), .ZN(_07484_ ) );
NAND4_X1 _28323_ ( .A1(_06721_ ), .A2(_06835_ ), .A3(_05249_ ), .A4(_06741_ ), .ZN(_07485_ ) );
AOI22_X1 _28324_ ( .A1(_07055_ ), .A2(_05251_ ), .B1(_01099_ ), .B2(_06694_ ), .ZN(_07486_ ) );
NAND3_X1 _28325_ ( .A1(_07484_ ), .A2(_07485_ ), .A3(_07486_ ), .ZN(_07487_ ) );
NAND3_X1 _28326_ ( .A1(_06694_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06606_ ), .ZN(_07488_ ) );
AOI21_X1 _28327_ ( .A(_07459_ ), .B1(_07487_ ), .B2(_07488_ ), .ZN(_07489_ ) );
NAND4_X1 _28328_ ( .A1(_06850_ ), .A2(_06711_ ), .A3(_05256_ ), .A4(_06597_ ), .ZN(_07490_ ) );
OR2_X1 _28329_ ( .A1(_06930_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07491_ ) );
NAND3_X1 _28330_ ( .A1(_07489_ ), .A2(_07490_ ), .A3(_07491_ ), .ZN(_07492_ ) );
OAI21_X1 _28331_ ( .A(_06933_ ), .B1(_06717_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07493_ ) );
OAI21_X1 _28332_ ( .A(_07458_ ), .B1(_07492_ ), .B2(_07493_ ), .ZN(_07494_ ) );
NAND4_X1 _28333_ ( .A1(_06947_ ), .A2(_07071_ ), .A3(_05263_ ), .A4(_06885_ ), .ZN(_07495_ ) );
OR2_X1 _28334_ ( .A1(_06732_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07496_ ) );
AND4_X1 _28335_ ( .A1(_06738_ ), .A2(_07494_ ), .A3(_07495_ ), .A4(_07496_ ), .ZN(_07497_ ) );
AND4_X1 _28336_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_07058_ ), .A3(_06937_ ), .A4(_01102_ ), .ZN(_07498_ ) );
OAI21_X1 _28337_ ( .A(_07457_ ), .B1(_07497_ ), .B2(_07498_ ), .ZN(_07499_ ) );
NOR2_X1 _28338_ ( .A1(_06870_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07500_ ) );
OAI21_X1 _28339_ ( .A(_07134_ ), .B1(_06872_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07501_ ) );
NOR3_X1 _28340_ ( .A1(_07499_ ), .A2(_07500_ ), .A3(_07501_ ), .ZN(_07502_ ) );
OAI211_X1 _28341_ ( .A(_06875_ ), .B(_06877_ ), .C1(_05272_ ), .C2(_06600_ ), .ZN(_07503_ ) );
OAI211_X1 _28342_ ( .A(_07454_ ), .B(_07456_ ), .C1(_07502_ ), .C2(_07503_ ), .ZN(\idu.io_out_bits_rs2_data [29] ) );
OAI21_X1 _28343_ ( .A(_06767_ ), .B1(_02728_ ), .B2(_02729_ ), .ZN(_07504_ ) );
AND4_X1 _28344_ ( .A1(\wbu.io_in_bits_rd_wdata [11] ), .A2(_06782_ ), .A3(_07138_ ), .A4(_06780_ ), .ZN(_07505_ ) );
AOI21_X1 _28345_ ( .A(_07505_ ), .B1(\lsu.io_out_bits_rd_wdata [11] ), .B2(_06784_ ), .ZN(_07506_ ) );
NAND3_X1 _28346_ ( .A1(_06604_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06728_ ), .ZN(_07507_ ) );
AND4_X1 _28347_ ( .A1(_05312_ ), .A2(_06669_ ), .A3(_06909_ ), .A4(_06611_ ), .ZN(_07508_ ) );
OR3_X1 _28348_ ( .A1(_06827_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10620_ ), .ZN(_07509_ ) );
OR3_X1 _28349_ ( .A1(_11126_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10620_ ), .ZN(_07510_ ) );
NAND4_X1 _28350_ ( .A1(_06586_ ), .A2(_06682_ ), .A3(_05296_ ), .A4(_11049_ ), .ZN(_07511_ ) );
AND3_X1 _28351_ ( .A1(_07509_ ), .A2(_07510_ ), .A3(_07511_ ), .ZN(_07512_ ) );
OR3_X1 _28352_ ( .A1(_06624_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10783_ ), .ZN(_07513_ ) );
NAND3_X1 _28353_ ( .A1(_07512_ ), .A2(_06971_ ), .A3(_07513_ ), .ZN(_07514_ ) );
NAND3_X1 _28354_ ( .A1(_06703_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06653_ ), .ZN(_07515_ ) );
NAND2_X1 _28355_ ( .A1(_07514_ ), .A2(_07515_ ), .ZN(_07516_ ) );
OAI21_X1 _28356_ ( .A(_07516_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06633_ ), .ZN(_07517_ ) );
NOR3_X1 _28357_ ( .A1(_06636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11122_ ), .ZN(_07518_ ) );
AND4_X1 _28358_ ( .A1(_05290_ ), .A2(_06601_ ), .A3(_06683_ ), .A4(_11051_ ), .ZN(_07519_ ) );
OR3_X1 _28359_ ( .A1(_07517_ ), .A2(_07518_ ), .A3(_07519_ ), .ZN(_07520_ ) );
NOR2_X1 _28360_ ( .A1(_06646_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07521_ ) );
AND4_X1 _28361_ ( .A1(_05304_ ), .A2(_06668_ ), .A3(_06723_ ), .A4(_06814_ ), .ZN(_07522_ ) );
OR3_X1 _28362_ ( .A1(_07520_ ), .A2(_07521_ ), .A3(_07522_ ), .ZN(_07523_ ) );
NOR2_X1 _28363_ ( .A1(_06809_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07524_ ) );
OAI21_X1 _28364_ ( .A(_06988_ ), .B1(_07106_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07525_ ) );
OR3_X1 _28365_ ( .A1(_07523_ ), .A2(_07524_ ), .A3(_07525_ ), .ZN(_07526_ ) );
NAND3_X1 _28366_ ( .A1(_06749_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06846_ ), .ZN(_07527_ ) );
AOI21_X1 _28367_ ( .A(_07508_ ), .B1(_07526_ ), .B2(_07527_ ), .ZN(_07528_ ) );
OR2_X1 _28368_ ( .A1(_06677_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07529_ ) );
OR2_X1 _28369_ ( .A1(_06687_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07530_ ) );
NAND3_X1 _28370_ ( .A1(_07528_ ), .A2(_07529_ ), .A3(_07530_ ), .ZN(_07531_ ) );
AND4_X1 _28371_ ( .A1(_05317_ ), .A2(_06720_ ), .A3(_06834_ ), .A4(_06595_ ), .ZN(_07532_ ) );
NOR3_X1 _28372_ ( .A1(_06918_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06919_ ), .ZN(_07533_ ) );
NOR3_X1 _28373_ ( .A1(_07531_ ), .A2(_07532_ ), .A3(_07533_ ), .ZN(_07534_ ) );
NAND3_X1 _28374_ ( .A1(_06694_ ), .A2(_05321_ ), .A3(_06606_ ), .ZN(_07535_ ) );
NAND4_X1 _28375_ ( .A1(_06710_ ), .A2(_07066_ ), .A3(_05289_ ), .A4(_06750_ ), .ZN(_07536_ ) );
AND3_X1 _28376_ ( .A1(_07534_ ), .A2(_07535_ ), .A3(_07536_ ), .ZN(_07537_ ) );
OR2_X1 _28377_ ( .A1(_06706_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07538_ ) );
NAND4_X1 _28378_ ( .A1(_06755_ ), .A2(_07232_ ), .A3(_05327_ ), .A4(_06865_ ), .ZN(_07539_ ) );
NAND3_X1 _28379_ ( .A1(_07537_ ), .A2(_07538_ ), .A3(_07539_ ), .ZN(_07540_ ) );
OAI21_X1 _28380_ ( .A(_06933_ ), .B1(_06717_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07541_ ) );
OAI21_X1 _28381_ ( .A(_07507_ ), .B1(_07540_ ), .B2(_07541_ ), .ZN(_07542_ ) );
NAND4_X1 _28382_ ( .A1(_06947_ ), .A2(_07010_ ), .A3(_05333_ ), .A4(_07011_ ), .ZN(_07543_ ) );
OR2_X1 _28383_ ( .A1(_06940_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07544_ ) );
AND3_X1 _28384_ ( .A1(_07542_ ), .A2(_07543_ ), .A3(_07544_ ), .ZN(_07545_ ) );
NAND4_X1 _28385_ ( .A1(_07058_ ), .A2(_06937_ ), .A3(_05337_ ), .A4(_07018_ ), .ZN(_07546_ ) );
OR2_X1 _28386_ ( .A1(_06943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07547_ ) );
NAND3_X1 _28387_ ( .A1(_07545_ ), .A2(_07546_ ), .A3(_07547_ ), .ZN(_07548_ ) );
NOR2_X1 _28388_ ( .A1(_06870_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07549_ ) );
OAI21_X1 _28389_ ( .A(_07134_ ), .B1(_06872_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07550_ ) );
NOR3_X1 _28390_ ( .A1(_07548_ ), .A2(_07549_ ), .A3(_07550_ ), .ZN(_07551_ ) );
OAI211_X1 _28391_ ( .A(_06875_ ), .B(_06877_ ), .C1(_05344_ ), .C2(_06600_ ), .ZN(_07552_ ) );
OAI211_X1 _28392_ ( .A(_07504_ ), .B(_07506_ ), .C1(_07551_ ), .C2(_07552_ ), .ZN(\idu.io_out_bits_rs2_data [11] ) );
NAND2_X1 _28393_ ( .A1(\exu.io_out_bits_rd_wdata [10] ), .A2(_06879_ ), .ZN(_07553_ ) );
AND4_X1 _28394_ ( .A1(\wbu.io_in_bits_rd_wdata [10] ), .A2(_06782_ ), .A3(_07138_ ), .A4(_06779_ ), .ZN(_07554_ ) );
AOI21_X1 _28395_ ( .A(_07554_ ), .B1(\lsu.io_out_bits_rd_wdata [10] ), .B2(_06783_ ), .ZN(_07555_ ) );
NOR2_X1 _28396_ ( .A1(_06676_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07556_ ) );
NOR2_X1 _28397_ ( .A1(_06651_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07557_ ) );
NOR3_X1 _28398_ ( .A1(_11126_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10783_ ), .ZN(_07558_ ) );
AND3_X1 _28399_ ( .A1(_10651_ ), .A2(_05363_ ), .A3(_11049_ ), .ZN(_07559_ ) );
AND4_X1 _28400_ ( .A1(_05366_ ), .A2(_06586_ ), .A3(_06682_ ), .A4(_11049_ ), .ZN(_07560_ ) );
NOR3_X1 _28401_ ( .A1(_07558_ ), .A2(_07559_ ), .A3(_07560_ ), .ZN(_07561_ ) );
OR3_X1 _28402_ ( .A1(_06624_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10783_ ), .ZN(_07562_ ) );
NAND3_X1 _28403_ ( .A1(_06702_ ), .A2(_05370_ ), .A3(_11050_ ), .ZN(_07563_ ) );
AND3_X1 _28404_ ( .A1(_07561_ ), .A2(_07562_ ), .A3(_07563_ ), .ZN(_07564_ ) );
MUX2_X1 _28405_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_07564_ ), .S(_06633_ ), .Z(_07565_ ) );
NAND4_X1 _28406_ ( .A1(_06897_ ), .A2(_07210_ ), .A3(_05375_ ), .A4(_06674_ ), .ZN(_07566_ ) );
OR3_X1 _28407_ ( .A1(_06641_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06592_ ), .ZN(_07567_ ) );
AND3_X1 _28408_ ( .A1(_07565_ ), .A2(_07566_ ), .A3(_07567_ ), .ZN(_07568_ ) );
OR2_X1 _28409_ ( .A1(_06647_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07569_ ) );
NAND3_X1 _28410_ ( .A1(_07568_ ), .A2(_06655_ ), .A3(_07569_ ), .ZN(_07570_ ) );
NAND3_X1 _28411_ ( .A1(_06730_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06811_ ), .ZN(_07571_ ) );
AOI21_X1 _28412_ ( .A(_07557_ ), .B1(_07570_ ), .B2(_07571_ ), .ZN(_07572_ ) );
NAND4_X1 _28413_ ( .A1(_06909_ ), .A2(_06699_ ), .A3(_05383_ ), .A4(_06845_ ), .ZN(_07573_ ) );
AOI22_X1 _28414_ ( .A1(_06986_ ), .A2(_05386_ ), .B1(_06816_ ), .B2(_06745_ ), .ZN(_07574_ ) );
NAND3_X1 _28415_ ( .A1(_07572_ ), .A2(_07573_ ), .A3(_07574_ ), .ZN(_07575_ ) );
NAND3_X1 _28416_ ( .A1(_06745_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06817_ ), .ZN(_07576_ ) );
AOI21_X1 _28417_ ( .A(_07556_ ), .B1(_07575_ ), .B2(_07576_ ), .ZN(_07577_ ) );
NAND3_X1 _28418_ ( .A1(_06684_ ), .A2(_05390_ ), .A3(_06595_ ), .ZN(_07578_ ) );
NAND4_X1 _28419_ ( .A1(_06720_ ), .A2(_06834_ ), .A3(_05393_ ), .A4(_06595_ ), .ZN(_07579_ ) );
NAND3_X1 _28420_ ( .A1(_07577_ ), .A2(_07578_ ), .A3(_07579_ ), .ZN(_07580_ ) );
NOR3_X1 _28421_ ( .A1(_06918_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07199_ ), .ZN(_07581_ ) );
OAI21_X1 _28422_ ( .A(_06923_ ), .B1(_06840_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07582_ ) );
NOR3_X1 _28423_ ( .A1(_07580_ ), .A2(_07581_ ), .A3(_07582_ ), .ZN(_07583_ ) );
AOI21_X1 _28424_ ( .A(_07583_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06922_ ), .ZN(_07584_ ) );
NOR2_X1 _28425_ ( .A1(_06706_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07585_ ) );
AND3_X1 _28426_ ( .A1(_06631_ ), .A2(_05401_ ), .A3(_06750_ ), .ZN(_07586_ ) );
NOR3_X1 _28427_ ( .A1(_07584_ ), .A2(_07585_ ), .A3(_07586_ ), .ZN(_07587_ ) );
NAND4_X1 _28428_ ( .A1(_07058_ ), .A2(_06926_ ), .A3(_05404_ ), .A4(_06607_ ), .ZN(_07588_ ) );
OR3_X1 _28429_ ( .A1(_06804_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03837_ ), .ZN(_07589_ ) );
AND3_X1 _28430_ ( .A1(_07587_ ), .A2(_07588_ ), .A3(_07589_ ), .ZN(_07590_ ) );
NAND4_X1 _28431_ ( .A1(_06936_ ), .A2(_06937_ ), .A3(_05408_ ), .A4(_06938_ ), .ZN(_07591_ ) );
NAND4_X1 _28432_ ( .A1(_06756_ ), .A2(_07010_ ), .A3(_05410_ ), .A4(_07011_ ), .ZN(_07592_ ) );
NAND3_X1 _28433_ ( .A1(_07590_ ), .A2(_07591_ ), .A3(_07592_ ), .ZN(_07593_ ) );
NOR2_X1 _28434_ ( .A1(_06944_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07594_ ) );
NOR2_X1 _28435_ ( .A1(_06943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07595_ ) );
NOR3_X1 _28436_ ( .A1(_07593_ ), .A2(_07594_ ), .A3(_07595_ ), .ZN(_07596_ ) );
NAND4_X1 _28437_ ( .A1(_06948_ ), .A2(_06949_ ), .A3(_05415_ ), .A4(_06952_ ), .ZN(_07597_ ) );
AOI22_X1 _28438_ ( .A1(_06747_ ), .A2(_05418_ ), .B1(_06952_ ), .B2(_06953_ ), .ZN(_07598_ ) );
AND3_X1 _28439_ ( .A1(_07596_ ), .A2(_07597_ ), .A3(_07598_ ), .ZN(_07599_ ) );
NAND3_X1 _28440_ ( .A1(_07251_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_07080_ ), .ZN(_07600_ ) );
NAND4_X1 _28441_ ( .A1(_06956_ ), .A2(_06957_ ), .A3(_07250_ ), .A4(_07600_ ), .ZN(_07601_ ) );
OAI211_X1 _28442_ ( .A(_07553_ ), .B(_07555_ ), .C1(_07599_ ), .C2(_07601_ ), .ZN(\idu.io_out_bits_rs2_data [10] ) );
NAND2_X1 _28443_ ( .A1(\exu.io_out_bits_rd_wdata [9] ), .A2(_06879_ ), .ZN(_07602_ ) );
AND4_X1 _28444_ ( .A1(\wbu.io_in_bits_rd_wdata [9] ), .A2(_06782_ ), .A3(_07138_ ), .A4(_06779_ ), .ZN(_07603_ ) );
AOI21_X1 _28445_ ( .A(_07603_ ), .B1(\lsu.io_out_bits_rd_wdata [9] ), .B2(_06783_ ), .ZN(_07604_ ) );
OR2_X1 _28446_ ( .A1(_06940_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07605_ ) );
NAND3_X1 _28447_ ( .A1(_06614_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06811_ ), .ZN(_07606_ ) );
NAND3_X1 _28448_ ( .A1(_06703_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11052_ ), .ZN(_07607_ ) );
OR3_X1 _28449_ ( .A1(_06828_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10812_ ), .ZN(_07608_ ) );
OR3_X1 _28450_ ( .A1(_11126_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10812_ ), .ZN(_07609_ ) );
NAND4_X1 _28451_ ( .A1(_06587_ ), .A2(_06833_ ), .A3(_05442_ ), .A4(_06673_ ), .ZN(_07610_ ) );
NAND3_X1 _28452_ ( .A1(_07608_ ), .A2(_07609_ ), .A3(_07610_ ), .ZN(_07611_ ) );
OAI21_X1 _28453_ ( .A(_06972_ ), .B1(_07264_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07612_ ) );
OAI21_X1 _28454_ ( .A(_07607_ ), .B1(_07611_ ), .B2(_07612_ ), .ZN(_07613_ ) );
NAND4_X1 _28455_ ( .A1(_06668_ ), .A2(_07210_ ), .A3(_05447_ ), .A4(_06814_ ), .ZN(_07614_ ) );
OR3_X1 _28456_ ( .A1(_06636_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06592_ ), .ZN(_07615_ ) );
AND3_X1 _28457_ ( .A1(_07613_ ), .A2(_07614_ ), .A3(_07615_ ), .ZN(_07616_ ) );
OR3_X1 _28458_ ( .A1(_06641_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11123_ ), .ZN(_07617_ ) );
NAND4_X1 _28459_ ( .A1(_06663_ ), .A2(_07156_ ), .A3(_05452_ ), .A4(_06815_ ), .ZN(_07618_ ) );
NAND3_X1 _28460_ ( .A1(_07616_ ), .A2(_07617_ ), .A3(_07618_ ), .ZN(_07619_ ) );
OAI21_X1 _28461_ ( .A(_06651_ ), .B1(_06655_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07620_ ) );
OAI21_X1 _28462_ ( .A(_07606_ ), .B1(_07619_ ), .B2(_07620_ ), .ZN(_07621_ ) );
NAND4_X1 _28463_ ( .A1(_06909_ ), .A2(_06699_ ), .A3(_05457_ ), .A4(_06816_ ), .ZN(_07622_ ) );
OR2_X1 _28464_ ( .A1(_06988_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07623_ ) );
NAND3_X1 _28465_ ( .A1(_07621_ ), .A2(_07622_ ), .A3(_07623_ ), .ZN(_07624_ ) );
NOR3_X1 _28466_ ( .A1(_07110_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06690_ ), .ZN(_07625_ ) );
OAI21_X1 _28467_ ( .A(_06686_ ), .B1(_06676_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07626_ ) );
NOR3_X1 _28468_ ( .A1(_07624_ ), .A2(_07625_ ), .A3(_07626_ ), .ZN(_07627_ ) );
AOI21_X1 _28469_ ( .A(_07627_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06685_ ), .ZN(_07628_ ) );
NOR3_X1 _28470_ ( .A1(_06830_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06919_ ), .ZN(_07629_ ) );
AND3_X1 _28471_ ( .A1(_06966_ ), .A2(_05467_ ), .A3(_06691_ ), .ZN(_07630_ ) );
NOR3_X1 _28472_ ( .A1(_07628_ ), .A2(_07629_ ), .A3(_07630_ ), .ZN(_07631_ ) );
NAND4_X1 _28473_ ( .A1(_07058_ ), .A2(_06916_ ), .A3(_05469_ ), .A4(_06750_ ), .ZN(_07632_ ) );
OR3_X1 _28474_ ( .A1(_06843_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03836_ ), .ZN(_07633_ ) );
AND3_X1 _28475_ ( .A1(_07631_ ), .A2(_07632_ ), .A3(_07633_ ), .ZN(_07634_ ) );
NAND4_X1 _28476_ ( .A1(_06850_ ), .A2(_07232_ ), .A3(_05473_ ), .A4(_06865_ ), .ZN(_07635_ ) );
NAND4_X1 _28477_ ( .A1(_06709_ ), .A2(_07232_ ), .A3(_05476_ ), .A4(_06865_ ), .ZN(_07636_ ) );
NAND3_X1 _28478_ ( .A1(_07634_ ), .A2(_07635_ ), .A3(_07636_ ), .ZN(_07637_ ) );
NOR3_X1 _28479_ ( .A1(_06855_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07007_ ), .ZN(_07638_ ) );
OAI21_X1 _28480_ ( .A(_06860_ ), .B1(_06933_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07639_ ) );
NOR3_X1 _28481_ ( .A1(_07637_ ), .A2(_07638_ ), .A3(_07639_ ), .ZN(_07640_ ) );
AND3_X1 _28482_ ( .A1(_06858_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06728_ ), .ZN(_07641_ ) );
OAI21_X1 _28483_ ( .A(_07605_ ), .B1(_07640_ ), .B2(_07641_ ), .ZN(_07642_ ) );
AND3_X1 _28484_ ( .A1(_06735_ ), .A2(_05484_ ), .A3(_06938_ ), .ZN(_07643_ ) );
NOR2_X1 _28485_ ( .A1(_06943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07644_ ) );
NOR3_X1 _28486_ ( .A1(_07642_ ), .A2(_07643_ ), .A3(_07644_ ), .ZN(_07645_ ) );
NAND4_X1 _28487_ ( .A1(_06948_ ), .A2(_06949_ ), .A3(_05488_ ), .A4(_06952_ ), .ZN(_07646_ ) );
AOI22_X1 _28488_ ( .A1(_06747_ ), .A2(_05491_ ), .B1(_06952_ ), .B2(_06591_ ), .ZN(_07647_ ) );
AND3_X1 _28489_ ( .A1(_07645_ ), .A2(_07646_ ), .A3(_07647_ ), .ZN(_07648_ ) );
NAND3_X1 _28490_ ( .A1(_07251_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_07080_ ), .ZN(_07649_ ) );
NAND4_X1 _28491_ ( .A1(_06956_ ), .A2(_06957_ ), .A3(_07250_ ), .A4(_07649_ ), .ZN(_07650_ ) );
OAI211_X1 _28492_ ( .A(_07602_ ), .B(_07604_ ), .C1(_07648_ ), .C2(_07650_ ), .ZN(\idu.io_out_bits_rs2_data [9] ) );
NAND2_X1 _28493_ ( .A1(\exu.io_out_bits_rd_wdata [8] ), .A2(_06560_ ), .ZN(_07651_ ) );
AND4_X1 _28494_ ( .A1(\wbu.io_in_bits_rd_wdata [8] ), .A2(_07084_ ), .A3(_03990_ ), .A4(_06576_ ), .ZN(_07652_ ) );
AOI21_X1 _28495_ ( .A(_07652_ ), .B1(\lsu.io_out_bits_rd_wdata [8] ), .B2(_06581_ ), .ZN(_07653_ ) );
NAND3_X1 _28496_ ( .A1(_06761_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(\idu.immI [4] ), .ZN(_07654_ ) );
NAND3_X1 _28497_ ( .A1(_06858_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06728_ ), .ZN(_07655_ ) );
NAND3_X1 _28498_ ( .A1(_06679_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01099_ ), .ZN(_07656_ ) );
OR3_X1 _28499_ ( .A1(_06640_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11122_ ), .ZN(_07657_ ) );
OR3_X1 _28500_ ( .A1(_11126_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10783_ ), .ZN(_07658_ ) );
OAI21_X1 _28501_ ( .A(_07658_ ), .B1(_06791_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_07659_ ) );
NOR2_X1 _28502_ ( .A1(_07094_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07660_ ) );
AOI211_X1 _28503_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_06625_ ), .C1(\idu.io_in_bits_inst [24] ), .C2(_10646_ ), .ZN(_07661_ ) );
NOR3_X1 _28504_ ( .A1(_07659_ ), .A2(_07660_ ), .A3(_07661_ ), .ZN(_07662_ ) );
OR2_X1 _28505_ ( .A1(_06971_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07663_ ) );
NOR2_X1 _28506_ ( .A1(_06633_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07664_ ) );
NOR2_X1 _28507_ ( .A1(_07664_ ), .A2(_07036_ ), .ZN(_07665_ ) );
AND3_X1 _28508_ ( .A1(_07662_ ), .A2(_07663_ ), .A3(_07665_ ), .ZN(_07666_ ) );
AND3_X1 _28509_ ( .A1(_06635_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03832_ ), .ZN(_07667_ ) );
OAI21_X1 _28510_ ( .A(_07657_ ), .B1(_07666_ ), .B2(_07667_ ), .ZN(_07668_ ) );
AND3_X1 _28511_ ( .A1(_06858_ ), .A2(_05522_ ), .A3(_06796_ ), .ZN(_07669_ ) );
AND4_X1 _28512_ ( .A1(_05524_ ), .A2(_10685_ ), .A3(_06601_ ), .A4(_03832_ ), .ZN(_07670_ ) );
OR3_X1 _28513_ ( .A1(_07668_ ), .A2(_07669_ ), .A3(_07670_ ), .ZN(_07671_ ) );
NOR2_X1 _28514_ ( .A1(_06651_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07672_ ) );
OAI21_X1 _28515_ ( .A(_06988_ ), .B1(_07106_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07673_ ) );
NOR3_X1 _28516_ ( .A1(_07671_ ), .A2(_07672_ ), .A3(_07673_ ), .ZN(_07674_ ) );
AND3_X1 _28517_ ( .A1(_06749_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03834_ ), .ZN(_07675_ ) );
NOR2_X1 _28518_ ( .A1(_07674_ ), .A2(_07675_ ), .ZN(_07676_ ) );
AOI211_X1 _28519_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_07110_ ), .C1(\idu.io_in_bits_inst [24] ), .C2(_04003_ ), .ZN(_07677_ ) );
NOR2_X1 _28520_ ( .A1(_06676_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07678_ ) );
OR3_X1 _28521_ ( .A1(_07676_ ), .A2(_07677_ ), .A3(_07678_ ), .ZN(_07679_ ) );
OAI21_X1 _28522_ ( .A(_06681_ ), .B1(_06824_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07680_ ) );
OAI21_X1 _28523_ ( .A(_07656_ ), .B1(_07679_ ), .B2(_07680_ ), .ZN(_07681_ ) );
NAND4_X1 _28524_ ( .A1(_06708_ ), .A2(_06916_ ), .A3(_05537_ ), .A4(_06596_ ), .ZN(_07682_ ) );
OR2_X1 _28525_ ( .A1(_06840_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07683_ ) );
NAND3_X1 _28526_ ( .A1(_07681_ ), .A2(_07682_ ), .A3(_07683_ ), .ZN(_07684_ ) );
AND4_X1 _28527_ ( .A1(_05541_ ), .A2(_06698_ ), .A3(_06699_ ), .A4(_06741_ ), .ZN(_07685_ ) );
NOR2_X1 _28528_ ( .A1(_06706_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07686_ ) );
NOR3_X1 _28529_ ( .A1(_07684_ ), .A2(_07685_ ), .A3(_07686_ ), .ZN(_07687_ ) );
NAND4_X1 _28530_ ( .A1(_06709_ ), .A2(_06711_ ), .A3(_05545_ ), .A4(_06597_ ), .ZN(_07688_ ) );
OR3_X1 _28531_ ( .A1(_06802_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06847_ ), .ZN(_07689_ ) );
NAND3_X1 _28532_ ( .A1(_07687_ ), .A2(_07688_ ), .A3(_07689_ ), .ZN(_07690_ ) );
OAI21_X1 _28533_ ( .A(_06860_ ), .B1(_06933_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07691_ ) );
OAI21_X1 _28534_ ( .A(_07655_ ), .B1(_07690_ ), .B2(_07691_ ), .ZN(_07692_ ) );
NAND4_X1 _28535_ ( .A1(_06755_ ), .A2(_07071_ ), .A3(_05552_ ), .A4(_06866_ ), .ZN(_07693_ ) );
OR2_X1 _28536_ ( .A1(_06737_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07694_ ) );
AND3_X1 _28537_ ( .A1(_07692_ ), .A2(_07693_ ), .A3(_07694_ ), .ZN(_07695_ ) );
OR2_X1 _28538_ ( .A1(_06743_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07696_ ) );
NAND4_X1 _28539_ ( .A1(_06948_ ), .A2(_06758_ ), .A3(_05558_ ), .A4(_06883_ ), .ZN(_07697_ ) );
NAND3_X1 _28540_ ( .A1(_07695_ ), .A2(_07696_ ), .A3(_07697_ ), .ZN(_07698_ ) );
OAI21_X1 _28541_ ( .A(_07134_ ), .B1(_06748_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07699_ ) );
OAI21_X1 _28542_ ( .A(_07654_ ), .B1(_07698_ ), .B2(_07699_ ), .ZN(_07700_ ) );
OAI221_X1 _28543_ ( .A(_07651_ ), .B1(_06560_ ), .B2(_07653_ ), .C1(_06584_ ), .C2(_07700_ ), .ZN(\idu.io_out_bits_rs2_data [8] ) );
NAND2_X1 _28544_ ( .A1(\exu.io_out_bits_rd_wdata [7] ), .A2(_06879_ ), .ZN(_07701_ ) );
AND4_X1 _28545_ ( .A1(\wbu.io_in_bits_rd_wdata [7] ), .A2(_06782_ ), .A3(_07138_ ), .A4(_06779_ ), .ZN(_07702_ ) );
AOI21_X1 _28546_ ( .A(_07702_ ), .B1(\lsu.io_out_bits_rd_wdata [7] ), .B2(_06783_ ), .ZN(_07703_ ) );
NAND3_X1 _28547_ ( .A1(_06658_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06817_ ), .ZN(_07704_ ) );
NAND3_X1 _28548_ ( .A1(_06603_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06811_ ), .ZN(_07705_ ) );
NOR3_X1 _28549_ ( .A1(_06843_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11123_ ), .ZN(_07706_ ) );
OR3_X1 _28550_ ( .A1(_11127_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06592_ ), .ZN(_07707_ ) );
OR3_X1 _28551_ ( .A1(_06829_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_06592_ ), .ZN(_07708_ ) );
NAND3_X1 _28552_ ( .A1(_07707_ ), .A2(_07094_ ), .A3(_07708_ ), .ZN(_07709_ ) );
NAND3_X1 _28553_ ( .A1(_06694_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03833_ ), .ZN(_07710_ ) );
AOI21_X1 _28554_ ( .A(_07706_ ), .B1(_07709_ ), .B2(_07710_ ), .ZN(_07711_ ) );
NAND4_X1 _28555_ ( .A1(_06664_ ), .A2(_06697_ ), .A3(_05580_ ), .A4(_06610_ ), .ZN(_07712_ ) );
OR2_X1 _28556_ ( .A1(_06799_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07713_ ) );
NAND3_X1 _28557_ ( .A1(_07711_ ), .A2(_07712_ ), .A3(_07713_ ), .ZN(_07714_ ) );
OAI21_X1 _28558_ ( .A(_07153_ ), .B1(_07037_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07715_ ) );
OAI21_X1 _28559_ ( .A(_07705_ ), .B1(_07714_ ), .B2(_07715_ ), .ZN(_07716_ ) );
NAND4_X1 _28560_ ( .A1(_06665_ ), .A2(_06725_ ), .A3(_05587_ ), .A4(_06845_ ), .ZN(_07717_ ) );
OR2_X1 _28561_ ( .A1(_06655_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07718_ ) );
NAND3_X1 _28562_ ( .A1(_07716_ ), .A2(_07717_ ), .A3(_07718_ ), .ZN(_07719_ ) );
OAI21_X1 _28563_ ( .A(_06661_ ), .B1(_06809_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07720_ ) );
OAI21_X1 _28564_ ( .A(_07704_ ), .B1(_07719_ ), .B2(_07720_ ), .ZN(_07721_ ) );
NAND4_X1 _28565_ ( .A1(_06907_ ), .A2(_06910_ ), .A3(_05573_ ), .A4(_06612_ ), .ZN(_07722_ ) );
OR3_X1 _28566_ ( .A1(_07188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06690_ ), .ZN(_07723_ ) );
NAND3_X1 _28567_ ( .A1(_07721_ ), .A2(_07722_ ), .A3(_07723_ ), .ZN(_07724_ ) );
AND4_X1 _28568_ ( .A1(_05596_ ), .A2(_07057_ ), .A3(_06666_ ), .A4(_06846_ ), .ZN(_07725_ ) );
NOR2_X1 _28569_ ( .A1(_06824_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07726_ ) );
NOR3_X1 _28570_ ( .A1(_07724_ ), .A2(_07725_ ), .A3(_07726_ ), .ZN(_07727_ ) );
OR3_X1 _28571_ ( .A1(_06830_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06919_ ), .ZN(_07728_ ) );
NAND4_X1 _28572_ ( .A1(_06708_ ), .A2(_06916_ ), .A3(_05602_ ), .A4(_06596_ ), .ZN(_07729_ ) );
NAND3_X1 _28573_ ( .A1(_07727_ ), .A2(_07728_ ), .A3(_07729_ ), .ZN(_07730_ ) );
NOR2_X1 _28574_ ( .A1(_06841_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07731_ ) );
NOR3_X1 _28575_ ( .A1(_06844_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03837_ ), .ZN(_07732_ ) );
NOR3_X1 _28576_ ( .A1(_07730_ ), .A2(_07731_ ), .A3(_07732_ ), .ZN(_07733_ ) );
NAND4_X1 _28577_ ( .A1(_06850_ ), .A2(_06926_ ), .A3(_05607_ ), .A4(_07001_ ), .ZN(_07734_ ) );
NAND4_X1 _28578_ ( .A1(_06755_ ), .A2(_07232_ ), .A3(_05610_ ), .A4(_07001_ ), .ZN(_07735_ ) );
NAND3_X1 _28579_ ( .A1(_07733_ ), .A2(_07734_ ), .A3(_07735_ ), .ZN(_07736_ ) );
NOR3_X1 _28580_ ( .A1(_06855_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07007_ ), .ZN(_07737_ ) );
NOR3_X1 _28581_ ( .A1(_07006_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07007_ ), .ZN(_07738_ ) );
NOR3_X1 _28582_ ( .A1(_07736_ ), .A2(_07737_ ), .A3(_07738_ ), .ZN(_07739_ ) );
NAND4_X1 _28583_ ( .A1(_06936_ ), .A2(_06937_ ), .A3(_05615_ ), .A4(_06938_ ), .ZN(_07740_ ) );
NAND4_X1 _28584_ ( .A1(_06756_ ), .A2(_07010_ ), .A3(_05618_ ), .A4(_07011_ ), .ZN(_07741_ ) );
NAND3_X1 _28585_ ( .A1(_07739_ ), .A2(_07740_ ), .A3(_07741_ ), .ZN(_07742_ ) );
NOR2_X1 _28586_ ( .A1(_06944_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07743_ ) );
AND3_X1 _28587_ ( .A1(_06740_ ), .A2(_05622_ ), .A3(_06938_ ), .ZN(_07744_ ) );
NOR3_X1 _28588_ ( .A1(_07742_ ), .A2(_07743_ ), .A3(_07744_ ), .ZN(_07745_ ) );
NAND4_X1 _28589_ ( .A1(_06948_ ), .A2(_06949_ ), .A3(_05624_ ), .A4(_06952_ ), .ZN(_07746_ ) );
AOI22_X1 _28590_ ( .A1(_06747_ ), .A2(_05627_ ), .B1(_07018_ ), .B2(_06591_ ), .ZN(_07747_ ) );
AND3_X1 _28591_ ( .A1(_07745_ ), .A2(_07746_ ), .A3(_07747_ ), .ZN(_07748_ ) );
NAND3_X1 _28592_ ( .A1(_07251_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_07080_ ), .ZN(_07749_ ) );
NAND4_X1 _28593_ ( .A1(_06956_ ), .A2(_06957_ ), .A3(_07250_ ), .A4(_07749_ ), .ZN(_07750_ ) );
OAI211_X1 _28594_ ( .A(_07701_ ), .B(_07703_ ), .C1(_07748_ ), .C2(_07750_ ), .ZN(\idu.io_out_bits_rs2_data [7] ) );
NAND2_X1 _28595_ ( .A1(\exu.io_out_bits_rd_wdata [6] ), .A2(_06879_ ), .ZN(_07751_ ) );
AND4_X1 _28596_ ( .A1(\wbu.io_in_bits_rd_wdata [6] ), .A2(_06782_ ), .A3(_07138_ ), .A4(_06779_ ), .ZN(_07752_ ) );
AOI21_X1 _28597_ ( .A(_07752_ ), .B1(\lsu.io_out_bits_rd_wdata [6] ), .B2(_06783_ ), .ZN(_07753_ ) );
NAND3_X1 _28598_ ( .A1(_06740_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06883_ ), .ZN(_07754_ ) );
NAND3_X1 _28599_ ( .A1(_06604_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06885_ ), .ZN(_07755_ ) );
NAND3_X1 _28600_ ( .A1(_06740_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06817_ ), .ZN(_07756_ ) );
OR3_X1 _28601_ ( .A1(_11127_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11122_ ), .ZN(_07757_ ) );
OAI21_X1 _28602_ ( .A(_07757_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .B2(_06791_ ), .ZN(_07758_ ) );
AND4_X1 _28603_ ( .A1(_05647_ ), .A2(_06587_ ), .A3(_06833_ ), .A4(_06796_ ), .ZN(_07759_ ) );
NOR3_X1 _28604_ ( .A1(_06794_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11123_ ), .ZN(_07760_ ) );
NOR3_X1 _28605_ ( .A1(_07758_ ), .A2(_07759_ ), .A3(_07760_ ), .ZN(_07761_ ) );
NAND4_X1 _28606_ ( .A1(_06664_ ), .A2(_06697_ ), .A3(_05651_ ), .A4(_06610_ ), .ZN(_07762_ ) );
OR2_X1 _28607_ ( .A1(_06799_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07763_ ) );
NAND3_X1 _28608_ ( .A1(_07761_ ), .A2(_07762_ ), .A3(_07763_ ), .ZN(_07764_ ) );
AND4_X1 _28609_ ( .A1(_05656_ ), .A2(_06897_ ), .A3(_06697_ ), .A4(_07258_ ), .ZN(_07765_ ) );
NOR3_X1 _28610_ ( .A1(_06804_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11124_ ), .ZN(_07766_ ) );
NOR3_X1 _28611_ ( .A1(_07764_ ), .A2(_07765_ ), .A3(_07766_ ), .ZN(_07767_ ) );
OR2_X1 _28612_ ( .A1(_06647_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07768_ ) );
OR2_X1 _28613_ ( .A1(_06655_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07769_ ) );
NAND3_X1 _28614_ ( .A1(_07767_ ), .A2(_07768_ ), .A3(_07769_ ), .ZN(_07770_ ) );
OAI21_X1 _28615_ ( .A(_06661_ ), .B1(_06809_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07771_ ) );
OAI21_X1 _28616_ ( .A(_07756_ ), .B1(_07770_ ), .B2(_07771_ ), .ZN(_07772_ ) );
NAND4_X1 _28617_ ( .A1(_06907_ ), .A2(_06910_ ), .A3(_05665_ ), .A4(_06612_ ), .ZN(_07773_ ) );
OR3_X1 _28618_ ( .A1(_07188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06690_ ), .ZN(_07774_ ) );
NAND3_X1 _28619_ ( .A1(_07772_ ), .A2(_07773_ ), .A3(_07774_ ), .ZN(_07775_ ) );
AND4_X1 _28620_ ( .A1(_05669_ ), .A2(_07057_ ), .A3(_06910_ ), .A4(_06846_ ), .ZN(_07776_ ) );
NOR2_X1 _28621_ ( .A1(_06824_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07777_ ) );
NOR3_X1 _28622_ ( .A1(_07775_ ), .A2(_07776_ ), .A3(_07777_ ), .ZN(_07778_ ) );
OR3_X1 _28623_ ( .A1(_06830_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06919_ ), .ZN(_07779_ ) );
NAND4_X1 _28624_ ( .A1(_06708_ ), .A2(_06916_ ), .A3(_05675_ ), .A4(_06596_ ), .ZN(_07780_ ) );
NAND3_X1 _28625_ ( .A1(_07778_ ), .A2(_07779_ ), .A3(_07780_ ), .ZN(_07781_ ) );
NOR2_X1 _28626_ ( .A1(_06841_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07782_ ) );
NOR3_X1 _28627_ ( .A1(_06844_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03837_ ), .ZN(_07783_ ) );
NOR3_X1 _28628_ ( .A1(_07781_ ), .A2(_07782_ ), .A3(_07783_ ), .ZN(_07784_ ) );
NAND4_X1 _28629_ ( .A1(_06722_ ), .A2(_06926_ ), .A3(_05681_ ), .A4(_07001_ ), .ZN(_07785_ ) );
OR2_X1 _28630_ ( .A1(_06930_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07786_ ) );
NAND3_X1 _28631_ ( .A1(_07784_ ), .A2(_07785_ ), .A3(_07786_ ), .ZN(_07787_ ) );
OAI21_X1 _28632_ ( .A(_06933_ ), .B1(_06717_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07788_ ) );
OAI21_X1 _28633_ ( .A(_07755_ ), .B1(_07787_ ), .B2(_07788_ ), .ZN(_07789_ ) );
NAND4_X1 _28634_ ( .A1(_06936_ ), .A2(_07010_ ), .A3(_05688_ ), .A4(_06938_ ), .ZN(_07790_ ) );
OR2_X1 _28635_ ( .A1(_06940_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07791_ ) );
NAND3_X1 _28636_ ( .A1(_07789_ ), .A2(_07790_ ), .A3(_07791_ ), .ZN(_07792_ ) );
OAI21_X1 _28637_ ( .A(_06943_ ), .B1(_06944_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07793_ ) );
OAI21_X1 _28638_ ( .A(_07754_ ), .B1(_07792_ ), .B2(_07793_ ), .ZN(_07794_ ) );
NAND4_X1 _28639_ ( .A1(_06948_ ), .A2(_06949_ ), .A3(_05695_ ), .A4(_06952_ ), .ZN(_07795_ ) );
AOI22_X1 _28640_ ( .A1(_06747_ ), .A2(_05697_ ), .B1(_07018_ ), .B2(_06591_ ), .ZN(_07796_ ) );
AND3_X1 _28641_ ( .A1(_07794_ ), .A2(_07795_ ), .A3(_07796_ ), .ZN(_07797_ ) );
NAND3_X1 _28642_ ( .A1(_07251_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_07080_ ), .ZN(_07798_ ) );
NAND4_X1 _28643_ ( .A1(_06956_ ), .A2(_07249_ ), .A3(_07250_ ), .A4(_07798_ ), .ZN(_07799_ ) );
OAI211_X1 _28644_ ( .A(_07751_ ), .B(_07753_ ), .C1(_07797_ ), .C2(_07799_ ), .ZN(\idu.io_out_bits_rs2_data [6] ) );
AND3_X1 _28645_ ( .A1(_03105_ ), .A2(_03106_ ), .A3(_06766_ ), .ZN(_07800_ ) );
NOR3_X1 _28646_ ( .A1(_07195_ ), .A2(_00484_ ), .A3(_07196_ ), .ZN(_07801_ ) );
OAI22_X1 _28647_ ( .A1(\lsu.io_out_bits_rd_wdata [5] ), .A2(_07193_ ), .B1(_07194_ ), .B2(_07801_ ), .ZN(_07802_ ) );
NAND3_X1 _28648_ ( .A1(_06740_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06883_ ), .ZN(_07803_ ) );
AND3_X1 _28649_ ( .A1(_06735_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01101_ ), .ZN(_07804_ ) );
AND4_X1 _28650_ ( .A1(_05705_ ), .A2(_06720_ ), .A3(_06834_ ), .A4(_11125_ ), .ZN(_07805_ ) );
OR3_X1 _28651_ ( .A1(_11126_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10783_ ), .ZN(_07806_ ) );
OAI21_X1 _28652_ ( .A(_07806_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .B2(_06791_ ), .ZN(_07807_ ) );
AOI21_X1 _28653_ ( .A(_07807_ ), .B1(_05711_ ), .B2(_06619_ ), .ZN(_07808_ ) );
OR3_X1 _28654_ ( .A1(_06625_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10812_ ), .ZN(_07809_ ) );
NAND4_X1 _28655_ ( .A1(_06627_ ), .A2(_06628_ ), .A3(_05714_ ), .A4(_06673_ ), .ZN(_07810_ ) );
AND3_X1 _28656_ ( .A1(_07808_ ), .A2(_07809_ ), .A3(_07810_ ), .ZN(_07811_ ) );
OR2_X1 _28657_ ( .A1(_06799_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07812_ ) );
NAND4_X1 _28658_ ( .A1(_06897_ ), .A2(_06696_ ), .A3(_05718_ ), .A4(_06814_ ), .ZN(_07813_ ) );
NAND3_X1 _28659_ ( .A1(_07811_ ), .A2(_07812_ ), .A3(_07813_ ), .ZN(_07814_ ) );
NOR3_X1 _28660_ ( .A1(_06641_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11123_ ), .ZN(_07815_ ) );
AND4_X1 _28661_ ( .A1(_05722_ ), .A2(_06627_ ), .A3(_06723_ ), .A4(_06796_ ), .ZN(_07816_ ) );
NOR3_X1 _28662_ ( .A1(_07814_ ), .A2(_07815_ ), .A3(_07816_ ), .ZN(_07817_ ) );
NAND4_X1 _28663_ ( .A1(_07215_ ), .A2(_06724_ ), .A3(_05725_ ), .A4(_06815_ ), .ZN(_07818_ ) );
OR2_X1 _28664_ ( .A1(_06650_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07819_ ) );
AND3_X1 _28665_ ( .A1(_07817_ ), .A2(_07818_ ), .A3(_07819_ ), .ZN(_07820_ ) );
OR2_X1 _28666_ ( .A1(_07106_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07821_ ) );
NAND4_X1 _28667_ ( .A1(_06664_ ), .A2(_06589_ ), .A3(_05707_ ), .A4(_06811_ ), .ZN(_07822_ ) );
NAND3_X1 _28668_ ( .A1(_07820_ ), .A2(_07821_ ), .A3(_07822_ ), .ZN(_07823_ ) );
NOR3_X1 _28669_ ( .A1(_07110_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06594_ ), .ZN(_07824_ ) );
OAI21_X1 _28670_ ( .A(_06686_ ), .B1(_06676_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07825_ ) );
OR3_X1 _28671_ ( .A1(_07823_ ), .A2(_07824_ ), .A3(_07825_ ), .ZN(_07826_ ) );
NAND3_X1 _28672_ ( .A1(_06684_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06605_ ), .ZN(_07827_ ) );
AOI21_X1 _28673_ ( .A(_07805_ ), .B1(_07826_ ), .B2(_07827_ ), .ZN(_07828_ ) );
OR3_X1 _28674_ ( .A1(_06918_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07199_ ), .ZN(_07829_ ) );
NAND4_X1 _28675_ ( .A1(_07057_ ), .A2(_06916_ ), .A3(_05738_ ), .A4(_06596_ ), .ZN(_07830_ ) );
NAND3_X1 _28676_ ( .A1(_07828_ ), .A2(_07829_ ), .A3(_07830_ ), .ZN(_07831_ ) );
NOR3_X1 _28677_ ( .A1(_06844_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06847_ ), .ZN(_07832_ ) );
AND4_X1 _28678_ ( .A1(_05742_ ), .A2(_06907_ ), .A3(_06698_ ), .A4(_01099_ ), .ZN(_07833_ ) );
NOR3_X1 _28679_ ( .A1(_07831_ ), .A2(_07832_ ), .A3(_07833_ ), .ZN(_07834_ ) );
NAND4_X1 _28680_ ( .A1(_06709_ ), .A2(_06711_ ), .A3(_05745_ ), .A4(_06597_ ), .ZN(_07835_ ) );
OR3_X1 _28681_ ( .A1(_06802_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06847_ ), .ZN(_07836_ ) );
NAND3_X1 _28682_ ( .A1(_07834_ ), .A2(_07835_ ), .A3(_07836_ ), .ZN(_07837_ ) );
NOR3_X1 _28683_ ( .A1(_07006_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06856_ ), .ZN(_07838_ ) );
AND4_X1 _28684_ ( .A1(_05750_ ), .A2(_06721_ ), .A3(_06726_ ), .A4(_06852_ ), .ZN(_07839_ ) );
NOR3_X1 _28685_ ( .A1(_07837_ ), .A2(_07838_ ), .A3(_07839_ ), .ZN(_07840_ ) );
AOI22_X1 _28686_ ( .A1(_06731_ ), .A2(_05753_ ), .B1(_06885_ ), .B2(_06735_ ), .ZN(_07841_ ) );
AOI21_X1 _28687_ ( .A(_07804_ ), .B1(_07840_ ), .B2(_07841_ ), .ZN(_07842_ ) );
OAI21_X1 _28688_ ( .A(_07803_ ), .B1(_07842_ ), .B2(_06742_ ), .ZN(_07843_ ) );
OR2_X1 _28689_ ( .A1(_06752_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07844_ ) );
NOR3_X1 _28690_ ( .A1(_07188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03838_ ), .ZN(_07845_ ) );
NOR2_X1 _28691_ ( .A1(_07845_ ), .A2(_06598_ ), .ZN(_07846_ ) );
AND3_X1 _28692_ ( .A1(_07843_ ), .A2(_07844_ ), .A3(_07846_ ), .ZN(_07847_ ) );
NAND3_X1 _28693_ ( .A1(_06953_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_06950_ ), .ZN(_07848_ ) );
NAND4_X1 _28694_ ( .A1(_07248_ ), .A2(_07249_ ), .A3(_07250_ ), .A4(_07848_ ), .ZN(_07849_ ) );
OAI22_X1 _28695_ ( .A1(_07800_ ), .A2(_07802_ ), .B1(_07847_ ), .B2(_07849_ ), .ZN(\idu.io_out_bits_rs2_data [5] ) );
AND3_X1 _28696_ ( .A1(_03165_ ), .A2(_03166_ ), .A3(_06766_ ), .ZN(_07850_ ) );
NOR3_X1 _28697_ ( .A1(_07195_ ), .A2(_00485_ ), .A3(_07196_ ), .ZN(_07851_ ) );
OAI22_X1 _28698_ ( .A1(\lsu.io_out_bits_rd_wdata [4] ), .A2(_07193_ ), .B1(_07194_ ), .B2(_07851_ ), .ZN(_07852_ ) );
AND3_X1 _28699_ ( .A1(_06635_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01100_ ), .ZN(_07853_ ) );
OR2_X1 _28700_ ( .A1(_06651_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07854_ ) );
OR2_X1 _28701_ ( .A1(_07094_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07855_ ) );
OR3_X1 _28702_ ( .A1(_06828_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_10812_ ), .ZN(_07856_ ) );
OR3_X1 _28703_ ( .A1(_11127_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10812_ ), .ZN(_07857_ ) );
NAND3_X1 _28704_ ( .A1(_07855_ ), .A2(_07856_ ), .A3(_07857_ ), .ZN(_07858_ ) );
AOI211_X1 _28705_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_06625_ ), .C1(\idu.io_in_bits_inst [24] ), .C2(_11030_ ), .ZN(_07859_ ) );
NOR2_X1 _28706_ ( .A1(_06972_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07860_ ) );
NOR3_X1 _28707_ ( .A1(_07858_ ), .A2(_07859_ ), .A3(_07860_ ), .ZN(_07861_ ) );
NAND3_X1 _28708_ ( .A1(_06631_ ), .A2(_05792_ ), .A3(_06674_ ), .ZN(_07862_ ) );
NAND4_X1 _28709_ ( .A1(_06897_ ), .A2(_07210_ ), .A3(_05794_ ), .A4(_06674_ ), .ZN(_07863_ ) );
NAND3_X1 _28710_ ( .A1(_07861_ ), .A2(_07862_ ), .A3(_07863_ ), .ZN(_07864_ ) );
NOR3_X1 _28711_ ( .A1(_06641_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06593_ ), .ZN(_07865_ ) );
OAI21_X1 _28712_ ( .A(_06655_ ), .B1(_06646_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07866_ ) );
NOR3_X1 _28713_ ( .A1(_07864_ ), .A2(_07865_ ), .A3(_07866_ ), .ZN(_07867_ ) );
AND3_X1 _28714_ ( .A1(_06652_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07258_ ), .ZN(_07868_ ) );
OAI21_X1 _28715_ ( .A(_07854_ ), .B1(_07867_ ), .B2(_07868_ ), .ZN(_07869_ ) );
AND3_X1 _28716_ ( .A1(_06658_ ), .A2(_05803_ ), .A3(_06787_ ), .ZN(_07870_ ) );
AND4_X1 _28717_ ( .A1(_05805_ ), .A2(_06664_ ), .A3(_06589_ ), .A4(_06815_ ), .ZN(_07871_ ) );
NOR3_X1 _28718_ ( .A1(_07869_ ), .A2(_07870_ ), .A3(_07871_ ), .ZN(_07872_ ) );
OR3_X1 _28719_ ( .A1(_07110_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11124_ ), .ZN(_07873_ ) );
OR2_X1 _28720_ ( .A1(_06676_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07874_ ) );
AND3_X1 _28721_ ( .A1(_07872_ ), .A2(_07873_ ), .A3(_07874_ ), .ZN(_07875_ ) );
NAND4_X1 _28722_ ( .A1(_06835_ ), .A2(_06699_ ), .A3(_05811_ ), .A4(_06595_ ), .ZN(_07876_ ) );
OR3_X1 _28723_ ( .A1(_06829_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03835_ ), .ZN(_07877_ ) );
NAND3_X1 _28724_ ( .A1(_07875_ ), .A2(_07876_ ), .A3(_07877_ ), .ZN(_07878_ ) );
NOR3_X1 _28725_ ( .A1(_06918_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07199_ ), .ZN(_07879_ ) );
NOR2_X1 _28726_ ( .A1(_06840_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07880_ ) );
NOR3_X1 _28727_ ( .A1(_07878_ ), .A2(_07879_ ), .A3(_07880_ ), .ZN(_07881_ ) );
NAND4_X1 _28728_ ( .A1(_06710_ ), .A2(_07066_ ), .A3(_05818_ ), .A4(_06596_ ), .ZN(_07882_ ) );
OR2_X1 _28729_ ( .A1(_06705_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07883_ ) );
AND3_X1 _28730_ ( .A1(_07881_ ), .A2(_07882_ ), .A3(_07883_ ), .ZN(_07884_ ) );
NOR2_X1 _28731_ ( .A1(_06930_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07885_ ) );
NOR2_X1 _28732_ ( .A1(_07885_ ), .A2(_06716_ ), .ZN(_07886_ ) );
AOI21_X1 _28733_ ( .A(_07853_ ), .B1(_07884_ ), .B2(_07886_ ), .ZN(_07887_ ) );
NOR3_X1 _28734_ ( .A1(_07006_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06856_ ), .ZN(_07888_ ) );
AND3_X1 _28735_ ( .A1(_06858_ ), .A2(_05826_ ), .A3(_06865_ ), .ZN(_07889_ ) );
NOR3_X1 _28736_ ( .A1(_07887_ ), .A2(_07888_ ), .A3(_07889_ ), .ZN(_07890_ ) );
OR2_X1 _28737_ ( .A1(_06940_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07891_ ) );
OR2_X1 _28738_ ( .A1(_06737_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07892_ ) );
NAND3_X1 _28739_ ( .A1(_07890_ ), .A2(_07891_ ), .A3(_07892_ ), .ZN(_07893_ ) );
AND4_X1 _28740_ ( .A1(_05831_ ), .A2(_06757_ ), .A3(_07067_ ), .A4(_06885_ ), .ZN(_07894_ ) );
NOR2_X1 _28741_ ( .A1(_06752_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07895_ ) );
NOR3_X1 _28742_ ( .A1(_07893_ ), .A2(_07894_ ), .A3(_07895_ ), .ZN(_07896_ ) );
OR3_X1 _28743_ ( .A1(_07188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03838_ ), .ZN(_07897_ ) );
AND3_X1 _28744_ ( .A1(_07896_ ), .A2(_06600_ ), .A3(_07897_ ), .ZN(_07898_ ) );
NAND3_X1 _28745_ ( .A1(_06953_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_06950_ ), .ZN(_07899_ ) );
NAND4_X1 _28746_ ( .A1(_07248_ ), .A2(_07249_ ), .A3(_07250_ ), .A4(_07899_ ), .ZN(_07900_ ) );
OAI22_X1 _28747_ ( .A1(_07850_ ), .A2(_07852_ ), .B1(_07898_ ), .B2(_07900_ ), .ZN(\idu.io_out_bits_rs2_data [4] ) );
AND3_X1 _28748_ ( .A1(_03225_ ), .A2(_03226_ ), .A3(_06766_ ), .ZN(_07901_ ) );
NOR3_X1 _28749_ ( .A1(_07195_ ), .A2(_00566_ ), .A3(_07196_ ), .ZN(_07902_ ) );
OAI22_X1 _28750_ ( .A1(\lsu.io_out_bits_rd_wdata [3] ), .A2(_07193_ ), .B1(_07194_ ), .B2(_07902_ ), .ZN(_07903_ ) );
OR3_X1 _28751_ ( .A1(_06829_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06811_ ), .ZN(_07904_ ) );
OR3_X1 _28752_ ( .A1(_11126_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11121_ ), .ZN(_07905_ ) );
OAI21_X1 _28753_ ( .A(_07905_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .B2(_06791_ ), .ZN(_07906_ ) );
AND4_X1 _28754_ ( .A1(_05856_ ), .A2(_06586_ ), .A3(_06682_ ), .A4(_11050_ ), .ZN(_07907_ ) );
NOR3_X1 _28755_ ( .A1(_06625_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10812_ ), .ZN(_07908_ ) );
NOR3_X1 _28756_ ( .A1(_07906_ ), .A2(_07907_ ), .A3(_07908_ ), .ZN(_07909_ ) );
NAND4_X1 _28757_ ( .A1(_06627_ ), .A2(_06628_ ), .A3(_05859_ ), .A4(_03832_ ), .ZN(_07910_ ) );
OR2_X1 _28758_ ( .A1(_06633_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07911_ ) );
NAND3_X1 _28759_ ( .A1(_07909_ ), .A2(_07910_ ), .A3(_07911_ ), .ZN(_07912_ ) );
AND4_X1 _28760_ ( .A1(_05863_ ), .A2(_06587_ ), .A3(_06628_ ), .A4(_06673_ ), .ZN(_07913_ ) );
NOR3_X1 _28761_ ( .A1(_06641_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06638_ ), .ZN(_07914_ ) );
NOR3_X1 _28762_ ( .A1(_07912_ ), .A2(_07913_ ), .A3(_07914_ ), .ZN(_07915_ ) );
NAND4_X1 _28763_ ( .A1(_06663_ ), .A2(_06723_ ), .A3(_05867_ ), .A4(_06609_ ), .ZN(_07916_ ) );
NAND4_X1 _28764_ ( .A1(_06668_ ), .A2(_06723_ ), .A3(_05870_ ), .A4(_06609_ ), .ZN(_07917_ ) );
NAND3_X1 _28765_ ( .A1(_07915_ ), .A2(_07916_ ), .A3(_07917_ ), .ZN(_07918_ ) );
NOR2_X1 _28766_ ( .A1(_06650_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07919_ ) );
NOR2_X1 _28767_ ( .A1(_07106_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07920_ ) );
NOR3_X1 _28768_ ( .A1(_07918_ ), .A2(_07919_ ), .A3(_07920_ ), .ZN(_07921_ ) );
NAND4_X1 _28769_ ( .A1(_06664_ ), .A2(_06589_ ), .A3(_05875_ ), .A4(_06787_ ), .ZN(_07922_ ) );
AOI22_X1 _28770_ ( .A1(_06819_ ), .A2(_05878_ ), .B1(_06787_ ), .B2(_06590_ ), .ZN(_07923_ ) );
NAND3_X1 _28771_ ( .A1(_07921_ ), .A2(_07922_ ), .A3(_07923_ ), .ZN(_07924_ ) );
NAND3_X1 _28772_ ( .A1(_06590_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06845_ ), .ZN(_07925_ ) );
AOI21_X1 _28773_ ( .A(_06685_ ), .B1(_07924_ ), .B2(_07925_ ), .ZN(_07926_ ) );
AND3_X1 _28774_ ( .A1(_06684_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06594_ ), .ZN(_07927_ ) );
OAI21_X1 _28775_ ( .A(_07904_ ), .B1(_07926_ ), .B2(_07927_ ), .ZN(_07928_ ) );
AND4_X1 _28776_ ( .A1(_05885_ ), .A2(_06670_ ), .A3(_06834_ ), .A4(_06690_ ), .ZN(_07929_ ) );
NOR2_X1 _28777_ ( .A1(_06839_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07930_ ) );
NOR3_X1 _28778_ ( .A1(_07928_ ), .A2(_07929_ ), .A3(_07930_ ), .ZN(_07931_ ) );
NAND4_X1 _28779_ ( .A1(_06698_ ), .A2(_06699_ ), .A3(_05889_ ), .A4(_06691_ ), .ZN(_07932_ ) );
NAND4_X1 _28780_ ( .A1(_06907_ ), .A2(_06698_ ), .A3(_05891_ ), .A4(_06691_ ), .ZN(_07933_ ) );
NAND3_X1 _28781_ ( .A1(_07931_ ), .A2(_07932_ ), .A3(_07933_ ), .ZN(_07934_ ) );
NOR2_X1 _28782_ ( .A1(_06929_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07935_ ) );
NOR3_X1 _28783_ ( .A1(_06802_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03836_ ), .ZN(_07936_ ) );
NOR3_X1 _28784_ ( .A1(_07934_ ), .A2(_07935_ ), .A3(_07936_ ), .ZN(_07937_ ) );
NAND4_X1 _28785_ ( .A1(_06726_ ), .A2(_07066_ ), .A3(_05897_ ), .A4(_01100_ ), .ZN(_07938_ ) );
NAND4_X1 _28786_ ( .A1(_06721_ ), .A2(_06726_ ), .A3(_05899_ ), .A4(_06606_ ), .ZN(_07939_ ) );
AND4_X1 _28787_ ( .A1(_06732_ ), .A2(_07937_ ), .A3(_07938_ ), .A4(_07939_ ), .ZN(_07940_ ) );
AOI21_X1 _28788_ ( .A(_07940_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06731_ ), .ZN(_07941_ ) );
NOR2_X1 _28789_ ( .A1(_06738_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07942_ ) );
AND4_X1 _28790_ ( .A1(_05904_ ), .A2(_06757_ ), .A3(_07067_ ), .A4(_01101_ ), .ZN(_07943_ ) );
OR3_X1 _28791_ ( .A1(_07941_ ), .A2(_07942_ ), .A3(_07943_ ), .ZN(_07944_ ) );
NOR2_X1 _28792_ ( .A1(_06870_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07945_ ) );
OAI21_X1 _28793_ ( .A(_07134_ ), .B1(_06748_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07946_ ) );
NOR3_X1 _28794_ ( .A1(_07944_ ), .A2(_07945_ ), .A3(_07946_ ), .ZN(_07947_ ) );
NAND3_X1 _28795_ ( .A1(_06953_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_06950_ ), .ZN(_07948_ ) );
NAND4_X1 _28796_ ( .A1(_07248_ ), .A2(_07249_ ), .A3(_06876_ ), .A4(_07948_ ), .ZN(_07949_ ) );
OAI22_X1 _28797_ ( .A1(_07901_ ), .A2(_07903_ ), .B1(_07947_ ), .B2(_07949_ ), .ZN(\idu.io_out_bits_rs2_data [3] ) );
OR3_X1 _28798_ ( .A1(_03284_ ), .A2(_03285_ ), .A3(_06773_ ), .ZN(_07950_ ) );
AND4_X1 _28799_ ( .A1(\wbu.io_in_bits_rd_wdata [2] ), .A2(_06782_ ), .A3(_06772_ ), .A4(_06779_ ), .ZN(_07951_ ) );
AOI21_X1 _28800_ ( .A(_07951_ ), .B1(\lsu.io_out_bits_rd_wdata [2] ), .B2(_06783_ ), .ZN(_07952_ ) );
NAND3_X1 _28801_ ( .A1(_06761_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(\idu.immI [4] ), .ZN(_07953_ ) );
NAND3_X1 _28802_ ( .A1(_06604_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06607_ ), .ZN(_07954_ ) );
AND4_X1 _28803_ ( .A1(_05927_ ), .A2(_10685_ ), .A3(_06696_ ), .A4(_11052_ ), .ZN(_07955_ ) );
OR3_X1 _28804_ ( .A1(_06828_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_11121_ ), .ZN(_07956_ ) );
OAI21_X1 _28805_ ( .A(_07956_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_10688_ ), .ZN(_07957_ ) );
AND4_X1 _28806_ ( .A1(_05931_ ), .A2(_06586_ ), .A3(_06682_ ), .A4(_06653_ ), .ZN(_07958_ ) );
OAI21_X1 _28807_ ( .A(_06971_ ), .B1(_07264_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07959_ ) );
OR3_X1 _28808_ ( .A1(_07957_ ), .A2(_07958_ ), .A3(_07959_ ), .ZN(_07960_ ) );
NAND3_X1 _28809_ ( .A1(_06703_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06609_ ), .ZN(_07961_ ) );
AOI21_X1 _28810_ ( .A(_07955_ ), .B1(_07960_ ), .B2(_07961_ ), .ZN(_07962_ ) );
OR3_X1 _28811_ ( .A1(_06637_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06638_ ), .ZN(_07963_ ) );
NAND4_X1 _28812_ ( .A1(_07156_ ), .A2(_06683_ ), .A3(_05925_ ), .A4(_07258_ ), .ZN(_07964_ ) );
NAND3_X1 _28813_ ( .A1(_07962_ ), .A2(_07963_ ), .A3(_07964_ ), .ZN(_07965_ ) );
NOR2_X1 _28814_ ( .A1(_06647_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07966_ ) );
AND4_X1 _28815_ ( .A1(_05944_ ), .A2(_07215_ ), .A3(_07156_ ), .A4(_03833_ ), .ZN(_07967_ ) );
NOR3_X1 _28816_ ( .A1(_07965_ ), .A2(_07966_ ), .A3(_07967_ ), .ZN(_07968_ ) );
NAND4_X1 _28817_ ( .A1(_06898_ ), .A2(_06725_ ), .A3(_05947_ ), .A4(_06816_ ), .ZN(_07969_ ) );
OR2_X1 _28818_ ( .A1(_07106_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07970_ ) );
NAND3_X1 _28819_ ( .A1(_07968_ ), .A2(_07969_ ), .A3(_07970_ ), .ZN(_07971_ ) );
NOR2_X1 _28820_ ( .A1(_06988_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07972_ ) );
AND4_X1 _28821_ ( .A1(_05952_ ), .A2(_06669_ ), .A3(_06589_ ), .A4(_06811_ ), .ZN(_07973_ ) );
NOR3_X1 _28822_ ( .A1(_07971_ ), .A2(_07972_ ), .A3(_07973_ ), .ZN(_07974_ ) );
OR2_X1 _28823_ ( .A1(_06676_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07975_ ) );
OR2_X1 _28824_ ( .A1(_06687_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07976_ ) );
NAND3_X1 _28825_ ( .A1(_07974_ ), .A2(_07975_ ), .A3(_07976_ ), .ZN(_07977_ ) );
NOR3_X1 _28826_ ( .A1(_06830_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06831_ ), .ZN(_07978_ ) );
AND4_X1 _28827_ ( .A1(_05958_ ), .A2(_06670_ ), .A3(_06834_ ), .A4(_11125_ ), .ZN(_07979_ ) );
NOR3_X1 _28828_ ( .A1(_07977_ ), .A2(_07978_ ), .A3(_07979_ ), .ZN(_07980_ ) );
NAND4_X1 _28829_ ( .A1(_07057_ ), .A2(_06835_ ), .A3(_05961_ ), .A4(_06741_ ), .ZN(_07981_ ) );
OR3_X1 _28830_ ( .A1(_06843_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06831_ ), .ZN(_07982_ ) );
AND3_X1 _28831_ ( .A1(_07980_ ), .A2(_07981_ ), .A3(_07982_ ), .ZN(_07983_ ) );
OR2_X1 _28832_ ( .A1(_06706_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07984_ ) );
NAND4_X1 _28833_ ( .A1(_06709_ ), .A2(_06711_ ), .A3(_05966_ ), .A4(_06852_ ), .ZN(_07985_ ) );
NAND3_X1 _28834_ ( .A1(_07983_ ), .A2(_07984_ ), .A3(_07985_ ), .ZN(_07986_ ) );
OAI21_X1 _28835_ ( .A(_06933_ ), .B1(_06717_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07987_ ) );
OAI21_X1 _28836_ ( .A(_07954_ ), .B1(_07986_ ), .B2(_07987_ ), .ZN(_07988_ ) );
NAND4_X1 _28837_ ( .A1(_06722_ ), .A2(_06727_ ), .A3(_05972_ ), .A4(_06728_ ), .ZN(_07989_ ) );
OR2_X1 _28838_ ( .A1(_06732_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07990_ ) );
NAND3_X1 _28839_ ( .A1(_07988_ ), .A2(_07989_ ), .A3(_07990_ ), .ZN(_07991_ ) );
NOR2_X1 _28840_ ( .A1(_06738_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07992_ ) );
AND4_X1 _28841_ ( .A1(_05977_ ), .A2(_06757_ ), .A3(_07067_ ), .A4(_01101_ ), .ZN(_07993_ ) );
NOR3_X1 _28842_ ( .A1(_07991_ ), .A2(_07992_ ), .A3(_07993_ ), .ZN(_07994_ ) );
AOI22_X1 _28843_ ( .A1(_06751_ ), .A2(_05980_ ), .B1(_01102_ ), .B2(_06745_ ), .ZN(_07995_ ) );
AOI22_X1 _28844_ ( .A1(_07994_ ), .A2(_07995_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06747_ ), .ZN(_07996_ ) );
OAI21_X1 _28845_ ( .A(_07953_ ), .B1(_07996_ ), .B2(_06598_ ), .ZN(_07997_ ) );
OAI211_X1 _28846_ ( .A(_07950_ ), .B(_07952_ ), .C1(_06584_ ), .C2(_07997_ ), .ZN(\idu.io_out_bits_rs2_data [2] ) );
AND3_X1 _28847_ ( .A1(_03334_ ), .A2(_03335_ ), .A3(_06766_ ), .ZN(_07998_ ) );
NOR3_X1 _28848_ ( .A1(_07195_ ), .A2(_00639_ ), .A3(_07196_ ), .ZN(_07999_ ) );
OAI22_X1 _28849_ ( .A1(\lsu.io_out_bits_rd_wdata [28] ), .A2(_07193_ ), .B1(_07194_ ), .B2(_07999_ ), .ZN(_08000_ ) );
AND4_X1 _28850_ ( .A1(_06045_ ), .A2(_06757_ ), .A3(_07067_ ), .A4(_06885_ ), .ZN(_08001_ ) );
AND3_X1 _28851_ ( .A1(_06730_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03834_ ), .ZN(_08002_ ) );
NAND3_X1 _28852_ ( .A1(_06703_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03833_ ), .ZN(_08003_ ) );
OR2_X1 _28853_ ( .A1(_07094_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08004_ ) );
OR3_X1 _28854_ ( .A1(_06828_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .A3(_11122_ ), .ZN(_08005_ ) );
OR3_X1 _28855_ ( .A1(_11127_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11122_ ), .ZN(_08006_ ) );
NAND3_X1 _28856_ ( .A1(_08004_ ), .A2(_08005_ ), .A3(_08006_ ), .ZN(_08007_ ) );
OAI21_X1 _28857_ ( .A(_06972_ ), .B1(_07264_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08008_ ) );
OAI21_X1 _28858_ ( .A(_08003_ ), .B1(_08007_ ), .B2(_08008_ ), .ZN(_08009_ ) );
NAND4_X1 _28859_ ( .A1(_07215_ ), .A2(_06697_ ), .A3(_06004_ ), .A4(_06815_ ), .ZN(_08010_ ) );
OR3_X1 _28860_ ( .A1(_06637_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11123_ ), .ZN(_08011_ ) );
NAND3_X1 _28861_ ( .A1(_08009_ ), .A2(_08010_ ), .A3(_08011_ ), .ZN(_08012_ ) );
NOR3_X1 _28862_ ( .A1(_06804_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11124_ ), .ZN(_08013_ ) );
NOR2_X1 _28863_ ( .A1(_08012_ ), .A2(_08013_ ), .ZN(_08014_ ) );
NOR2_X1 _28864_ ( .A1(_06647_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08015_ ) );
NOR2_X1 _28865_ ( .A1(_08015_ ), .A2(_06654_ ), .ZN(_08016_ ) );
AOI21_X1 _28866_ ( .A(_08002_ ), .B1(_08014_ ), .B2(_08016_ ), .ZN(_08017_ ) );
NOR2_X1 _28867_ ( .A1(_06809_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08018_ ) );
AND3_X1 _28868_ ( .A1(_06658_ ), .A2(_06014_ ), .A3(_06816_ ), .ZN(_08019_ ) );
NOR3_X1 _28869_ ( .A1(_08017_ ), .A2(_08018_ ), .A3(_08019_ ), .ZN(_08020_ ) );
NAND4_X1 _28870_ ( .A1(_06720_ ), .A2(_06910_ ), .A3(_06017_ ), .A4(_06846_ ), .ZN(_08021_ ) );
OR3_X1 _28871_ ( .A1(_07110_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06690_ ), .ZN(_08022_ ) );
NAND3_X1 _28872_ ( .A1(_08020_ ), .A2(_08021_ ), .A3(_08022_ ), .ZN(_08023_ ) );
NOR2_X1 _28873_ ( .A1(_06677_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08024_ ) );
NOR2_X1 _28874_ ( .A1(_06824_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08025_ ) );
NOR3_X1 _28875_ ( .A1(_08023_ ), .A2(_08024_ ), .A3(_08025_ ), .ZN(_08026_ ) );
OR3_X1 _28876_ ( .A1(_06830_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07199_ ), .ZN(_08027_ ) );
NAND4_X1 _28877_ ( .A1(_06708_ ), .A2(_06916_ ), .A3(_06024_ ), .A4(_06596_ ), .ZN(_08028_ ) );
NAND3_X1 _28878_ ( .A1(_08026_ ), .A2(_08027_ ), .A3(_08028_ ), .ZN(_08029_ ) );
NOR2_X1 _28879_ ( .A1(_06841_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08030_ ) );
NOR3_X1 _28880_ ( .A1(_06844_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06847_ ), .ZN(_08031_ ) );
NOR3_X1 _28881_ ( .A1(_08029_ ), .A2(_08030_ ), .A3(_08031_ ), .ZN(_08032_ ) );
NAND4_X1 _28882_ ( .A1(_06850_ ), .A2(_07232_ ), .A3(_06030_ ), .A4(_06865_ ), .ZN(_08033_ ) );
NAND4_X1 _28883_ ( .A1(_06709_ ), .A2(_07232_ ), .A3(_06032_ ), .A4(_06865_ ), .ZN(_08034_ ) );
NAND3_X1 _28884_ ( .A1(_08032_ ), .A2(_08033_ ), .A3(_08034_ ), .ZN(_08035_ ) );
NOR3_X1 _28885_ ( .A1(_06855_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07007_ ), .ZN(_08036_ ) );
NOR3_X1 _28886_ ( .A1(_07006_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06856_ ), .ZN(_08037_ ) );
NOR3_X1 _28887_ ( .A1(_08035_ ), .A2(_08036_ ), .A3(_08037_ ), .ZN(_08038_ ) );
NAND4_X1 _28888_ ( .A1(_06947_ ), .A2(_07071_ ), .A3(_06038_ ), .A4(_06866_ ), .ZN(_08039_ ) );
AOI22_X1 _28889_ ( .A1(_06731_ ), .A2(_06040_ ), .B1(_06885_ ), .B2(_06735_ ), .ZN(_08040_ ) );
NAND3_X1 _28890_ ( .A1(_08038_ ), .A2(_08039_ ), .A3(_08040_ ), .ZN(_08041_ ) );
NAND3_X1 _28891_ ( .A1(_06735_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01102_ ), .ZN(_08042_ ) );
AOI21_X1 _28892_ ( .A(_08001_ ), .B1(_08041_ ), .B2(_08042_ ), .ZN(_08043_ ) );
OR2_X1 _28893_ ( .A1(_06752_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08044_ ) );
NOR3_X1 _28894_ ( .A1(_07188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03838_ ), .ZN(_08045_ ) );
NOR2_X1 _28895_ ( .A1(_08045_ ), .A2(_06598_ ), .ZN(_08046_ ) );
AND3_X1 _28896_ ( .A1(_08043_ ), .A2(_08044_ ), .A3(_08046_ ), .ZN(_08047_ ) );
NAND3_X1 _28897_ ( .A1(_06953_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_06950_ ), .ZN(_08048_ ) );
NAND4_X1 _28898_ ( .A1(_07248_ ), .A2(_07249_ ), .A3(_06876_ ), .A4(_08048_ ), .ZN(_08049_ ) );
OAI22_X1 _28899_ ( .A1(_07998_ ), .A2(_08000_ ), .B1(_08047_ ), .B2(_08049_ ), .ZN(\idu.io_out_bits_rs2_data [28] ) );
NOR2_X1 _28900_ ( .A1(\exu.io_out_bits_rd_wdata [1] ), .A2(_06957_ ), .ZN(_08050_ ) );
NOR3_X1 _28901_ ( .A1(_07195_ ), .A2(_00640_ ), .A3(_07196_ ), .ZN(_08051_ ) );
OAI22_X1 _28902_ ( .A1(\lsu.io_out_bits_rd_wdata [1] ), .A2(_07193_ ), .B1(_07194_ ), .B2(_08051_ ), .ZN(_08052_ ) );
NOR2_X1 _28903_ ( .A1(_06738_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08053_ ) );
NOR3_X1 _28904_ ( .A1(_06802_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06856_ ), .ZN(_08054_ ) );
AND4_X1 _28905_ ( .A1(_06067_ ), .A2(_06720_ ), .A3(_06834_ ), .A4(_11125_ ), .ZN(_08055_ ) );
NAND3_X1 _28906_ ( .A1(_10651_ ), .A2(_06071_ ), .A3(_11050_ ), .ZN(_08056_ ) );
OAI21_X1 _28907_ ( .A(_08056_ ), .B1(_10688_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08057_ ) );
AOI21_X1 _28908_ ( .A(_08057_ ), .B1(_06075_ ), .B2(_06619_ ), .ZN(_08058_ ) );
OR3_X1 _28909_ ( .A1(_06625_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_10812_ ), .ZN(_08059_ ) );
NAND4_X1 _28910_ ( .A1(_06627_ ), .A2(_06628_ ), .A3(_06078_ ), .A4(_06673_ ), .ZN(_08060_ ) );
AND3_X1 _28911_ ( .A1(_08058_ ), .A2(_08059_ ), .A3(_08060_ ), .ZN(_08061_ ) );
OR2_X1 _28912_ ( .A1(_06799_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08062_ ) );
NAND4_X1 _28913_ ( .A1(_06897_ ), .A2(_06696_ ), .A3(_06082_ ), .A4(_06814_ ), .ZN(_08063_ ) );
NAND3_X1 _28914_ ( .A1(_08061_ ), .A2(_08062_ ), .A3(_08063_ ), .ZN(_08064_ ) );
NOR3_X1 _28915_ ( .A1(_06641_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11123_ ), .ZN(_08065_ ) );
AND4_X1 _28916_ ( .A1(_06086_ ), .A2(_06627_ ), .A3(_06723_ ), .A4(_06796_ ), .ZN(_08066_ ) );
NOR3_X1 _28917_ ( .A1(_08064_ ), .A2(_08065_ ), .A3(_08066_ ), .ZN(_08067_ ) );
OR2_X1 _28918_ ( .A1(_06655_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08068_ ) );
OR2_X1 _28919_ ( .A1(_06650_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08069_ ) );
AND3_X1 _28920_ ( .A1(_08067_ ), .A2(_08068_ ), .A3(_08069_ ), .ZN(_08070_ ) );
OR2_X1 _28921_ ( .A1(_07106_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08071_ ) );
NAND4_X1 _28922_ ( .A1(_06665_ ), .A2(_06909_ ), .A3(_06092_ ), .A4(_06811_ ), .ZN(_08072_ ) );
NAND3_X1 _28923_ ( .A1(_08070_ ), .A2(_08071_ ), .A3(_08072_ ), .ZN(_08073_ ) );
NOR3_X1 _28924_ ( .A1(_07110_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06690_ ), .ZN(_08074_ ) );
OAI21_X1 _28925_ ( .A(_06686_ ), .B1(_06676_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08075_ ) );
OR3_X1 _28926_ ( .A1(_08073_ ), .A2(_08074_ ), .A3(_08075_ ), .ZN(_08076_ ) );
NAND3_X1 _28927_ ( .A1(_06684_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06605_ ), .ZN(_08077_ ) );
AOI21_X1 _28928_ ( .A(_08055_ ), .B1(_08076_ ), .B2(_08077_ ), .ZN(_08078_ ) );
OR3_X1 _28929_ ( .A1(_06918_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06831_ ), .ZN(_08079_ ) );
OR2_X1 _28930_ ( .A1(_06840_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08080_ ) );
AND3_X1 _28931_ ( .A1(_08078_ ), .A2(_08079_ ), .A3(_08080_ ), .ZN(_08081_ ) );
NAND4_X1 _28932_ ( .A1(_06711_ ), .A2(_07066_ ), .A3(_06103_ ), .A4(_06852_ ), .ZN(_08082_ ) );
AOI22_X1 _28933_ ( .A1(_06704_ ), .A2(_06105_ ), .B1(_01100_ ), .B2(_06631_ ), .ZN(_08083_ ) );
NAND3_X1 _28934_ ( .A1(_08081_ ), .A2(_08082_ ), .A3(_08083_ ), .ZN(_08084_ ) );
NAND3_X1 _28935_ ( .A1(_06631_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06607_ ), .ZN(_08085_ ) );
AOI21_X1 _28936_ ( .A(_08054_ ), .B1(_08084_ ), .B2(_08085_ ), .ZN(_08086_ ) );
NAND3_X1 _28937_ ( .A1(_06604_ ), .A2(_06110_ ), .A3(_06885_ ), .ZN(_08087_ ) );
NAND4_X1 _28938_ ( .A1(_06722_ ), .A2(_06727_ ), .A3(_06112_ ), .A4(_06728_ ), .ZN(_08088_ ) );
NAND4_X1 _28939_ ( .A1(_08086_ ), .A2(_06940_ ), .A3(_08087_ ), .A4(_08088_ ), .ZN(_08089_ ) );
NAND4_X1 _28940_ ( .A1(_06756_ ), .A2(_06937_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_01102_ ), .ZN(_08090_ ) );
AOI21_X1 _28941_ ( .A(_08053_ ), .B1(_08089_ ), .B2(_08090_ ), .ZN(_08091_ ) );
NAND4_X1 _28942_ ( .A1(_06758_ ), .A2(_07067_ ), .A3(_06117_ ), .A4(_07018_ ), .ZN(_08092_ ) );
OR2_X1 _28943_ ( .A1(_06752_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08093_ ) );
NAND3_X1 _28944_ ( .A1(_08091_ ), .A2(_08092_ ), .A3(_08093_ ), .ZN(_08094_ ) );
NOR3_X1 _28945_ ( .A1(_07188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03838_ ), .ZN(_08095_ ) );
NOR3_X1 _28946_ ( .A1(_08094_ ), .A2(_06598_ ), .A3(_08095_ ), .ZN(_08096_ ) );
NAND3_X1 _28947_ ( .A1(_06953_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_06950_ ), .ZN(_08097_ ) );
NAND4_X1 _28948_ ( .A1(_07248_ ), .A2(_06773_ ), .A3(_06876_ ), .A4(_08097_ ), .ZN(_08098_ ) );
OAI22_X1 _28949_ ( .A1(_08050_ ), .A2(_08052_ ), .B1(_08096_ ), .B2(_08098_ ), .ZN(\idu.io_out_bits_rs2_data [1] ) );
NAND2_X1 _28950_ ( .A1(\exu.io_out_bits_rd_wdata [0] ), .A2(_06767_ ), .ZN(_08099_ ) );
AND4_X1 _28951_ ( .A1(_06565_ ), .A2(_06570_ ), .A3(_06573_ ), .A4(_06572_ ), .ZN(_08100_ ) );
NAND4_X1 _28952_ ( .A1(_08100_ ), .A2(_06566_ ), .A3(_06567_ ), .A4(_06571_ ), .ZN(_08101_ ) );
AOI21_X1 _28953_ ( .A(_08101_ ), .B1(_03966_ ), .B2(_03988_ ), .ZN(_08102_ ) );
NAND4_X1 _28954_ ( .A1(_06562_ ), .A2(_04235_ ), .A3(_06563_ ), .A4(_06569_ ), .ZN(_08103_ ) );
NOR2_X1 _28955_ ( .A1(_13276_ ), .A2(_08103_ ), .ZN(_08104_ ) );
NAND3_X1 _28956_ ( .A1(_08102_ ), .A2(\wbu.io_in_bits_rd_wdata [0] ), .A3(_08104_ ), .ZN(_08105_ ) );
OAI211_X1 _28957_ ( .A(_10786_ ), .B(_10755_ ), .C1(_03920_ ), .C2(_03922_ ), .ZN(_08106_ ) );
NOR2_X1 _28958_ ( .A1(_04657_ ), .A2(_08106_ ), .ZN(_08107_ ) );
MUX2_X1 _28959_ ( .A(_08105_ ), .B(_06161_ ), .S(_08107_ ), .Z(_08108_ ) );
AND3_X1 _28960_ ( .A1(_06730_ ), .A2(\wbu.rf_10 [0] ), .A3(_06847_ ), .ZN(_08109_ ) );
AND3_X1 _28961_ ( .A1(_06635_ ), .A2(\wbu.rf_7 [0] ), .A3(_03836_ ), .ZN(_08110_ ) );
OR2_X1 _28962_ ( .A1(_08109_ ), .A2(_08110_ ), .ZN(_08111_ ) );
AOI221_X4 _28963_ ( .A(_08111_ ), .B1(\wbu.rf_29 [0] ), .B2(_06751_ ), .C1(\wbu.rf_5 [0] ), .C2(_06970_ ), .ZN(_08112_ ) );
AND3_X1 _28964_ ( .A1(_06749_ ), .A2(\wbu.rf_13 [0] ), .A3(_03836_ ), .ZN(_08113_ ) );
AND3_X1 _28965_ ( .A1(_06604_ ), .A2(\wbu.rf_8 [0] ), .A3(_03836_ ), .ZN(_08114_ ) );
OR2_X1 _28966_ ( .A1(_08113_ ), .A2(_08114_ ), .ZN(_08115_ ) );
AOI221_X4 _28967_ ( .A(_08115_ ), .B1(\wbu.rf_25 [0] ), .B2(_06859_ ), .C1(\wbu.rf_6 [0] ), .C2(_06632_ ), .ZN(_08116_ ) );
AND3_X1 _28968_ ( .A1(_06966_ ), .A2(\wbu.rf_2 [0] ), .A3(_03836_ ), .ZN(_08117_ ) );
AND3_X1 _28969_ ( .A1(_06684_ ), .A2(\wbu.rf_16 [0] ), .A3(_06605_ ), .ZN(_08118_ ) );
OR2_X1 _28970_ ( .A1(_08117_ ), .A2(_08118_ ), .ZN(_08119_ ) );
AOI221_X4 _28971_ ( .A(_08119_ ), .B1(\wbu.rf_19 [0] ), .B2(_06838_ ), .C1(\wbu.rf_14 [0] ), .C2(_06819_ ), .ZN(_08120_ ) );
NAND3_X1 _28972_ ( .A1(_06735_ ), .A2(\wbu.rf_27 [0] ), .A3(_01100_ ), .ZN(_08121_ ) );
NAND3_X1 _28973_ ( .A1(_06740_ ), .A2(\wbu.rf_28 [0] ), .A3(_06606_ ), .ZN(_08122_ ) );
NAND2_X1 _28974_ ( .A1(_08121_ ), .A2(_08122_ ), .ZN(_08123_ ) );
AOI221_X4 _28975_ ( .A(_08123_ ), .B1(\wbu.rf_22 [0] ), .B2(_06928_ ), .C1(\wbu._GEN_71 [0] ), .C2(_10652_ ), .ZN(_08124_ ) );
NAND4_X1 _28976_ ( .A1(_08112_ ), .A2(_08116_ ), .A3(_08120_ ), .A4(_08124_ ), .ZN(_08125_ ) );
AOI22_X1 _28977_ ( .A1(\wbu.rf_30 [0] ), .A2(_06747_ ), .B1(_06731_ ), .B2(\wbu.rf_26 [0] ), .ZN(_08126_ ) );
AOI22_X1 _28978_ ( .A1(\wbu.rf_18 [0] ), .A2(_07055_ ), .B1(_06619_ ), .B2(\wbu.rf_3 [0] ), .ZN(_08127_ ) );
AOI22_X1 _28979_ ( .A1(\wbu.rf_23 [0] ), .A2(_06716_ ), .B1(_07263_ ), .B2(\wbu.rf_4 [0] ), .ZN(_08128_ ) );
AND3_X1 _28980_ ( .A1(_06679_ ), .A2(\wbu.rf_17 [0] ), .A3(_01101_ ), .ZN(_08129_ ) );
AOI21_X1 _28981_ ( .A(_08129_ ), .B1(\wbu.rf_24 [0] ), .B2(_06714_ ), .ZN(_08130_ ) );
NAND4_X1 _28982_ ( .A1(_08126_ ), .A2(_08127_ ), .A3(_08128_ ), .A4(_08130_ ), .ZN(_08131_ ) );
AND3_X1 _28983_ ( .A1(_06858_ ), .A2(\wbu.rf_9 [0] ), .A3(_03837_ ), .ZN(_08132_ ) );
AOI221_X4 _28984_ ( .A(_08132_ ), .B1(_06675_ ), .B2(\wbu.rf_15 [0] ), .C1(\wbu.rf_12 [0] ), .C2(_06659_ ), .ZN(_08133_ ) );
AOI22_X1 _28985_ ( .A1(\wbu.rf_21 [0] ), .A2(_06704_ ), .B1(_06922_ ), .B2(\wbu.rf_20 [0] ), .ZN(_08134_ ) );
AND3_X1 _28986_ ( .A1(_06591_ ), .A2(\wbu.rf_31 [0] ), .A3(_01101_ ), .ZN(_08135_ ) );
AOI21_X1 _28987_ ( .A(_08135_ ), .B1(\wbu.rf_11 [0] ), .B2(_06649_ ), .ZN(_08136_ ) );
NAND3_X1 _28988_ ( .A1(_08133_ ), .A2(_08134_ ), .A3(_08136_ ), .ZN(_08137_ ) );
NOR3_X1 _28989_ ( .A1(_08125_ ), .A2(_08131_ ), .A3(_08137_ ), .ZN(_08138_ ) );
OAI221_X1 _28990_ ( .A(_08099_ ), .B1(_06879_ ), .B2(_08108_ ), .C1(_06584_ ), .C2(_08138_ ), .ZN(\idu.io_out_bits_rs2_data [0] ) );
OAI21_X1 _28991_ ( .A(_06767_ ), .B1(_03581_ ), .B2(_03582_ ), .ZN(_08139_ ) );
OAI21_X1 _28992_ ( .A(_08107_ ), .B1(_06164_ ), .B2(_06165_ ), .ZN(_08140_ ) );
AND3_X1 _28993_ ( .A1(_08102_ ), .A2(\wbu.io_in_bits_rd_wdata [27] ), .A3(_08104_ ), .ZN(_08141_ ) );
OAI211_X1 _28994_ ( .A(_08140_ ), .B(_07249_ ), .C1(_08107_ ), .C2(_08141_ ), .ZN(_08142_ ) );
AND3_X1 _28995_ ( .A1(_06603_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11052_ ), .ZN(_08143_ ) );
NOR2_X1 _28996_ ( .A1(_06633_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08144_ ) );
NAND3_X1 _28997_ ( .A1(_10651_ ), .A2(_06177_ ), .A3(_10621_ ), .ZN(_08145_ ) );
MUX2_X1 _28998_ ( .A(_08145_ ), .B(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(_10687_ ), .Z(_08146_ ) );
MUX2_X1 _28999_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_08146_ ), .S(_06620_ ), .Z(_08147_ ) );
MUX2_X1 _29000_ ( .A(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_08147_ ), .S(_07264_ ), .Z(_08148_ ) );
NAND2_X1 _29001_ ( .A1(_08148_ ), .A2(_06972_ ), .ZN(_08149_ ) );
NAND4_X1 _29002_ ( .A1(_06627_ ), .A2(_06628_ ), .A3(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A4(_03832_ ), .ZN(_08150_ ) );
AOI21_X1 _29003_ ( .A(_08144_ ), .B1(_08149_ ), .B2(_08150_ ), .ZN(_08151_ ) );
NOR3_X1 _29004_ ( .A1(_06637_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06592_ ), .ZN(_08152_ ) );
NOR2_X1 _29005_ ( .A1(_08152_ ), .A2(_07152_ ), .ZN(_08153_ ) );
AOI21_X1 _29006_ ( .A(_08143_ ), .B1(_08151_ ), .B2(_08153_ ), .ZN(_08154_ ) );
NOR2_X1 _29007_ ( .A1(_06646_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08155_ ) );
AND3_X1 _29008_ ( .A1(_06652_ ), .A2(_06189_ ), .A3(_06674_ ), .ZN(_08156_ ) );
NOR3_X1 _29009_ ( .A1(_08154_ ), .A2(_08155_ ), .A3(_08156_ ), .ZN(_08157_ ) );
NAND4_X1 _29010_ ( .A1(_06898_ ), .A2(_06724_ ), .A3(_06192_ ), .A4(_06610_ ), .ZN(_08158_ ) );
OR2_X1 _29011_ ( .A1(_06660_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08159_ ) );
AND3_X1 _29012_ ( .A1(_08157_ ), .A2(_08158_ ), .A3(_08159_ ), .ZN(_08160_ ) );
NAND4_X1 _29013_ ( .A1(_06665_ ), .A2(_06909_ ), .A3(_06196_ ), .A4(_06845_ ), .ZN(_08161_ ) );
NAND4_X1 _29014_ ( .A1(_06669_ ), .A2(_06909_ ), .A3(_06198_ ), .A4(_06845_ ), .ZN(_08162_ ) );
NAND3_X1 _29015_ ( .A1(_08160_ ), .A2(_08161_ ), .A3(_08162_ ), .ZN(_08163_ ) );
NOR2_X1 _29016_ ( .A1(_06676_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08164_ ) );
NOR2_X1 _29017_ ( .A1(_06686_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08165_ ) );
NOR3_X1 _29018_ ( .A1(_08163_ ), .A2(_08164_ ), .A3(_08165_ ), .ZN(_08166_ ) );
OR3_X1 _29019_ ( .A1(_06829_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03835_ ), .ZN(_08167_ ) );
OR3_X1 _29020_ ( .A1(_11127_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03835_ ), .ZN(_08168_ ) );
NAND3_X1 _29021_ ( .A1(_08166_ ), .A2(_08167_ ), .A3(_08168_ ), .ZN(_08169_ ) );
NOR2_X1 _29022_ ( .A1(_06840_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08170_ ) );
NOR3_X1 _29023_ ( .A1(_06843_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07199_ ), .ZN(_08171_ ) );
NOR3_X1 _29024_ ( .A1(_08169_ ), .A2(_08170_ ), .A3(_08171_ ), .ZN(_08172_ ) );
OR2_X1 _29025_ ( .A1(_06705_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08173_ ) );
AND3_X1 _29026_ ( .A1(_08172_ ), .A2(_06930_ ), .A3(_08173_ ), .ZN(_08174_ ) );
AOI21_X1 _29027_ ( .A(_08174_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06928_ ), .ZN(_08175_ ) );
NOR3_X1 _29028_ ( .A1(_06855_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07007_ ), .ZN(_08176_ ) );
NOR3_X1 _29029_ ( .A1(_07006_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07007_ ), .ZN(_08177_ ) );
NOR3_X1 _29030_ ( .A1(_08175_ ), .A2(_08176_ ), .A3(_08177_ ), .ZN(_08178_ ) );
NAND4_X1 _29031_ ( .A1(_06947_ ), .A2(_07010_ ), .A3(_06212_ ), .A4(_07011_ ), .ZN(_08179_ ) );
NAND4_X1 _29032_ ( .A1(_06756_ ), .A2(_07071_ ), .A3(_06215_ ), .A4(_06866_ ), .ZN(_08180_ ) );
AND3_X1 _29033_ ( .A1(_08178_ ), .A2(_08179_ ), .A3(_08180_ ), .ZN(_08181_ ) );
OR2_X1 _29034_ ( .A1(_06944_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08182_ ) );
OR2_X1 _29035_ ( .A1(_06943_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08183_ ) );
NAND3_X1 _29036_ ( .A1(_08181_ ), .A2(_08182_ ), .A3(_08183_ ), .ZN(_08184_ ) );
AND4_X1 _29037_ ( .A1(_06220_ ), .A2(_06936_ ), .A3(_06758_ ), .A4(_06883_ ), .ZN(_08185_ ) );
OAI21_X1 _29038_ ( .A(_07134_ ), .B1(_06872_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08186_ ) );
NOR3_X1 _29039_ ( .A1(_08184_ ), .A2(_08185_ ), .A3(_08186_ ), .ZN(_08187_ ) );
NAND3_X1 _29040_ ( .A1(_07251_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_07080_ ), .ZN(_08188_ ) );
NAND4_X1 _29041_ ( .A1(_07248_ ), .A2(_07249_ ), .A3(_07250_ ), .A4(_08188_ ), .ZN(_08189_ ) );
OAI211_X1 _29042_ ( .A(_08139_ ), .B(_08142_ ), .C1(_08187_ ), .C2(_08189_ ), .ZN(\idu.io_out_bits_rs2_data [27] ) );
AND3_X1 _29043_ ( .A1(_03628_ ), .A2(_03629_ ), .A3(_06766_ ), .ZN(_08190_ ) );
NOR3_X1 _29044_ ( .A1(_07195_ ), .A2(_00808_ ), .A3(_07196_ ), .ZN(_08191_ ) );
OAI22_X1 _29045_ ( .A1(\lsu.io_out_bits_rd_wdata [26] ), .A2(_07193_ ), .B1(_07194_ ), .B2(_08191_ ), .ZN(_08192_ ) );
NAND3_X1 _29046_ ( .A1(_06761_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(\idu.immI [4] ), .ZN(_08193_ ) );
NOR2_X1 _29047_ ( .A1(_06687_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08194_ ) );
NAND3_X1 _29048_ ( .A1(_06679_ ), .A2(_06235_ ), .A3(_11052_ ), .ZN(_08195_ ) );
OAI21_X1 _29049_ ( .A(_08195_ ), .B1(_10688_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08196_ ) );
AND4_X1 _29050_ ( .A1(_06239_ ), .A2(_06587_ ), .A3(_06833_ ), .A4(_03832_ ), .ZN(_08197_ ) );
NOR3_X1 _29051_ ( .A1(_06794_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06638_ ), .ZN(_08198_ ) );
NOR3_X1 _29052_ ( .A1(_08196_ ), .A2(_08197_ ), .A3(_08198_ ), .ZN(_08199_ ) );
NAND4_X1 _29053_ ( .A1(_06663_ ), .A2(_07210_ ), .A3(_06242_ ), .A4(_03833_ ), .ZN(_08200_ ) );
OR2_X1 _29054_ ( .A1(_06799_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08201_ ) );
NAND3_X1 _29055_ ( .A1(_08199_ ), .A2(_08200_ ), .A3(_08201_ ), .ZN(_08202_ ) );
AND4_X1 _29056_ ( .A1(_06246_ ), .A2(_06897_ ), .A3(_07210_ ), .A4(_03833_ ), .ZN(_08203_ ) );
NOR3_X1 _29057_ ( .A1(_06804_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06593_ ), .ZN(_08204_ ) );
NOR3_X1 _29058_ ( .A1(_08202_ ), .A2(_08203_ ), .A3(_08204_ ), .ZN(_08205_ ) );
NAND4_X1 _29059_ ( .A1(_06664_ ), .A2(_06724_ ), .A3(_06250_ ), .A4(_03834_ ), .ZN(_08206_ ) );
NAND4_X1 _29060_ ( .A1(_06669_ ), .A2(_06724_ ), .A3(_06252_ ), .A4(_03834_ ), .ZN(_08207_ ) );
NAND3_X1 _29061_ ( .A1(_08205_ ), .A2(_08206_ ), .A3(_08207_ ), .ZN(_08208_ ) );
NOR2_X1 _29062_ ( .A1(_06809_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08209_ ) );
NOR2_X1 _29063_ ( .A1(_06661_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08210_ ) );
NOR3_X1 _29064_ ( .A1(_08208_ ), .A2(_08209_ ), .A3(_08210_ ), .ZN(_08211_ ) );
NAND4_X1 _29065_ ( .A1(_06665_ ), .A2(_06666_ ), .A3(_06258_ ), .A4(_03835_ ), .ZN(_08212_ ) );
AOI22_X1 _29066_ ( .A1(_06819_ ), .A2(_06260_ ), .B1(_03835_ ), .B2(_06590_ ), .ZN(_08213_ ) );
NAND3_X1 _29067_ ( .A1(_08211_ ), .A2(_08212_ ), .A3(_08213_ ), .ZN(_08214_ ) );
NAND3_X1 _29068_ ( .A1(_06590_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06831_ ), .ZN(_08215_ ) );
AOI21_X1 _29069_ ( .A(_08194_ ), .B1(_08214_ ), .B2(_08215_ ), .ZN(_08216_ ) );
OR3_X1 _29070_ ( .A1(_06829_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06612_ ), .ZN(_08217_ ) );
NAND4_X1 _29071_ ( .A1(_06708_ ), .A2(_06835_ ), .A3(_06267_ ), .A4(_01099_ ), .ZN(_08218_ ) );
NAND3_X1 _29072_ ( .A1(_08216_ ), .A2(_08217_ ), .A3(_08218_ ), .ZN(_08219_ ) );
NOR2_X1 _29073_ ( .A1(_06841_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08220_ ) );
NOR3_X1 _29074_ ( .A1(_06844_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06847_ ), .ZN(_08221_ ) );
NOR3_X1 _29075_ ( .A1(_08219_ ), .A2(_08220_ ), .A3(_08221_ ), .ZN(_08222_ ) );
NAND4_X1 _29076_ ( .A1(_06850_ ), .A2(_06710_ ), .A3(_06273_ ), .A4(_01100_ ), .ZN(_08223_ ) );
NAND4_X1 _29077_ ( .A1(_06708_ ), .A2(_06710_ ), .A3(_06275_ ), .A4(_01100_ ), .ZN(_08224_ ) );
NAND3_X1 _29078_ ( .A1(_08222_ ), .A2(_08223_ ), .A3(_08224_ ), .ZN(_08225_ ) );
NOR3_X1 _29079_ ( .A1(_06802_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06856_ ), .ZN(_08226_ ) );
NOR3_X1 _29080_ ( .A1(_06804_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03837_ ), .ZN(_08227_ ) );
NOR3_X1 _29081_ ( .A1(_08225_ ), .A2(_08226_ ), .A3(_08227_ ), .ZN(_08228_ ) );
NAND4_X1 _29082_ ( .A1(_06722_ ), .A2(_06727_ ), .A3(_06281_ ), .A4(_06728_ ), .ZN(_08229_ ) );
OR2_X1 _29083_ ( .A1(_06732_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08230_ ) );
NAND3_X1 _29084_ ( .A1(_08228_ ), .A2(_08229_ ), .A3(_08230_ ), .ZN(_08231_ ) );
NOR2_X1 _29085_ ( .A1(_06738_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08232_ ) );
NOR2_X1 _29086_ ( .A1(_06743_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08233_ ) );
NOR3_X1 _29087_ ( .A1(_08231_ ), .A2(_08232_ ), .A3(_08233_ ), .ZN(_08234_ ) );
OAI21_X1 _29088_ ( .A(_08234_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06870_ ), .ZN(_08235_ ) );
OAI21_X1 _29089_ ( .A(_07134_ ), .B1(_06748_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08236_ ) );
OAI21_X1 _29090_ ( .A(_08193_ ), .B1(_08235_ ), .B2(_08236_ ), .ZN(_08237_ ) );
OAI22_X1 _29091_ ( .A1(_08190_ ), .A2(_08192_ ), .B1(_06584_ ), .B2(_08237_ ), .ZN(\idu.io_out_bits_rs2_data [26] ) );
AND3_X1 _29092_ ( .A1(_03676_ ), .A2(_03677_ ), .A3(_06766_ ), .ZN(_08238_ ) );
NOR3_X1 _29093_ ( .A1(_07195_ ), .A2(_00845_ ), .A3(_07196_ ), .ZN(_08239_ ) );
OAI22_X1 _29094_ ( .A1(\lsu.io_out_bits_rd_wdata [25] ), .A2(_07193_ ), .B1(_07194_ ), .B2(_08239_ ), .ZN(_08240_ ) );
NAND3_X1 _29095_ ( .A1(_06604_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06728_ ), .ZN(_08241_ ) );
AND4_X1 _29096_ ( .A1(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A2(_06723_ ), .A3(_06683_ ), .A4(_06609_ ), .ZN(_08242_ ) );
AND4_X1 _29097_ ( .A1(_06305_ ), .A2(_06668_ ), .A3(_06696_ ), .A4(_06796_ ), .ZN(_08243_ ) );
NAND3_X1 _29098_ ( .A1(_06966_ ), .A2(_06307_ ), .A3(_11050_ ), .ZN(_08244_ ) );
OAI21_X1 _29099_ ( .A(_08244_ ), .B1(_06791_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_08245_ ) );
MUX2_X1 _29100_ ( .A(_06311_ ), .B(_08245_ ), .S(_07094_ ), .Z(_08246_ ) );
NOR3_X1 _29101_ ( .A1(_06794_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11122_ ), .ZN(_08247_ ) );
OR3_X1 _29102_ ( .A1(_08246_ ), .A2(_06970_ ), .A3(_08247_ ), .ZN(_08248_ ) );
NAND3_X1 _29103_ ( .A1(_06703_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03833_ ), .ZN(_08249_ ) );
AOI21_X1 _29104_ ( .A(_08243_ ), .B1(_08248_ ), .B2(_08249_ ), .ZN(_08250_ ) );
OR3_X1 _29105_ ( .A1(_06637_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06638_ ), .ZN(_08251_ ) );
AND2_X1 _29106_ ( .A1(_08251_ ), .A2(_07153_ ), .ZN(_08252_ ) );
AOI21_X1 _29107_ ( .A(_08242_ ), .B1(_08250_ ), .B2(_08252_ ), .ZN(_08253_ ) );
NOR2_X1 _29108_ ( .A1(_06647_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08254_ ) );
AND4_X1 _29109_ ( .A1(_06320_ ), .A2(_07215_ ), .A3(_07156_ ), .A4(_07258_ ), .ZN(_08255_ ) );
NOR3_X1 _29110_ ( .A1(_08253_ ), .A2(_08254_ ), .A3(_08255_ ), .ZN(_08256_ ) );
NAND4_X1 _29111_ ( .A1(_06898_ ), .A2(_06725_ ), .A3(_06322_ ), .A4(_06611_ ), .ZN(_08257_ ) );
OR2_X1 _29112_ ( .A1(_06661_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08258_ ) );
NAND3_X1 _29113_ ( .A1(_08256_ ), .A2(_08257_ ), .A3(_08258_ ), .ZN(_08259_ ) );
NOR2_X1 _29114_ ( .A1(_06988_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08260_ ) );
AND4_X1 _29115_ ( .A1(_06327_ ), .A2(_06669_ ), .A3(_06909_ ), .A4(_06816_ ), .ZN(_08261_ ) );
NOR3_X1 _29116_ ( .A1(_08259_ ), .A2(_08260_ ), .A3(_08261_ ), .ZN(_08262_ ) );
NAND4_X1 _29117_ ( .A1(_07057_ ), .A2(_06757_ ), .A3(_06329_ ), .A4(_06831_ ), .ZN(_08263_ ) );
OR2_X1 _29118_ ( .A1(_06687_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08264_ ) );
NAND3_X1 _29119_ ( .A1(_08262_ ), .A2(_08263_ ), .A3(_08264_ ), .ZN(_08265_ ) );
NOR3_X1 _29120_ ( .A1(_06830_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06919_ ), .ZN(_08266_ ) );
AND4_X1 _29121_ ( .A1(_06334_ ), .A2(_06670_ ), .A3(_06834_ ), .A4(_06595_ ), .ZN(_08267_ ) );
NOR3_X1 _29122_ ( .A1(_08265_ ), .A2(_08266_ ), .A3(_08267_ ), .ZN(_08268_ ) );
NAND4_X1 _29123_ ( .A1(_07058_ ), .A2(_06916_ ), .A3(_06336_ ), .A4(_06750_ ), .ZN(_08269_ ) );
OR3_X1 _29124_ ( .A1(_06843_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06919_ ), .ZN(_08270_ ) );
AND3_X1 _29125_ ( .A1(_08268_ ), .A2(_08269_ ), .A3(_08270_ ), .ZN(_08271_ ) );
OR2_X1 _29126_ ( .A1(_06706_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08272_ ) );
NAND4_X1 _29127_ ( .A1(_06709_ ), .A2(_07232_ ), .A3(_06342_ ), .A4(_06865_ ), .ZN(_08273_ ) );
NAND3_X1 _29128_ ( .A1(_08271_ ), .A2(_08272_ ), .A3(_08273_ ), .ZN(_08274_ ) );
OAI21_X1 _29129_ ( .A(_06933_ ), .B1(_06717_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08275_ ) );
OAI21_X1 _29130_ ( .A(_08241_ ), .B1(_08274_ ), .B2(_08275_ ), .ZN(_08276_ ) );
NAND4_X1 _29131_ ( .A1(_06947_ ), .A2(_07071_ ), .A3(_06347_ ), .A4(_06866_ ), .ZN(_08277_ ) );
OR2_X1 _29132_ ( .A1(_06732_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08278_ ) );
AND3_X1 _29133_ ( .A1(_08276_ ), .A2(_08277_ ), .A3(_08278_ ), .ZN(_08279_ ) );
NAND4_X1 _29134_ ( .A1(_07058_ ), .A2(_06937_ ), .A3(_06351_ ), .A4(_07018_ ), .ZN(_08280_ ) );
OR2_X1 _29135_ ( .A1(_06743_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08281_ ) );
NAND3_X1 _29136_ ( .A1(_08279_ ), .A2(_08280_ ), .A3(_08281_ ), .ZN(_08282_ ) );
AND4_X1 _29137_ ( .A1(_06355_ ), .A2(_06936_ ), .A3(_06758_ ), .A4(_06883_ ), .ZN(_08283_ ) );
OAI21_X1 _29138_ ( .A(_07134_ ), .B1(_06748_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08284_ ) );
NOR3_X1 _29139_ ( .A1(_08282_ ), .A2(_08283_ ), .A3(_08284_ ), .ZN(_08285_ ) );
NAND3_X1 _29140_ ( .A1(_06953_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_06950_ ), .ZN(_08286_ ) );
NAND4_X1 _29141_ ( .A1(_07248_ ), .A2(_06773_ ), .A3(_06876_ ), .A4(_08286_ ), .ZN(_08287_ ) );
OAI22_X1 _29142_ ( .A1(_08238_ ), .A2(_08240_ ), .B1(_08285_ ), .B2(_08287_ ), .ZN(\idu.io_out_bits_rs2_data [25] ) );
AND3_X1 _29143_ ( .A1(_03722_ ), .A2(_03723_ ), .A3(_06766_ ), .ZN(_08288_ ) );
NOR3_X1 _29144_ ( .A1(_07195_ ), .A2(_00885_ ), .A3(_07196_ ), .ZN(_08289_ ) );
OAI22_X1 _29145_ ( .A1(\lsu.io_out_bits_rd_wdata [24] ), .A2(_07193_ ), .B1(_07194_ ), .B2(_08289_ ), .ZN(_08290_ ) );
AND3_X1 _29146_ ( .A1(_06631_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06750_ ), .ZN(_08291_ ) );
NAND3_X1 _29147_ ( .A1(_06679_ ), .A2(_06371_ ), .A3(_03832_ ), .ZN(_08292_ ) );
OAI21_X1 _29148_ ( .A(_08292_ ), .B1(_10688_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08293_ ) );
AND4_X1 _29149_ ( .A1(_06374_ ), .A2(_06587_ ), .A3(_06833_ ), .A4(_03832_ ), .ZN(_08294_ ) );
NOR3_X1 _29150_ ( .A1(_06794_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06638_ ), .ZN(_08295_ ) );
NOR3_X1 _29151_ ( .A1(_08293_ ), .A2(_08294_ ), .A3(_08295_ ), .ZN(_08296_ ) );
NAND4_X1 _29152_ ( .A1(_06663_ ), .A2(_07210_ ), .A3(_06377_ ), .A4(_06609_ ), .ZN(_08297_ ) );
OR2_X1 _29153_ ( .A1(_06799_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08298_ ) );
NAND3_X1 _29154_ ( .A1(_08296_ ), .A2(_08297_ ), .A3(_08298_ ), .ZN(_08299_ ) );
NOR3_X1 _29155_ ( .A1(_06637_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06593_ ), .ZN(_08300_ ) );
AND4_X1 _29156_ ( .A1(_06383_ ), .A2(_06723_ ), .A3(_06683_ ), .A4(_06674_ ), .ZN(_08301_ ) );
NOR3_X1 _29157_ ( .A1(_08299_ ), .A2(_08300_ ), .A3(_08301_ ), .ZN(_08302_ ) );
NAND4_X1 _29158_ ( .A1(_06664_ ), .A2(_06724_ ), .A3(_06385_ ), .A4(_03834_ ), .ZN(_08303_ ) );
NAND4_X1 _29159_ ( .A1(_06669_ ), .A2(_06724_ ), .A3(_06388_ ), .A4(_06787_ ), .ZN(_08304_ ) );
NAND3_X1 _29160_ ( .A1(_08302_ ), .A2(_08303_ ), .A3(_08304_ ), .ZN(_08305_ ) );
NOR2_X1 _29161_ ( .A1(_06809_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08306_ ) );
AND4_X1 _29162_ ( .A1(_06392_ ), .A2(_06589_ ), .A3(_06683_ ), .A4(_06787_ ), .ZN(_08307_ ) );
NOR3_X1 _29163_ ( .A1(_08305_ ), .A2(_08306_ ), .A3(_08307_ ), .ZN(_08308_ ) );
NAND4_X1 _29164_ ( .A1(_06665_ ), .A2(_06666_ ), .A3(_06394_ ), .A4(_03835_ ), .ZN(_08309_ ) );
OR3_X1 _29165_ ( .A1(_07110_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06594_ ), .ZN(_08310_ ) );
NAND3_X1 _29166_ ( .A1(_08308_ ), .A2(_08309_ ), .A3(_08310_ ), .ZN(_08311_ ) );
NOR2_X1 _29167_ ( .A1(_06677_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08312_ ) );
AND4_X1 _29168_ ( .A1(_06400_ ), .A2(_06833_ ), .A3(_06699_ ), .A4(_06690_ ), .ZN(_08313_ ) );
NOR3_X1 _29169_ ( .A1(_08311_ ), .A2(_08312_ ), .A3(_08313_ ), .ZN(_08314_ ) );
NAND4_X1 _29170_ ( .A1(_06907_ ), .A2(_06835_ ), .A3(_06402_ ), .A4(_06605_ ), .ZN(_08315_ ) );
OR3_X1 _29171_ ( .A1(_11127_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06846_ ), .ZN(_08316_ ) );
NAND3_X1 _29172_ ( .A1(_08314_ ), .A2(_08315_ ), .A3(_08316_ ), .ZN(_08317_ ) );
NOR2_X1 _29173_ ( .A1(_06840_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08318_ ) );
AND4_X1 _29174_ ( .A1(_06408_ ), .A2(_06698_ ), .A3(_06699_ ), .A4(_06691_ ), .ZN(_08319_ ) );
NOR3_X1 _29175_ ( .A1(_08317_ ), .A2(_08318_ ), .A3(_08319_ ), .ZN(_08320_ ) );
AOI22_X1 _29176_ ( .A1(_06704_ ), .A2(_06410_ ), .B1(_06606_ ), .B2(_06631_ ), .ZN(_08321_ ) );
AOI21_X1 _29177_ ( .A(_08291_ ), .B1(_08320_ ), .B2(_08321_ ), .ZN(_08322_ ) );
NOR3_X1 _29178_ ( .A1(_06802_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03837_ ), .ZN(_08323_ ) );
AND4_X1 _29179_ ( .A1(_06415_ ), .A2(_06726_ ), .A3(_07066_ ), .A4(_06606_ ), .ZN(_08324_ ) );
NOR3_X1 _29180_ ( .A1(_08322_ ), .A2(_08323_ ), .A3(_08324_ ), .ZN(_08325_ ) );
NAND4_X1 _29181_ ( .A1(_06722_ ), .A2(_06727_ ), .A3(_06417_ ), .A4(_01101_ ), .ZN(_08326_ ) );
NAND4_X1 _29182_ ( .A1(_06755_ ), .A2(_06727_ ), .A3(_06420_ ), .A4(_01101_ ), .ZN(_08327_ ) );
NAND3_X1 _29183_ ( .A1(_08325_ ), .A2(_08326_ ), .A3(_08327_ ), .ZN(_08328_ ) );
NOR2_X1 _29184_ ( .A1(_06738_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08329_ ) );
NOR3_X1 _29185_ ( .A1(_08328_ ), .A2(_06742_ ), .A3(_08329_ ), .ZN(_08330_ ) );
AOI21_X1 _29186_ ( .A(_08330_ ), .B1(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_06742_ ), .ZN(_08331_ ) );
NOR2_X1 _29187_ ( .A1(_06870_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08332_ ) );
OAI21_X1 _29188_ ( .A(_06599_ ), .B1(_06748_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08333_ ) );
NOR3_X1 _29189_ ( .A1(_08331_ ), .A2(_08332_ ), .A3(_08333_ ), .ZN(_08334_ ) );
NAND3_X1 _29190_ ( .A1(_06953_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_06950_ ), .ZN(_08335_ ) );
NAND4_X1 _29191_ ( .A1(_06771_ ), .A2(_06773_ ), .A3(_06876_ ), .A4(_08335_ ), .ZN(_08336_ ) );
OAI22_X1 _29192_ ( .A1(_08288_ ), .A2(_08290_ ), .B1(_08334_ ), .B2(_08336_ ), .ZN(\idu.io_out_bits_rs2_data [24] ) );
NAND2_X1 _29193_ ( .A1(\exu.io_out_bits_rd_wdata [23] ), .A2(_06767_ ), .ZN(_08337_ ) );
AND4_X1 _29194_ ( .A1(\wbu.io_in_bits_rd_wdata [23] ), .A2(_06782_ ), .A3(_06772_ ), .A4(_06779_ ), .ZN(_08338_ ) );
AOI21_X1 _29195_ ( .A(_08338_ ), .B1(\lsu.io_out_bits_rd_wdata [23] ), .B2(_06783_ ), .ZN(_08339_ ) );
NAND3_X1 _29196_ ( .A1(_06740_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06883_ ), .ZN(_08340_ ) );
NAND3_X1 _29197_ ( .A1(_06604_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06885_ ), .ZN(_08341_ ) );
AND3_X1 _29198_ ( .A1(_06730_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03834_ ), .ZN(_08342_ ) );
NAND3_X1 _29199_ ( .A1(_06703_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07258_ ), .ZN(_08343_ ) );
NAND3_X1 _29200_ ( .A1(_06966_ ), .A2(_06442_ ), .A3(_06673_ ), .ZN(_08344_ ) );
OAI21_X1 _29201_ ( .A(_08344_ ), .B1(_06791_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_08345_ ) );
MUX2_X1 _29202_ ( .A(_06445_ ), .B(_08345_ ), .S(_07094_ ), .Z(_08346_ ) );
OAI21_X1 _29203_ ( .A(_06972_ ), .B1(_07264_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08347_ ) );
OAI21_X1 _29204_ ( .A(_08343_ ), .B1(_08346_ ), .B2(_08347_ ), .ZN(_08348_ ) );
NAND4_X1 _29205_ ( .A1(_07215_ ), .A2(_06697_ ), .A3(_06450_ ), .A4(_06610_ ), .ZN(_08349_ ) );
OR3_X1 _29206_ ( .A1(_06637_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06593_ ), .ZN(_08350_ ) );
NAND3_X1 _29207_ ( .A1(_08348_ ), .A2(_08349_ ), .A3(_08350_ ), .ZN(_08351_ ) );
NOR3_X1 _29208_ ( .A1(_06804_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_11124_ ), .ZN(_08352_ ) );
NOR2_X1 _29209_ ( .A1(_08351_ ), .A2(_08352_ ), .ZN(_08353_ ) );
NOR2_X1 _29210_ ( .A1(_06647_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08354_ ) );
NOR2_X1 _29211_ ( .A1(_08354_ ), .A2(_06654_ ), .ZN(_08355_ ) );
AOI21_X1 _29212_ ( .A(_08342_ ), .B1(_08353_ ), .B2(_08355_ ), .ZN(_08356_ ) );
NOR2_X1 _29213_ ( .A1(_06809_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08357_ ) );
AND3_X1 _29214_ ( .A1(_06658_ ), .A2(_06460_ ), .A3(_06611_ ), .ZN(_08358_ ) );
NOR3_X1 _29215_ ( .A1(_08356_ ), .A2(_08357_ ), .A3(_08358_ ), .ZN(_08359_ ) );
NAND4_X1 _29216_ ( .A1(_06907_ ), .A2(_06910_ ), .A3(_06462_ ), .A4(_06612_ ), .ZN(_08360_ ) );
OR3_X1 _29217_ ( .A1(_07188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06690_ ), .ZN(_08361_ ) );
NAND3_X1 _29218_ ( .A1(_08359_ ), .A2(_08360_ ), .A3(_08361_ ), .ZN(_08362_ ) );
AND4_X1 _29219_ ( .A1(_06466_ ), .A2(_07057_ ), .A3(_06910_ ), .A4(_06846_ ), .ZN(_08363_ ) );
NOR2_X1 _29220_ ( .A1(_06824_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08364_ ) );
NOR3_X1 _29221_ ( .A1(_08362_ ), .A2(_08363_ ), .A3(_08364_ ), .ZN(_08365_ ) );
OR3_X1 _29222_ ( .A1(_06830_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06919_ ), .ZN(_08366_ ) );
OR3_X1 _29223_ ( .A1(_06918_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06919_ ), .ZN(_08367_ ) );
NAND3_X1 _29224_ ( .A1(_08365_ ), .A2(_08366_ ), .A3(_08367_ ), .ZN(_08368_ ) );
NOR2_X1 _29225_ ( .A1(_06841_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08369_ ) );
NOR3_X1 _29226_ ( .A1(_06844_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03837_ ), .ZN(_08370_ ) );
NOR3_X1 _29227_ ( .A1(_08368_ ), .A2(_08369_ ), .A3(_08370_ ), .ZN(_08371_ ) );
NAND4_X1 _29228_ ( .A1(_06722_ ), .A2(_06926_ ), .A3(_06474_ ), .A4(_07001_ ), .ZN(_08372_ ) );
OR2_X1 _29229_ ( .A1(_06930_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08373_ ) );
NAND3_X1 _29230_ ( .A1(_08371_ ), .A2(_08372_ ), .A3(_08373_ ), .ZN(_08374_ ) );
OAI21_X1 _29231_ ( .A(_06933_ ), .B1(_06717_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08375_ ) );
OAI21_X1 _29232_ ( .A(_08341_ ), .B1(_08374_ ), .B2(_08375_ ), .ZN(_08376_ ) );
NAND4_X1 _29233_ ( .A1(_06936_ ), .A2(_07010_ ), .A3(_06481_ ), .A4(_06938_ ), .ZN(_08377_ ) );
OR2_X1 _29234_ ( .A1(_06940_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08378_ ) );
NAND3_X1 _29235_ ( .A1(_08376_ ), .A2(_08377_ ), .A3(_08378_ ), .ZN(_08379_ ) );
OAI21_X1 _29236_ ( .A(_06943_ ), .B1(_06944_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08380_ ) );
OAI21_X1 _29237_ ( .A(_08340_ ), .B1(_08379_ ), .B2(_08380_ ), .ZN(_08381_ ) );
NAND4_X1 _29238_ ( .A1(_06948_ ), .A2(_06949_ ), .A3(_06488_ ), .A4(_06952_ ), .ZN(_08382_ ) );
AOI22_X1 _29239_ ( .A1(_06747_ ), .A2(_06491_ ), .B1(_07018_ ), .B2(_06591_ ), .ZN(_08383_ ) );
AND3_X1 _29240_ ( .A1(_08381_ ), .A2(_08382_ ), .A3(_08383_ ), .ZN(_08384_ ) );
NAND3_X1 _29241_ ( .A1(_07251_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_07080_ ), .ZN(_08385_ ) );
NAND4_X1 _29242_ ( .A1(_07248_ ), .A2(_07249_ ), .A3(_07250_ ), .A4(_08385_ ), .ZN(_08386_ ) );
OAI211_X1 _29243_ ( .A(_08337_ ), .B(_08339_ ), .C1(_08384_ ), .C2(_08386_ ), .ZN(\idu.io_out_bits_rs2_data [23] ) );
NAND2_X1 _29244_ ( .A1(\exu.io_out_bits_rd_wdata [22] ), .A2(_06767_ ), .ZN(_08387_ ) );
NOR3_X1 _29245_ ( .A1(_07195_ ), .A2(_00965_ ), .A3(_07196_ ), .ZN(_08388_ ) );
AOI22_X1 _29246_ ( .A1(\lsu.io_out_bits_rd_wdata [22] ), .A2(_06783_ ), .B1(_06875_ ), .B2(_08388_ ), .ZN(_08389_ ) );
AND4_X1 _29247_ ( .A1(_06553_ ), .A2(_06757_ ), .A3(_07067_ ), .A4(_06866_ ), .ZN(_08390_ ) );
OR2_X1 _29248_ ( .A1(_06930_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08391_ ) );
NAND3_X1 _29249_ ( .A1(_06679_ ), .A2(_06505_ ), .A3(_06814_ ), .ZN(_08392_ ) );
OAI21_X1 _29250_ ( .A(_08392_ ), .B1(_10688_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08393_ ) );
AND4_X1 _29251_ ( .A1(_06508_ ), .A2(_06587_ ), .A3(_06833_ ), .A4(_06796_ ), .ZN(_08394_ ) );
NOR3_X1 _29252_ ( .A1(_06794_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06638_ ), .ZN(_08395_ ) );
NOR3_X1 _29253_ ( .A1(_08393_ ), .A2(_08394_ ), .A3(_08395_ ), .ZN(_08396_ ) );
NAND4_X1 _29254_ ( .A1(_06663_ ), .A2(_06697_ ), .A3(_06511_ ), .A4(_06815_ ), .ZN(_08397_ ) );
OR2_X1 _29255_ ( .A1(_06799_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08398_ ) );
NAND3_X1 _29256_ ( .A1(_08396_ ), .A2(_08397_ ), .A3(_08398_ ), .ZN(_08399_ ) );
AND4_X1 _29257_ ( .A1(_06515_ ), .A2(_06897_ ), .A3(_07210_ ), .A4(_07258_ ), .ZN(_08400_ ) );
NOR3_X1 _29258_ ( .A1(_06804_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06593_ ), .ZN(_08401_ ) );
NOR3_X1 _29259_ ( .A1(_08399_ ), .A2(_08400_ ), .A3(_08401_ ), .ZN(_08402_ ) );
NAND4_X1 _29260_ ( .A1(_06665_ ), .A2(_06725_ ), .A3(_06519_ ), .A4(_06845_ ), .ZN(_08403_ ) );
NAND4_X1 _29261_ ( .A1(_06669_ ), .A2(_06725_ ), .A3(_06522_ ), .A4(_06845_ ), .ZN(_08404_ ) );
NAND3_X1 _29262_ ( .A1(_08402_ ), .A2(_08403_ ), .A3(_08404_ ), .ZN(_08405_ ) );
NOR2_X1 _29263_ ( .A1(_06809_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08406_ ) );
NOR2_X1 _29264_ ( .A1(_06661_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08407_ ) );
NOR3_X1 _29265_ ( .A1(_08405_ ), .A2(_08406_ ), .A3(_08407_ ), .ZN(_08408_ ) );
NAND4_X1 _29266_ ( .A1(_06720_ ), .A2(_06910_ ), .A3(_06527_ ), .A4(_06612_ ), .ZN(_08409_ ) );
NAND4_X1 _29267_ ( .A1(_06670_ ), .A2(_06910_ ), .A3(_06530_ ), .A4(_06612_ ), .ZN(_08410_ ) );
NAND3_X1 _29268_ ( .A1(_08408_ ), .A2(_08409_ ), .A3(_08410_ ), .ZN(_08411_ ) );
NOR2_X1 _29269_ ( .A1(_06677_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08412_ ) );
NOR2_X1 _29270_ ( .A1(_06824_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08413_ ) );
NOR3_X1 _29271_ ( .A1(_08411_ ), .A2(_08412_ ), .A3(_08413_ ), .ZN(_08414_ ) );
OR3_X1 _29272_ ( .A1(_06830_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07199_ ), .ZN(_08415_ ) );
OR3_X1 _29273_ ( .A1(_06918_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07199_ ), .ZN(_08416_ ) );
NAND3_X1 _29274_ ( .A1(_08414_ ), .A2(_08415_ ), .A3(_08416_ ), .ZN(_08417_ ) );
NOR2_X1 _29275_ ( .A1(_06841_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08418_ ) );
OAI21_X1 _29276_ ( .A(_06706_ ), .B1(_06923_ ), .B2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08419_ ) );
NOR3_X1 _29277_ ( .A1(_08417_ ), .A2(_08418_ ), .A3(_08419_ ), .ZN(_08420_ ) );
AND3_X1 _29278_ ( .A1(_06703_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06852_ ), .ZN(_08421_ ) );
OAI21_X1 _29279_ ( .A(_08391_ ), .B1(_08420_ ), .B2(_08421_ ), .ZN(_08422_ ) );
AND3_X1 _29280_ ( .A1(_06635_ ), .A2(_06543_ ), .A3(_06607_ ), .ZN(_08423_ ) );
NOR3_X1 _29281_ ( .A1(_07006_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_07007_ ), .ZN(_08424_ ) );
NOR3_X1 _29282_ ( .A1(_08422_ ), .A2(_08423_ ), .A3(_08424_ ), .ZN(_08425_ ) );
NAND4_X1 _29283_ ( .A1(_06936_ ), .A2(_06937_ ), .A3(_06547_ ), .A4(_06938_ ), .ZN(_08426_ ) );
AOI22_X1 _29284_ ( .A1(_06731_ ), .A2(_06549_ ), .B1(_06866_ ), .B2(_06735_ ), .ZN(_08427_ ) );
NAND3_X1 _29285_ ( .A1(_08425_ ), .A2(_08426_ ), .A3(_08427_ ), .ZN(_08428_ ) );
NAND3_X1 _29286_ ( .A1(_06735_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06883_ ), .ZN(_08429_ ) );
AOI21_X1 _29287_ ( .A(_08390_ ), .B1(_08428_ ), .B2(_08429_ ), .ZN(_08430_ ) );
OR2_X1 _29288_ ( .A1(_06752_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_08431_ ) );
NOR3_X1 _29289_ ( .A1(_07188_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03838_ ), .ZN(_08432_ ) );
NOR2_X1 _29290_ ( .A1(_08432_ ), .A2(_06598_ ), .ZN(_08433_ ) );
AND3_X1 _29291_ ( .A1(_08430_ ), .A2(_08431_ ), .A3(_08433_ ), .ZN(_08434_ ) );
NAND3_X1 _29292_ ( .A1(_07251_ ), .A2(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_06950_ ), .ZN(_08435_ ) );
NAND4_X1 _29293_ ( .A1(_07248_ ), .A2(_07249_ ), .A3(_07250_ ), .A4(_08435_ ), .ZN(_08436_ ) );
OAI211_X1 _29294_ ( .A(_08387_ ), .B(_08389_ ), .C1(_08434_ ), .C2(_08436_ ), .ZN(\idu.io_out_bits_rs2_data [22] ) );
OR2_X1 _29295_ ( .A1(\idu.io_out_bits_ori ), .A2(\idu.io_out_bits_addi ), .ZN(_08437_ ) );
AOI211_X1 _29296_ ( .A(\idu.io_out_bits_andi ), .B(_08437_ ), .C1(_11041_ ), .C2(_10998_ ), .ZN(_08438_ ) );
AND4_X1 _29297_ ( .A1(_10696_ ), .A2(_08438_ ), .A3(_11000_ ), .A4(_11037_ ), .ZN(_08439_ ) );
OR2_X1 _29298_ ( .A1(_03848_ ), .A2(_03846_ ), .ZN(_08440_ ) );
NAND2_X1 _29299_ ( .A1(_08440_ ), .A2(_03847_ ), .ZN(_08441_ ) );
NOR3_X1 _29300_ ( .A1(_08441_ ), .A2(\idu.io_out_bits_slli ), .A3(\idu.io_out_bits_sra ), .ZN(_08442_ ) );
INV_X1 _29301_ ( .A(\idu.io_out_bits_srai ), .ZN(_08443_ ) );
AND4_X1 _29302_ ( .A1(_10664_ ), .A2(_11013_ ), .A3(_11058_ ), .A4(_08443_ ), .ZN(_08444_ ) );
INV_X1 _29303_ ( .A(\idu.io_out_bits_xor ), .ZN(_08445_ ) );
OAI211_X1 _29304_ ( .A(_03843_ ), .B(_03842_ ), .C1(_10996_ ), .C2(_10999_ ), .ZN(_08446_ ) );
OAI211_X1 _29305_ ( .A(_03843_ ), .B(_03842_ ), .C1(_10695_ ), .C2(_10680_ ), .ZN(_08447_ ) );
OAI211_X1 _29306_ ( .A(_03843_ ), .B(_03842_ ), .C1(_10670_ ), .C2(_10681_ ), .ZN(_08448_ ) );
AND4_X1 _29307_ ( .A1(_08445_ ), .A2(_08446_ ), .A3(_08447_ ), .A4(_08448_ ), .ZN(_08449_ ) );
NAND4_X1 _29308_ ( .A1(_08439_ ), .A2(_08442_ ), .A3(_08444_ ), .A4(_08449_ ), .ZN(\idu.io_out_bits_wen_rd ) );
INV_X1 _29309_ ( .A(_11898_ ), .ZN(\ifu.io_out_bits_pc [1] ) );
INV_X1 _29310_ ( .A(_12549_ ), .ZN(\ifu.io_out_bits_pc [0] ) );
AOI21_X1 _29311_ ( .A(fanout_net_27 ), .B1(_12656_ ), .B2(_12658_ ), .ZN(_08450_ ) );
INV_X1 _29312_ ( .A(_08450_ ), .ZN(\ifu.ren_REG_$_DFF_P__Q_D ) );
NAND3_X1 _29313_ ( .A1(_10712_ ), .A2(_10987_ ), .A3(\ifu.state [1] ), .ZN(_08451_ ) );
NAND4_X1 _29314_ ( .A1(_12200_ ), .A2(\ifu.state [0] ), .A3(_12201_ ), .A4(_12048_ ), .ZN(_08452_ ) );
NAND2_X1 _29315_ ( .A1(_08451_ ), .A2(_08452_ ), .ZN(\ifu.state_$_DFF_P__Q_1_D ) );
AOI22_X1 _29316_ ( .A1(_10829_ ), .A2(_10830_ ), .B1(_10700_ ), .B2(_10702_ ), .ZN(_08453_ ) );
AND2_X1 _29317_ ( .A1(_10711_ ), .A2(_08453_ ), .ZN(_08454_ ) );
INV_X1 _29318_ ( .A(_08454_ ), .ZN(_08455_ ) );
NAND2_X1 _29319_ ( .A1(_10710_ ), .A2(_12048_ ), .ZN(_08456_ ) );
NAND4_X1 _29320_ ( .A1(_08455_ ), .A2(_10922_ ), .A3(\ifu.state [0] ), .A4(_08456_ ), .ZN(_08457_ ) );
NAND3_X1 _29321_ ( .A1(_idu_io_in_bits_T ), .A2(_10922_ ), .A3(\ifu.state [1] ), .ZN(_08458_ ) );
NAND4_X1 _29322_ ( .A1(_10829_ ), .A2(_10922_ ), .A3(_10830_ ), .A4(\ifu.state [2] ), .ZN(_08459_ ) );
NAND4_X1 _29323_ ( .A1(_08457_ ), .A2(_08458_ ), .A3(\ifu.ren_REG_$_DFF_P__Q_D_$_NAND__Y_B ), .A4(_08459_ ), .ZN(\ifu.state_$_DFF_P__Q_2_D ) );
NAND3_X1 _29324_ ( .A1(_08450_ ), .A2(\ifu.state [1] ), .A3(_12657_ ), .ZN(_08460_ ) );
NAND3_X1 _29325_ ( .A1(_10832_ ), .A2(_11892_ ), .A3(\ifu.state [2] ), .ZN(_08461_ ) );
NAND3_X1 _29326_ ( .A1(_10711_ ), .A2(\ifu.state [0] ), .A3(_08453_ ), .ZN(_08462_ ) );
NAND3_X1 _29327_ ( .A1(_08460_ ), .A2(_08461_ ), .A3(_08462_ ), .ZN(\ifu.state_$_DFF_P__Q_D ) );
OR3_X1 _29328_ ( .A1(_01067_ ), .A2(io_master_wready_$_ANDNOT__B_Y_$_OR__A_B ), .A3(_10708_ ), .ZN(_08463_ ) );
OR3_X1 _29329_ ( .A1(_08463_ ), .A2(\lsu.state [1] ), .A3(_10823_ ), .ZN(_08464_ ) );
BUF_X4 _29330_ ( .A(_08464_ ), .Z(_08465_ ) );
BUF_X4 _29331_ ( .A(_08465_ ), .Z(_08466_ ) );
AOI21_X1 _29332_ ( .A(_09772_ ), .B1(_08466_ ), .B2(_01065_ ), .ZN(_08467_ ) );
AOI21_X1 _29333_ ( .A(_00973_ ), .B1(_04982_ ), .B2(_04983_ ), .ZN(_08468_ ) );
NOR2_X2 _29334_ ( .A1(_08468_ ), .A2(\arbiter._io_axi_araddr_T ), .ZN(_08469_ ) );
BUF_X4 _29335_ ( .A(_08469_ ), .Z(_08470_ ) );
MUX2_X1 _29336_ ( .A(\io_master_awaddr [31] ), .B(_08467_ ), .S(_08470_ ), .Z(\io_master_araddr [31] ) );
AOI21_X1 _29337_ ( .A(_09717_ ), .B1(_08466_ ), .B2(_01065_ ), .ZN(_08471_ ) );
MUX2_X1 _29338_ ( .A(\io_master_awaddr [30] ), .B(_08471_ ), .S(_08470_ ), .Z(\io_master_araddr [30] ) );
AND2_X1 _29339_ ( .A1(_08465_ ), .A2(_01063_ ), .ZN(_08472_ ) );
INV_X1 _29340_ ( .A(_08469_ ), .ZN(_08473_ ) );
NOR2_X1 _29341_ ( .A1(_08472_ ), .A2(_08473_ ), .ZN(_08474_ ) );
INV_X2 _29342_ ( .A(_08474_ ), .ZN(_08475_ ) );
BUF_X4 _29343_ ( .A(_08475_ ), .Z(_08476_ ) );
INV_X1 _29344_ ( .A(_09611_ ), .ZN(_08477_ ) );
BUF_X4 _29345_ ( .A(_08469_ ), .Z(_08478_ ) );
OAI22_X1 _29346_ ( .A1(_08476_ ), .A2(_08477_ ), .B1(_08549_ ), .B2(_08478_ ), .ZN(\io_master_araddr [21] ) );
OAI22_X1 _29347_ ( .A1(_08476_ ), .A2(_10057_ ), .B1(_08550_ ), .B2(_08478_ ), .ZN(\io_master_araddr [20] ) );
BUF_X4 _29348_ ( .A(_08469_ ), .Z(_08479_ ) );
OAI22_X1 _29349_ ( .A1(_08476_ ), .A2(_09969_ ), .B1(_08553_ ), .B2(_08479_ ), .ZN(\io_master_araddr [19] ) );
OAI22_X1 _29350_ ( .A1(_08476_ ), .A2(_10013_ ), .B1(_08554_ ), .B2(_08479_ ), .ZN(\io_master_araddr [18] ) );
AOI21_X1 _29351_ ( .A(_10104_ ), .B1(_08466_ ), .B2(_01065_ ), .ZN(_08480_ ) );
BUF_X4 _29352_ ( .A(_08469_ ), .Z(_08481_ ) );
MUX2_X1 _29353_ ( .A(\io_master_awaddr [17] ), .B(_08480_ ), .S(_08481_ ), .Z(\io_master_araddr [17] ) );
AOI21_X1 _29354_ ( .A(_09918_ ), .B1(_08466_ ), .B2(_01064_ ), .ZN(_08482_ ) );
MUX2_X1 _29355_ ( .A(\io_master_awaddr [16] ), .B(_08482_ ), .S(_08481_ ), .Z(\io_master_araddr [16] ) );
AOI21_X1 _29356_ ( .A(_09869_ ), .B1(_08465_ ), .B2(_01064_ ), .ZN(_08483_ ) );
MUX2_X1 _29357_ ( .A(\io_master_awaddr [15] ), .B(_08483_ ), .S(_08481_ ), .Z(\io_master_araddr [15] ) );
AOI21_X1 _29358_ ( .A(_10153_ ), .B1(_08465_ ), .B2(_01064_ ), .ZN(_08484_ ) );
MUX2_X1 _29359_ ( .A(\io_master_awaddr [14] ), .B(_08484_ ), .S(_08481_ ), .Z(\io_master_araddr [14] ) );
OAI22_X1 _29360_ ( .A1(_08476_ ), .A2(_10202_ ), .B1(_03866_ ), .B2(_08479_ ), .ZN(\io_master_araddr [13] ) );
AOI21_X1 _29361_ ( .A(_11483_ ), .B1(_08465_ ), .B2(_01064_ ), .ZN(_08485_ ) );
MUX2_X1 _29362_ ( .A(\io_master_awaddr [12] ), .B(_08485_ ), .S(_08481_ ), .Z(\io_master_araddr [12] ) );
OAI22_X1 _29363_ ( .A1(_08476_ ), .A2(_11312_ ), .B1(_08541_ ), .B2(_08479_ ), .ZN(\io_master_araddr [29] ) );
AOI21_X1 _29364_ ( .A(_10349_ ), .B1(_08465_ ), .B2(_01064_ ), .ZN(_08486_ ) );
MUX2_X1 _29365_ ( .A(\io_master_awaddr [11] ), .B(_08486_ ), .S(_08481_ ), .Z(\io_master_araddr [11] ) );
OAI22_X1 _29366_ ( .A1(_08476_ ), .A2(_11484_ ), .B1(_03867_ ), .B2(_08479_ ), .ZN(\io_master_araddr [10] ) );
OAI22_X1 _29367_ ( .A1(_08476_ ), .A2(_11482_ ), .B1(_04745_ ), .B2(_08479_ ), .ZN(\io_master_araddr [9] ) );
AOI21_X1 _29368_ ( .A(_11326_ ), .B1(_08465_ ), .B2(_01064_ ), .ZN(_08487_ ) );
MUX2_X1 _29369_ ( .A(\io_master_awaddr [8] ), .B(_08487_ ), .S(_08481_ ), .Z(\io_master_araddr [8] ) );
OAI22_X1 _29370_ ( .A1(_08475_ ), .A2(_11327_ ), .B1(_04740_ ), .B2(_08479_ ), .ZN(\io_master_araddr [7] ) );
OAI22_X1 _29371_ ( .A1(_08475_ ), .A2(_11954_ ), .B1(_04747_ ), .B2(_08479_ ), .ZN(\io_master_araddr [6] ) );
OAI22_X1 _29372_ ( .A1(_08475_ ), .A2(_11956_ ), .B1(_08536_ ), .B2(_08479_ ), .ZN(\io_master_araddr [5] ) );
OAI22_X1 _29373_ ( .A1(_08475_ ), .A2(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__A_Y ), .B1(_08537_ ), .B2(_08479_ ), .ZN(\io_master_araddr [4] ) );
NAND3_X1 _29374_ ( .A1(_11581_ ), .A2(_11997_ ), .A3(_11583_ ), .ZN(_08488_ ) );
AOI21_X1 _29375_ ( .A(_08488_ ), .B1(_08466_ ), .B2(_01065_ ), .ZN(_08489_ ) );
NAND2_X1 _29376_ ( .A1(_08489_ ), .A2(_08470_ ), .ZN(_08490_ ) );
OAI21_X1 _29377_ ( .A(_08490_ ), .B1(_08538_ ), .B2(_08478_ ), .ZN(\io_master_araddr [3] ) );
NAND3_X1 _29378_ ( .A1(_11581_ ), .A2(_11994_ ), .A3(_11583_ ), .ZN(_08491_ ) );
AOI21_X1 _29379_ ( .A(_08491_ ), .B1(_08466_ ), .B2(_01065_ ), .ZN(_08492_ ) );
NAND2_X1 _29380_ ( .A1(_08492_ ), .A2(_08470_ ), .ZN(_08493_ ) );
OAI21_X1 _29381_ ( .A(_08493_ ), .B1(_00981_ ), .B2(_08478_ ), .ZN(\io_master_araddr [2] ) );
OAI22_X1 _29382_ ( .A1(_08475_ ), .A2(_09406_ ), .B1(_04741_ ), .B2(_08470_ ), .ZN(\io_master_araddr [28] ) );
NAND4_X1 _29383_ ( .A1(_11488_ ), .A2(_11363_ ), .A3(_11364_ ), .A4(_11492_ ), .ZN(_08494_ ) );
AOI21_X1 _29384_ ( .A(_08494_ ), .B1(_08466_ ), .B2(_01065_ ), .ZN(_08495_ ) );
NAND2_X1 _29385_ ( .A1(_08495_ ), .A2(_08470_ ), .ZN(_08496_ ) );
OAI21_X1 _29386_ ( .A(_08496_ ), .B1(_03872_ ), .B2(_08478_ ), .ZN(\io_master_araddr [1] ) );
NAND4_X1 _29387_ ( .A1(_11488_ ), .A2(_11403_ ), .A3(_11404_ ), .A4(_11492_ ), .ZN(_08497_ ) );
AOI21_X1 _29388_ ( .A(_08497_ ), .B1(_08466_ ), .B2(_01065_ ), .ZN(_08498_ ) );
NAND2_X1 _29389_ ( .A1(_08498_ ), .A2(_08470_ ), .ZN(_08499_ ) );
OAI21_X1 _29390_ ( .A(_08499_ ), .B1(_04469_ ), .B2(_08478_ ), .ZN(\io_master_araddr [0] ) );
AND3_X1 _29391_ ( .A1(_09465_ ), .A2(_09466_ ), .A3(_09467_ ), .ZN(_08500_ ) );
AOI221_X4 _29392_ ( .A(_08500_ ), .B1(\ifu.io_out_bits_pc_$_NOT__Y_A_$_MUX__Y_B ), .B2(\ifu._start_T ), .C1(_08465_ ), .C2(_01064_ ), .ZN(_08501_ ) );
MUX2_X1 _29393_ ( .A(\io_master_awaddr [27] ), .B(_08501_ ), .S(_08481_ ), .Z(\io_master_araddr [27] ) );
INV_X1 _29394_ ( .A(_09189_ ), .ZN(_08502_ ) );
OAI22_X1 _29395_ ( .A1(_08475_ ), .A2(_08502_ ), .B1(_08533_ ), .B2(_08470_ ), .ZN(\io_master_araddr [26] ) );
INV_X1 _29396_ ( .A(_11304_ ), .ZN(_08503_ ) );
OAI22_X1 _29397_ ( .A1(_08475_ ), .A2(_08503_ ), .B1(_03860_ ), .B2(_08470_ ), .ZN(\io_master_araddr [25] ) );
OAI22_X1 _29398_ ( .A1(_08475_ ), .A2(_11303_ ), .B1(_08534_ ), .B2(_08470_ ), .ZN(\io_master_araddr [24] ) );
AOI21_X1 _29399_ ( .A(_11308_ ), .B1(_08465_ ), .B2(_01064_ ), .ZN(_08504_ ) );
MUX2_X1 _29400_ ( .A(\io_master_awaddr [23] ), .B(_08504_ ), .S(_08481_ ), .Z(\io_master_araddr [23] ) );
AOI21_X1 _29401_ ( .A(_09563_ ), .B1(_08465_ ), .B2(_01064_ ), .ZN(_08505_ ) );
MUX2_X1 _29402_ ( .A(\io_master_awaddr [22] ), .B(_08505_ ), .S(_08481_ ), .Z(\io_master_araddr [22] ) );
NAND3_X1 _29403_ ( .A1(_08466_ ), .A2(_01065_ ), .A3(_08478_ ), .ZN(\io_master_arburst [0] ) );
AOI211_X1 _29404_ ( .A(_12090_ ), .B(_08473_ ), .C1(_08466_ ), .C2(_01065_ ), .ZN(\io_master_arlen [0] ) );
NOR3_X1 _29405_ ( .A1(_08478_ ), .A2(\arbiter.io_lsu_arsize [1] ), .A3(_04902_ ), .ZN(\io_master_arsize [0] ) );
OAI21_X1 _29406_ ( .A(_08476_ ), .B1(_03900_ ), .B2(_08478_ ), .ZN(\io_master_arsize [1] ) );
INV_X1 _29407_ ( .A(_01057_ ), .ZN(_08506_ ) );
OAI22_X1 _29408_ ( .A1(_08463_ ), .A2(_08506_ ), .B1(_04750_ ), .B2(_00973_ ), .ZN(io_master_arvalid ) );
OAI21_X1 _29409_ ( .A(\arbiter._clink_io_axi_araddr_T ), .B1(_10824_ ), .B2(\lsu._io_axi_awvalid_T_1 ), .ZN(_08507_ ) );
AND4_X1 _29410_ ( .A1(_08541_ ), .A2(_08540_ ), .A3(_08542_ ), .A4(_08545_ ), .ZN(_08508_ ) );
AND3_X1 _29411_ ( .A1(_08556_ ), .A2(_08557_ ), .A3(_08558_ ), .ZN(_08509_ ) );
AOI21_X1 _29412_ ( .A(_08507_ ), .B1(_08508_ ), .B2(_08509_ ), .ZN(io_master_awvalid ) );
OAI21_X1 _29413_ ( .A(_08476_ ), .B1(_03919_ ), .B2(_08478_ ), .ZN(io_master_rready ) );
OR3_X1 _29414_ ( .A1(\io_master_awaddr [0] ), .A2(\io_master_awsize [1] ), .A3(\io_master_awsize [0] ), .ZN(_08510_ ) );
OR3_X1 _29415_ ( .A1(\io_master_awsize [1] ), .A2(\lsu._GEN_1 [0] ), .A3(\io_master_awsize [0] ), .ZN(_08511_ ) );
AND3_X1 _29416_ ( .A1(_08510_ ), .A2(_08511_ ), .A3(io_master_wstrb_$_ANDNOT__Y_A ), .ZN(\io_master_wstrb [1] ) );
AND3_X1 _29417_ ( .A1(_08511_ ), .A2(_03872_ ), .A3(lsu_io_in_bits_r_sb_$_ANDNOT__B_Y_$_ANDNOT__B_A ), .ZN(\io_master_wstrb [0] ) );
OR2_X1 _29418_ ( .A1(\io_master_awaddr [1] ), .A2(\io_master_awsize [1] ), .ZN(_08512_ ) );
AND3_X1 _29419_ ( .A1(_08510_ ), .A2(_08511_ ), .A3(_08512_ ), .ZN(\io_master_wstrb [3] ) );
AOI21_X1 _29420_ ( .A(_03872_ ), .B1(_08511_ ), .B2(lsu_io_in_bits_r_sb_$_ANDNOT__B_Y_$_ANDNOT__B_A ), .ZN(_08513_ ) );
AOI211_X1 _29421_ ( .A(\io_master_awaddr [1] ), .B(\io_master_awsize [1] ), .C1(\io_master_awaddr [0] ), .C2(\io_master_awsize [0] ), .ZN(_08514_ ) );
NOR2_X1 _29422_ ( .A1(_08513_ ), .A2(_08514_ ), .ZN(\io_master_wstrb [2] ) );
AND2_X1 _29423_ ( .A1(io_slave_wvalid ), .A2(io_slave_awvalid ), .ZN(io_slave_bvalid ) );
AND2_X1 _29424_ ( .A1(io_master_awready ), .A2(io_master_wready ), .ZN(_08515_ ) );
OAI21_X1 _29425_ ( .A(\arbiter._clink_io_axi_araddr_T ), .B1(_08562_ ), .B2(_08515_ ), .ZN(_08516_ ) );
NOR2_X1 _29426_ ( .A1(_08516_ ), .A2(io_master_wready_$_ANDNOT__B_Y_$_OR__A_B ), .ZN(_08517_ ) );
NOR2_X1 _29427_ ( .A1(\lsu._io_axi_awvalid_T_1 ), .A2(\lsu._io_in_ready_T ), .ZN(_08518_ ) );
NOR4_X1 _29428_ ( .A1(_08517_ ), .A2(fanout_net_27 ), .A3(_01056_ ), .A4(_08518_ ), .ZN(\lsu.state_$_DFF_P__Q_1_D ) );
OAI21_X1 _29429_ ( .A(\arbiter._clink_io_axi_araddr_T ), .B1(_08563_ ), .B2(\arbiter.clink.io_axi_rvalid_REG_$_NOT__A_Y ), .ZN(_08519_ ) );
AOI21_X1 _29430_ ( .A(io_master_arready ), .B1(_04982_ ), .B2(_04983_ ), .ZN(_08520_ ) );
NOR2_X1 _29431_ ( .A1(_08519_ ), .A2(_08520_ ), .ZN(_08521_ ) );
INV_X1 _29432_ ( .A(_10824_ ), .ZN(_08522_ ) );
OAI211_X1 _29433_ ( .A(\lsu._io_in_ready_T ), .B(_10823_ ), .C1(_08517_ ), .C2(_08522_ ), .ZN(_08523_ ) );
INV_X1 _29434_ ( .A(\lsu.state [1] ), .ZN(_08524_ ) );
AOI211_X1 _29435_ ( .A(fanout_net_27 ), .B(_08521_ ), .C1(_08523_ ), .C2(_08524_ ), .ZN(\lsu.state_$_DFF_P__Q_2_D ) );
OAI211_X1 _29436_ ( .A(_10991_ ), .B(\ifu.ren_REG_$_DFF_P__Q_D_$_NAND__Y_B ), .C1(_03919_ ), .C2(_01070_ ), .ZN(\lsu.state_$_DFF_P__Q_3_D ) );
NOR3_X1 _29437_ ( .A1(_03919_ ), .A2(fanout_net_27 ), .A3(\arbiter.lsu_end ), .ZN(_08525_ ) );
NOR2_X1 _29438_ ( .A1(_10825_ ), .A2(fanout_net_27 ), .ZN(_08526_ ) );
OAI211_X1 _29439_ ( .A(\lsu._io_in_ready_T ), .B(_08526_ ), .C1(_08517_ ), .C2(_08522_ ), .ZN(_08527_ ) );
INV_X1 _29440_ ( .A(_08521_ ), .ZN(_08528_ ) );
AOI21_X1 _29441_ ( .A(_08527_ ), .B1(_10823_ ), .B2(_08528_ ), .ZN(_08529_ ) );
AND3_X1 _29442_ ( .A1(_08517_ ), .A2(_10845_ ), .A3(\lsu._io_axi_awvalid_T_1 ), .ZN(_08530_ ) );
NOR4_X1 _29443_ ( .A1(_08519_ ), .A2(fanout_net_27 ), .A3(_08524_ ), .A4(_08520_ ), .ZN(_08531_ ) );
OR4_X1 _29444_ ( .A1(_08525_ ), .A2(_08529_ ), .A3(_08530_ ), .A4(_08531_ ), .ZN(\lsu.state_$_DFF_P__Q_D ) );
NOR2_X1 _29445_ ( .A1(_12855_ ), .A2(\wbu.io_in_bits_csr_waddr [0] ), .ZN(wbu_io_in_bits_csr_waddr_$_ANDNOT__A_Y ) );
AND3_X1 _29446_ ( .A1(\wbu.io_in_bits_ecall ), .A2(\wbu.io_in_bits_wen_csr ), .A3(\ifu.io_valid ), .ZN(\wbu.csr_0_$_SDFFE_PP0P__Q_E ) );
AND4_X1 _29447_ ( .A1(fanout_net_36 ), .A2(_13181_ ), .A3(_13474_ ), .A4(_13183_ ), .ZN(\wbu.rf_31_$_SDFFE_PP0P__Q_E ) );
CLKGATE_X1 _29448_ ( .CK(clock ), .E(_wbu_io_in_bits_T ), .GCK(_13931_ ) );
CLKGATE_X1 _29449_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_13932_ ) );
CLKGATE_X1 _29450_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_Y ), .GCK(_13933_ ) );
CLKGATE_X1 _29451_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_Y ), .GCK(_13934_ ) );
CLKGATE_X1 _29452_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .GCK(_13935_ ) );
CLKGATE_X1 _29453_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_13936_ ) );
CLKGATE_X1 _29454_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_13937_ ) );
CLKGATE_X1 _29455_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_Y ), .GCK(_13938_ ) );
CLKGATE_X1 _29456_ ( .CK(clock ), .E(\wbu.rf_31_$_SDFFE_PP0P__Q_E ), .GCK(_13939_ ) );
CLKGATE_X1 _29457_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .GCK(_13940_ ) );
CLKGATE_X1 _29458_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .GCK(_13941_ ) );
CLKGATE_X1 _29459_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .GCK(_13942_ ) );
CLKGATE_X1 _29460_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_1_Y ), .GCK(_13943_ ) );
CLKGATE_X1 _29461_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .GCK(_13944_ ) );
CLKGATE_X1 _29462_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_Y_$_ANDNOT__B_1_Y ), .GCK(_13945_ ) );
CLKGATE_X1 _29463_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .GCK(_13946_ ) );
CLKGATE_X1 _29464_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_Y_$_ANDNOT__B_1_Y ), .GCK(_13947_ ) );
CLKGATE_X1 _29465_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .GCK(_13948_ ) );
CLKGATE_X1 _29466_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .GCK(_13949_ ) );
CLKGATE_X1 _29467_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__A_Y_$_ANDNOT__B_1_Y ), .GCK(_13950_ ) );
CLKGATE_X1 _29468_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .GCK(_13951_ ) );
CLKGATE_X1 _29469_ ( .CK(clock ), .E(_00000_ ), .GCK(_13952_ ) );
CLKGATE_X1 _29470_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_2_Y_$_ANDNOT__B_1_Y ), .GCK(_13953_ ) );
CLKGATE_X1 _29471_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_1_Y_$_ANDNOT__B_1_Y ), .GCK(_13954_ ) );
CLKGATE_X1 _29472_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_13955_ ) );
CLKGATE_X1 _29473_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_ANDNOT__B_Y ), .GCK(_13956_ ) );
CLKGATE_X1 _29474_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_1_Y ), .GCK(_13957_ ) );
CLKGATE_X1 _29475_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_13958_ ) );
CLKGATE_X1 _29476_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__A_B_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_13959_ ) );
CLKGATE_X1 _29477_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_13960_ ) );
CLKGATE_X1 _29478_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_1_Y_$_ANDNOT__B_Y ), .GCK(_13961_ ) );
CLKGATE_X1 _29479_ ( .CK(clock ), .E(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_1_A_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_13962_ ) );
CLKGATE_X1 _29480_ ( .CK(clock ), .E(wbu_io_in_bits_csr_waddr_$_AND__A_Y ), .GCK(_13963_ ) );
CLKGATE_X1 _29481_ ( .CK(clock ), .E(wbu_io_in_bits_csr_waddr_$_ANDNOT__A_Y ), .GCK(_13964_ ) );
CLKGATE_X1 _29482_ ( .CK(clock ), .E(_00001_ ), .GCK(_13965_ ) );
CLKGATE_X1 _29483_ ( .CK(clock ), .E(\wbu.csr_0_$_SDFFE_PP0P__Q_E ), .GCK(_13966_ ) );
CLKGATE_X1 _29484_ ( .CK(clock ), .E(_lsu_io_in_bits_T ), .GCK(_13967_ ) );
CLKGATE_X1 _29485_ ( .CK(clock ), .E(\ifu._start_T ), .GCK(_13968_ ) );
CLKGATE_X1 _29486_ ( .CK(clock ), .E(\ifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_13969_ ) );
CLKGATE_X1 _29487_ ( .CK(clock ), .E(_idu_io_in_bits_T ), .GCK(_13970_ ) );
CLKGATE_X1 _29488_ ( .CK(clock ), .E(\arbiter.io_ifu_araddr [4] ), .GCK(_13971_ ) );
CLKGATE_X1 _29489_ ( .CK(clock ), .E(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__A_Y ), .GCK(_13972_ ) );
CLKGATE_X1 _29490_ ( .CK(clock ), .E(\icache.valid_reg_1_$_MUX__A_Y_$_OR__B_A_$_ANDNOT__A_Y ), .GCK(_13973_ ) );
CLKGATE_X1 _29491_ ( .CK(clock ), .E(\icache.valid_reg_1_$_MUX__A_Y_$_OR__B_A_$_ANDNOT__A_1_Y ), .GCK(_13974_ ) );
CLKGATE_X1 _29492_ ( .CK(clock ), .E(\icache.offset_buf_$_SDFFE_PP0P__Q_E ), .GCK(_13975_ ) );
CLKGATE_X1 _29493_ ( .CK(clock ), .E(\icache.icache_reg_1_3_$_SDFFE_PP0P__Q_E ), .GCK(_13976_ ) );
CLKGATE_X1 _29494_ ( .CK(clock ), .E(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_NOR__A_Y ), .GCK(_13977_ ) );
CLKGATE_X1 _29495_ ( .CK(clock ), .E(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_NOR__A_Y ), .GCK(_13978_ ) );
CLKGATE_X1 _29496_ ( .CK(clock ), .E(\icache.offset_buf_$_OR__A_Y_$_NOR__A_Y ), .GCK(_13979_ ) );
CLKGATE_X1 _29497_ ( .CK(clock ), .E(\icache.offset_buf_$_NAND__A_Y_$_ANDNOT__B_Y ), .GCK(_13980_ ) );
CLKGATE_X1 _29498_ ( .CK(clock ), .E(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_A_$_ANDNOT__B_Y ), .GCK(_13981_ ) );
CLKGATE_X1 _29499_ ( .CK(clock ), .E(\icache.offset_buf_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_AND__Y_B_$_ANDNOT__B_Y ), .GCK(_13982_ ) );
CLKGATE_X1 _29500_ ( .CK(clock ), .E(\icache.offset_buf_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_13983_ ) );
CLKGATE_X1 _29501_ ( .CK(clock ), .E(_exu_io_in_bits_T ), .GCK(_13984_ ) );
LOGIC1_X1 _29502_ ( .Z(\io_master_awburst [0] ) );
LOGIC0_X1 _29503_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q ( .D(_00002_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [31] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_1 ( .D(_00003_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [30] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_1_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_10 ( .D(_00004_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [21] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_10_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_11 ( .D(_00005_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [20] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_11_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_12 ( .D(_00006_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [19] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_12_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_13 ( .D(_00007_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [18] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_13_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_14 ( .D(_00008_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [17] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_14_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_15 ( .D(_00009_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [16] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_15_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_16 ( .D(_00010_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [15] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_16_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_17 ( .D(_00011_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [14] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_17_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_18 ( .D(_00012_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [13] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_18_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_19 ( .D(_00013_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [12] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_19_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_2 ( .D(_00014_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [29] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_2_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_20 ( .D(_00015_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [11] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_20_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_21 ( .D(_00016_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [10] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_21_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_22 ( .D(_00017_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [9] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_22_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_23 ( .D(_00018_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [8] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_23_B_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_24 ( .D(_00019_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [7] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_8_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_25 ( .D(_00020_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [6] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_9_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_26 ( .D(_00021_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [5] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_10_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_27 ( .D(_00022_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [4] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_11_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_28 ( .D(_00023_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [3] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_12_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_29 ( .D(_00024_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [2] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_13_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_3 ( .D(_00025_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [28] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_3_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_30 ( .D(_00026_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [1] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_14_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_31 ( .D(_00027_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [0] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_15_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_4 ( .D(_00028_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [27] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_4_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_5 ( .D(_00029_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [26] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_5_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_6 ( .D(_00030_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [25] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_6_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_7 ( .D(_00031_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [24] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_7_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_8 ( .D(_00032_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [23] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_8_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rdata_REG_$_SDFF_PN0__Q_9 ( .D(_00033_ ), .CK(clock ), .Q(\arbiter.clink.io_axi_rdata [22] ), .QN(lsu_io_out_bits_rd_wdata_$_MUX__Y_9_B_$_OR__Y_A_$_OR__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \arbiter.clink.io_axi_rvalid_REG_$_DFF_P__Q ( .D(\arbiter.clink.io_axi_arvalid ), .CK(clock ), .Q(\arbiter.clink.io_axi_rvalid ), .QN(\arbiter.clink.io_axi_rvalid_REG_$_NOT__A_Y ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q ( .D(_00034_ ), .CK(clock ), .Q(\arbiter.clink.mtime [63] ), .QN(_14583_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_1 ( .D(_00035_ ), .CK(clock ), .Q(\arbiter.clink.mtime [62] ), .QN(_14582_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_10 ( .D(_00036_ ), .CK(clock ), .Q(\arbiter.clink.mtime [53] ), .QN(_14581_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_11 ( .D(_00037_ ), .CK(clock ), .Q(\arbiter.clink.mtime [52] ), .QN(_14580_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_12 ( .D(_00038_ ), .CK(clock ), .Q(\arbiter.clink.mtime [51] ), .QN(_14579_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_13 ( .D(_00039_ ), .CK(clock ), .Q(\arbiter.clink.mtime [50] ), .QN(_14578_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_14 ( .D(_00040_ ), .CK(clock ), .Q(\arbiter.clink.mtime [49] ), .QN(_14577_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_15 ( .D(_00041_ ), .CK(clock ), .Q(\arbiter.clink.mtime [48] ), .QN(_14576_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_16 ( .D(_00042_ ), .CK(clock ), .Q(\arbiter.clink.mtime [47] ), .QN(_14575_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_17 ( .D(_00043_ ), .CK(clock ), .Q(\arbiter.clink.mtime [46] ), .QN(_14574_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_18 ( .D(_00044_ ), .CK(clock ), .Q(\arbiter.clink.mtime [45] ), .QN(_14573_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_19 ( .D(_00045_ ), .CK(clock ), .Q(\arbiter.clink.mtime [44] ), .QN(_14572_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_2 ( .D(_00046_ ), .CK(clock ), .Q(\arbiter.clink.mtime [61] ), .QN(_14571_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_20 ( .D(_00047_ ), .CK(clock ), .Q(\arbiter.clink.mtime [43] ), .QN(_14570_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_21 ( .D(_00048_ ), .CK(clock ), .Q(\arbiter.clink.mtime [42] ), .QN(_14569_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_22 ( .D(_00049_ ), .CK(clock ), .Q(\arbiter.clink.mtime [41] ), .QN(_14568_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_23 ( .D(_00050_ ), .CK(clock ), .Q(\arbiter.clink.mtime [40] ), .QN(_14567_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_24 ( .D(_00051_ ), .CK(clock ), .Q(\arbiter.clink.mtime [39] ), .QN(_14566_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_25 ( .D(_00052_ ), .CK(clock ), .Q(\arbiter.clink.mtime [38] ), .QN(_14565_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_26 ( .D(_00053_ ), .CK(clock ), .Q(\arbiter.clink.mtime [37] ), .QN(_14564_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_27 ( .D(_00054_ ), .CK(clock ), .Q(\arbiter.clink.mtime [36] ), .QN(_14563_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_28 ( .D(_00055_ ), .CK(clock ), .Q(\arbiter.clink.mtime [35] ), .QN(_14562_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_29 ( .D(_00056_ ), .CK(clock ), .Q(\arbiter.clink.mtime [34] ), .QN(_14561_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_3 ( .D(_00057_ ), .CK(clock ), .Q(\arbiter.clink.mtime [60] ), .QN(_14560_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_30 ( .D(_00058_ ), .CK(clock ), .Q(\arbiter.clink.mtime [33] ), .QN(_14559_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_31 ( .D(_00059_ ), .CK(clock ), .Q(\arbiter.clink.mtime [32] ), .QN(_14558_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_32 ( .D(_00060_ ), .CK(clock ), .Q(\arbiter.clink.mtime [31] ), .QN(_14557_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_33 ( .D(_00061_ ), .CK(clock ), .Q(\arbiter.clink.mtime [30] ), .QN(_14556_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_34 ( .D(_00062_ ), .CK(clock ), .Q(\arbiter.clink.mtime [29] ), .QN(_14555_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_35 ( .D(_00063_ ), .CK(clock ), .Q(\arbiter.clink.mtime [28] ), .QN(_14554_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_36 ( .D(_00064_ ), .CK(clock ), .Q(\arbiter.clink.mtime [27] ), .QN(_14553_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_37 ( .D(_00065_ ), .CK(clock ), .Q(\arbiter.clink.mtime [26] ), .QN(_14552_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_38 ( .D(_00066_ ), .CK(clock ), .Q(\arbiter.clink.mtime [25] ), .QN(_14551_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_39 ( .D(_00067_ ), .CK(clock ), .Q(\arbiter.clink.mtime [24] ), .QN(_14550_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_4 ( .D(_00068_ ), .CK(clock ), .Q(\arbiter.clink.mtime [59] ), .QN(_14549_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_40 ( .D(_00069_ ), .CK(clock ), .Q(\arbiter.clink.mtime [23] ), .QN(_14548_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_41 ( .D(_00070_ ), .CK(clock ), .Q(\arbiter.clink.mtime [22] ), .QN(_14547_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_42 ( .D(_00071_ ), .CK(clock ), .Q(\arbiter.clink.mtime [21] ), .QN(_14546_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_43 ( .D(_00072_ ), .CK(clock ), .Q(\arbiter.clink.mtime [20] ), .QN(_14545_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_44 ( .D(_00073_ ), .CK(clock ), .Q(\arbiter.clink.mtime [19] ), .QN(_14544_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_45 ( .D(_00074_ ), .CK(clock ), .Q(\arbiter.clink.mtime [18] ), .QN(_14543_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_46 ( .D(_00075_ ), .CK(clock ), .Q(\arbiter.clink.mtime [17] ), .QN(_14542_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_47 ( .D(_00076_ ), .CK(clock ), .Q(\arbiter.clink.mtime [16] ), .QN(_14541_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_48 ( .D(_00077_ ), .CK(clock ), .Q(\arbiter.clink.mtime [15] ), .QN(_14540_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_49 ( .D(_00078_ ), .CK(clock ), .Q(\arbiter.clink.mtime [14] ), .QN(_14539_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_5 ( .D(_00079_ ), .CK(clock ), .Q(\arbiter.clink.mtime [58] ), .QN(_14538_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_50 ( .D(_00080_ ), .CK(clock ), .Q(\arbiter.clink.mtime [13] ), .QN(_14537_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_51 ( .D(_00081_ ), .CK(clock ), .Q(\arbiter.clink.mtime [12] ), .QN(_14536_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_52 ( .D(_00082_ ), .CK(clock ), .Q(\arbiter.clink.mtime [11] ), .QN(_14535_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_53 ( .D(_00083_ ), .CK(clock ), .Q(\arbiter.clink.mtime [10] ), .QN(_14534_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_54 ( .D(_00084_ ), .CK(clock ), .Q(\arbiter.clink.mtime [9] ), .QN(_14533_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_55 ( .D(_00085_ ), .CK(clock ), .Q(\arbiter.clink.mtime [8] ), .QN(_14532_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_56 ( .D(_00086_ ), .CK(clock ), .Q(\arbiter.clink.mtime [7] ), .QN(_14531_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_57 ( .D(_00087_ ), .CK(clock ), .Q(\arbiter.clink.mtime [6] ), .QN(_14530_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_58 ( .D(_00088_ ), .CK(clock ), .Q(\arbiter.clink.mtime [5] ), .QN(_14529_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_59 ( .D(_00089_ ), .CK(clock ), .Q(\arbiter.clink.mtime [4] ), .QN(_14528_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_6 ( .D(_00090_ ), .CK(clock ), .Q(\arbiter.clink.mtime [57] ), .QN(_14527_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_60 ( .D(_00091_ ), .CK(clock ), .Q(\arbiter.clink.mtime [3] ), .QN(_14526_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_61 ( .D(_00092_ ), .CK(clock ), .Q(\arbiter.clink.mtime [2] ), .QN(_14525_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_62 ( .D(_00093_ ), .CK(clock ), .Q(\arbiter.clink.mtime [1] ), .QN(_14524_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_63 ( .D(_00094_ ), .CK(clock ), .Q(\arbiter.clink.mtime [0] ), .QN(\arbiter.clink._mtime_T_1 [0] ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_7 ( .D(_00095_ ), .CK(clock ), .Q(\arbiter.clink.mtime [56] ), .QN(_14523_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_8 ( .D(_00096_ ), .CK(clock ), .Q(\arbiter.clink.mtime [55] ), .QN(_14522_ ) );
DFF_X1 \arbiter.clink.mtime_$_SDFF_PP0__Q_9 ( .D(_00097_ ), .CK(clock ), .Q(\arbiter.clink.mtime [54] ), .QN(_14521_ ) );
DFF_X1 \arbiter.ifu_end_$_SDFF_PP0__Q ( .D(_00098_ ), .CK(clock ), .Q(\arbiter.ifu_end ), .QN(_14520_ ) );
DFF_X1 \arbiter.lsu_end_$_SDFF_PP0__Q ( .D(_00099_ ), .CK(clock ), .Q(\arbiter.lsu_end ), .QN(_14585_ ) );
DFF_X1 \arbiter.state_$_DFF_P__Q ( .D(\arbiter.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\arbiter._io_axi_araddr_T ), .QN(_14586_ ) );
DFF_X1 \arbiter.state_$_DFF_P__Q_1 ( .D(\arbiter.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\arbiter._io_axi_araddr_T_6 ), .QN(_14587_ ) );
DFF_X1 \arbiter.state_$_DFF_P__Q_2 ( .D(\arbiter.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\arbiter._clink_io_axi_araddr_T ), .QN(io_master_wready_$_ANDNOT__B_Y_$_OR__A_B ) );
DFF_X1 \exu.state_$_SDFF_PP0__Q ( .D(_00100_ ), .CK(clock ), .Q(\exu.state ), .QN(_14588_ ) );
DFF_X1 exu_io_in_bits_csr_waddr_$_DFFE_PP__Q ( .D(\idu._io_out_bits_csr_waddr_T_16 [1] ), .CK(_13984_ ), .Q(\exu.io_in_bits_csr_waddr [1] ), .QN(_14584_ ) );
DFF_X1 exu_io_in_bits_csr_waddr_$_DFFE_PP__Q_1 ( .D(\idu._io_out_bits_csr_waddr_T_16 [0] ), .CK(_13984_ ), .Q(\exu.io_in_bits_csr_waddr [0] ), .QN(_14589_ ) );
DFF_X1 exu_io_in_bits_r_add_$_DFFE_PP__Q ( .D(\idu.io_out_bits_add ), .CK(_13984_ ), .Q(\exu.add.io_is ), .QN(_14590_ ) );
DFF_X1 exu_io_in_bits_r_addi_$_DFFE_PP__Q ( .D(\idu.io_out_bits_addi ), .CK(_13984_ ), .Q(\exu.addi.io_is ), .QN(_14591_ ) );
DFF_X1 exu_io_in_bits_r_and_$_DFFE_PP__Q ( .D(\idu.io_out_bits_and ), .CK(_13984_ ), .Q(\exu.and_.io_is ), .QN(_14592_ ) );
DFF_X1 exu_io_in_bits_r_andi_$_DFFE_PP__Q ( .D(\idu.io_out_bits_andi ), .CK(_13984_ ), .Q(\exu.andi.io_is ), .QN(_14593_ ) );
DFF_X1 exu_io_in_bits_r_auipc_$_DFFE_PP__Q ( .D(\idu.io_out_bits_auipc ), .CK(_13984_ ), .Q(\exu.auipc.io_is ), .QN(_14594_ ) );
DFF_X1 exu_io_in_bits_r_beq_$_DFFE_PP__Q ( .D(\idu.io_out_bits_beq ), .CK(_13984_ ), .Q(\exu.beq.io_is ), .QN(_14595_ ) );
DFF_X1 exu_io_in_bits_r_bge_$_DFFE_PP__Q ( .D(\idu.io_out_bits_bge ), .CK(_13984_ ), .Q(\exu.bge.io_is ), .QN(_14596_ ) );
DFF_X1 exu_io_in_bits_r_bgeu_$_DFFE_PP__Q ( .D(\idu.io_out_bits_bgeu ), .CK(_13984_ ), .Q(\exu.bgeu.io_is ), .QN(_14597_ ) );
DFF_X1 exu_io_in_bits_r_blt_$_DFFE_PP__Q ( .D(\idu.io_out_bits_blt ), .CK(_13984_ ), .Q(\exu.blt.io_is ), .QN(_14598_ ) );
DFF_X1 exu_io_in_bits_r_bltu_$_DFFE_PP__Q ( .D(\idu.io_out_bits_bltu ), .CK(_13984_ ), .Q(\exu.bltu.io_is ), .QN(_14599_ ) );
DFF_X1 exu_io_in_bits_r_bne_$_DFFE_PP__Q ( .D(\idu.io_out_bits_bne ), .CK(_13984_ ), .Q(\exu.bne.io_is ), .QN(_14519_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q ( .D(_00101_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [30] ), .QN(\ifu.io_out_bits_pc_$_MUX__Y_13_A_$_MUX__Y_A_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_1 ( .D(_00102_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [28] ), .QN(_14518_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_10 ( .D(_00103_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [12] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_17_A_$_MUX__A_B_$_MUX__B_1_A_$_XOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_NOR__B_Y_$_XOR__A_B ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_11 ( .D(_00104_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [11] ), .QN(_14517_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_12 ( .D(_00105_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [8] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_9_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_13 ( .D(_00106_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [6] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_11_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_14 ( .D(_00107_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [4] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_15 ( .D(_00108_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [3] ), .QN(_14516_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_16 ( .D(_00109_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [29] ), .QN(_14515_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_17 ( .D(_00110_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [26] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_1_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_XOR__Y_B ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_18 ( .D(_00111_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [24] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_9_A_$_MUX__A_B_$_MUX__B_1_A_$_XOR__Y_A_$_NOR__A_Y_$_XOR__A_B ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_19 ( .D(_00112_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [19] ), .QN(_14514_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_2 ( .D(_00113_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [27] ), .QN(_14513_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_20 ( .D(_00114_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [9] ), .QN(_14512_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_21 ( .D(_00115_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [5] ), .QN(_14511_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_22 ( .D(_00116_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [1] ), .QN(_14510_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_23 ( .D(_00117_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [31] ), .QN(_14509_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_24 ( .D(_00118_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [25] ), .QN(_14508_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_25 ( .D(_00119_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [23] ), .QN(_14507_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_26 ( .D(_00120_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [18] ), .QN(_14506_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_27 ( .D(_00121_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [15] ), .QN(_14505_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_28 ( .D(_00122_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [10] ), .QN(_14504_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_29 ( .D(_00123_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [7] ), .QN(_14503_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_3 ( .D(_00124_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [22] ), .QN(_14502_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_30 ( .D(_00125_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [2] ), .QN(_14501_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_31 ( .D(_00126_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [0] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_4 ( .D(_00127_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [21] ), .QN(_14500_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_5 ( .D(_00128_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [20] ), .QN(_14499_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_6 ( .D(_00129_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [17] ), .QN(_14498_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_7 ( .D(_00130_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [16] ), .QN(_14497_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_8 ( .D(_00131_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [14] ), .QN(_14496_ ) );
DFF_X1 exu_io_in_bits_r_csr_rdata_$_SDFFCE_PP0P__Q_9 ( .D(_00132_ ), .CK(_13984_ ), .Q(\exu.csrrs.io_csr_rdata [13] ), .QN(_14600_ ) );
DFF_X1 exu_io_in_bits_r_csrrs_$_DFFE_PP__Q ( .D(\idu.io_out_bits_csrrs ), .CK(_13984_ ), .Q(\exu.csrrs.io_is ), .QN(_14601_ ) );
DFF_X1 exu_io_in_bits_r_csrrw_$_DFFE_PP__Q ( .D(\idu.io_out_bits_csrrw ), .CK(_13984_ ), .Q(\exu.csrrw.io_is ), .QN(_14602_ ) );
DFF_X1 exu_io_in_bits_r_ecall_$_DFFE_PP__Q ( .D(\idu._io_csr_raddr_T_14 [0] ), .CK(_13984_ ), .Q(\exu.ecall.io_is ), .QN(\ifu.io_out_bits_pc_$_MUX__Y_9_A_$_MUX__Y_A_$_OR__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 exu_io_in_bits_r_en_dnpc_$_DFFE_PP__Q ( .D(\idu.io_out_bits_en_dnpc ), .CK(_13984_ ), .Q(\exu.io_in_bits_en_dnpc ), .QN(exu_io_in_bits_r_en_dnpc_$_NOT__A_Y ) );
DFF_X1 exu_io_in_bits_r_fencei_$_DFFE_PP__Q ( .D(\idu.io_out_bits_fencei ), .CK(_13984_ ), .Q(\exu.io_in_bits_fencei ), .QN(_14603_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q ( .D(\idu.io_out_bits_imm [31] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [31] ), .QN(_14604_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_1 ( .D(\idu.io_out_bits_imm [30] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [30] ), .QN(_14605_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_10 ( .D(\idu.io_out_bits_imm [21] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [21] ), .QN(_14606_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_11 ( .D(\idu.io_out_bits_imm [20] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [20] ), .QN(_14607_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_12 ( .D(\idu.io_out_bits_imm [19] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [19] ), .QN(_14608_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_13 ( .D(\idu.io_out_bits_imm [18] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [18] ), .QN(_14609_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_14 ( .D(\idu.io_out_bits_imm [17] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [17] ), .QN(_14610_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_15 ( .D(\idu.io_out_bits_imm [16] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [16] ), .QN(_14611_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_16 ( .D(\idu.io_out_bits_imm [15] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [15] ), .QN(_14612_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_17 ( .D(\idu.io_out_bits_imm [14] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [14] ), .QN(_14613_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_18 ( .D(\idu.io_out_bits_imm [13] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [13] ), .QN(_14614_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_19 ( .D(\idu.io_out_bits_imm [12] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [12] ), .QN(_14615_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_2 ( .D(\idu.io_out_bits_imm [29] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [29] ), .QN(_14616_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_20 ( .D(\idu.io_out_bits_imm [11] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [11] ), .QN(_14617_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_21 ( .D(\idu.io_out_bits_imm [10] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [10] ), .QN(_14618_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_22 ( .D(\idu.io_out_bits_imm [9] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [9] ), .QN(_14619_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_23 ( .D(\idu.io_out_bits_imm [8] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [8] ), .QN(_14620_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_24 ( .D(\idu.io_out_bits_imm [7] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [7] ), .QN(_14621_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_25 ( .D(\idu.io_out_bits_imm [6] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [6] ), .QN(_14622_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_26 ( .D(\idu.io_out_bits_imm [5] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [5] ), .QN(_14623_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_27 ( .D(\idu.io_out_bits_imm [4] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [4] ), .QN(_14624_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_28 ( .D(\idu.io_out_bits_imm [3] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [3] ), .QN(_14625_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_29 ( .D(\idu.io_out_bits_imm [2] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [2] ), .QN(_14626_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_3 ( .D(\idu.io_out_bits_imm [28] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [28] ), .QN(_14627_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_30 ( .D(\idu.io_out_bits_imm [1] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [1] ), .QN(_14628_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_31 ( .D(\idu.io_out_bits_imm [0] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [0] ), .QN(_14629_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_4 ( .D(\idu.io_out_bits_imm [27] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [27] ), .QN(_14630_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_5 ( .D(\idu.io_out_bits_imm [26] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [26] ), .QN(_14631_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_6 ( .D(\idu.io_out_bits_imm [25] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [25] ), .QN(_14632_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_7 ( .D(\idu.io_out_bits_imm [24] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [24] ), .QN(_14633_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_8 ( .D(\idu.io_out_bits_imm [23] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [23] ), .QN(_14634_ ) );
DFF_X1 exu_io_in_bits_r_imm_$_DFFE_PP__Q_9 ( .D(\idu.io_out_bits_imm [22] ), .CK(_13984_ ), .Q(\exu.addi.io_imm [22] ), .QN(_14635_ ) );
DFF_X1 exu_io_in_bits_r_jal_$_DFFE_PP__Q ( .D(\idu.io_out_bits_jal ), .CK(_13984_ ), .Q(\exu.io_in_bits_jal ), .QN(_14636_ ) );
DFF_X1 exu_io_in_bits_r_jalr_$_DFFE_PP__Q ( .D(\idu.io_out_bits_jalr ), .CK(_13984_ ), .Q(\exu.io_in_bits_jalr ), .QN(_14637_ ) );
DFF_X1 exu_io_in_bits_r_lb_$_DFFE_PP__Q ( .D(\idu.io_out_bits_lb ), .CK(_13984_ ), .Q(\exu.io_in_bits_lb ), .QN(_14638_ ) );
DFF_X1 exu_io_in_bits_r_lbu_$_DFFE_PP__Q ( .D(\idu.io_out_bits_lbu ), .CK(_13984_ ), .Q(\exu.io_in_bits_lbu ), .QN(_14639_ ) );
DFF_X1 exu_io_in_bits_r_lh_$_DFFE_PP__Q ( .D(\idu.io_out_bits_lh ), .CK(_13984_ ), .Q(\exu.io_in_bits_lh ), .QN(_14640_ ) );
DFF_X1 exu_io_in_bits_r_lhu_$_DFFE_PP__Q ( .D(\idu.io_out_bits_lhu ), .CK(_13984_ ), .Q(\exu.io_in_bits_lhu ), .QN(_14641_ ) );
DFF_X1 exu_io_in_bits_r_lui_$_DFFE_PP__Q ( .D(\idu.io_out_bits_lui ), .CK(_13984_ ), .Q(\exu.io_in_bits_lui ), .QN(exu_io_in_bits_r_lui_$_NOT__A_Y ) );
DFF_X1 exu_io_in_bits_r_lw_$_DFFE_PP__Q ( .D(\idu.io_out_bits_lw ), .CK(_13984_ ), .Q(\exu.io_in_bits_lw ), .QN(_14642_ ) );
DFF_X1 exu_io_in_bits_r_mret_$_DFFE_PP__Q ( .D(\idu._io_csr_raddr_T_15 [1] ), .CK(_13984_ ), .Q(\exu.io_in_bits_mret ), .QN(_14643_ ) );
DFF_X1 exu_io_in_bits_r_or_$_DFFE_PP__Q ( .D(\idu.io_out_bits_or ), .CK(_13984_ ), .Q(\exu.io_in_bits_or ), .QN(_14644_ ) );
DFF_X1 exu_io_in_bits_r_ori_$_DFFE_PP__Q ( .D(\idu.io_out_bits_ori ), .CK(_13984_ ), .Q(\exu.io_in_bits_ori ), .QN(_14645_ ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q ( .D(\idu.io_in_bits_pc [31] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [31] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_1 ( .D(\idu.io_in_bits_pc [30] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [30] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_1_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_10 ( .D(\idu.io_in_bits_pc [21] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [21] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_10_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_11 ( .D(\idu.io_in_bits_pc [20] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [20] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_11_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_12 ( .D(\idu.io_in_bits_pc [19] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [19] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_12_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_13 ( .D(\idu.io_in_bits_pc [18] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [18] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_13_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_14 ( .D(\idu.io_in_bits_pc [17] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [17] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_14_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_15 ( .D(\idu.io_in_bits_pc [16] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [16] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_15_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_16 ( .D(\idu.io_in_bits_pc [15] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [15] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_16_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_17 ( .D(\idu.io_in_bits_pc [14] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [14] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_17_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_18 ( .D(\idu.io_in_bits_pc [13] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [13] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_18_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_19 ( .D(\idu.io_in_bits_pc [12] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [12] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_19_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_2 ( .D(\idu.io_in_bits_pc [29] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [29] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_2_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_20 ( .D(\idu.io_in_bits_pc [11] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [11] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_20_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_21 ( .D(\idu.io_in_bits_pc [10] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [10] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_21_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_22 ( .D(\idu.io_in_bits_pc [9] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [9] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_22_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_23 ( .D(\idu.io_in_bits_pc [8] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [8] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_23_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_24 ( .D(\idu.io_in_bits_pc [7] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [7] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_24_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_25 ( .D(\idu.io_in_bits_pc [6] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [6] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_25_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_26 ( .D(\idu.io_in_bits_pc [5] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [5] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_26_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_27 ( .D(\idu.io_in_bits_pc [4] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [4] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_27_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_28 ( .D(\idu.io_in_bits_pc [3] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [3] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_28_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_29 ( .D(\idu.io_in_bits_pc [2] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [2] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_29_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_3 ( .D(\idu.io_in_bits_pc [28] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [28] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_3_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_30 ( .D(\idu.io_in_bits_pc [1] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [1] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_MUX__Y_B_$_OR__Y_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_31 ( .D(\idu.io_in_bits_pc [0] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [0] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_4 ( .D(\idu.io_in_bits_pc [27] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [27] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_4_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_5 ( .D(\idu.io_in_bits_pc [26] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [26] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_5_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_6 ( .D(\idu.io_in_bits_pc [25] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [25] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_6_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_7 ( .D(\idu.io_in_bits_pc [24] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [24] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_7_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_8 ( .D(\idu.io_in_bits_pc [23] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [23] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_8_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_pc_$_DFFE_PP__Q_9 ( .D(\idu.io_in_bits_pc [22] ), .CK(_13984_ ), .Q(\exu.auipc.io_rs1_data [22] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_9_A_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_rd_$_DFFE_PP__Q ( .D(\idu.immB [4] ), .CK(_13984_ ), .Q(\exu.io_in_bits_rd [4] ), .QN(_14646_ ) );
DFF_X1 exu_io_in_bits_r_rd_$_DFFE_PP__Q_1 ( .D(\idu.immB [3] ), .CK(_13984_ ), .Q(\exu.io_in_bits_rd [3] ), .QN(_14647_ ) );
DFF_X1 exu_io_in_bits_r_rd_$_DFFE_PP__Q_2 ( .D(\idu.immB [2] ), .CK(_13984_ ), .Q(\exu.io_in_bits_rd [2] ), .QN(_14648_ ) );
DFF_X1 exu_io_in_bits_r_rd_$_DFFE_PP__Q_3 ( .D(\idu.immB [1] ), .CK(_13984_ ), .Q(\exu.io_in_bits_rd [1] ), .QN(_14649_ ) );
DFF_X1 exu_io_in_bits_r_rd_$_DFFE_PP__Q_4 ( .D(\idu.immB [11] ), .CK(_13984_ ), .Q(\exu.io_in_bits_rd [0] ), .QN(_14650_ ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q ( .D(\idu.io_out_bits_rs1_data [31] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [31] ), .QN(\exu.addi._io_rd_T_4_$_NOT__Y_A_$_XNOR__Y_B_$_OR__B_Y_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_1 ( .D(\idu.io_out_bits_rs1_data [30] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [30] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_10 ( .D(\idu.io_out_bits_rs1_data [21] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [21] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_11 ( .D(\idu.io_out_bits_rs1_data [20] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [20] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_12 ( .D(\idu.io_out_bits_rs1_data [19] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [19] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_13 ( .D(\idu.io_out_bits_rs1_data [18] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [18] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_14 ( .D(\idu.io_out_bits_rs1_data [17] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [17] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_15 ( .D(\idu.io_out_bits_rs1_data [16] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [16] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_16 ( .D(\idu.io_out_bits_rs1_data [15] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [15] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_17 ( .D(\idu.io_out_bits_rs1_data [14] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [14] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_18 ( .D(\idu.io_out_bits_rs1_data [13] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [13] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_19 ( .D(\idu.io_out_bits_rs1_data [12] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [12] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_2 ( .D(\idu.io_out_bits_rs1_data [29] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [29] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_20 ( .D(\idu.io_out_bits_rs1_data [11] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [11] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_21 ( .D(\idu.io_out_bits_rs1_data [10] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [10] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_22 ( .D(\idu.io_out_bits_rs1_data [9] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [9] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_23 ( .D(\idu.io_out_bits_rs1_data [8] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [8] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_24 ( .D(\idu.io_out_bits_rs1_data [7] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [7] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_25 ( .D(\idu.io_out_bits_rs1_data [6] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [6] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_26 ( .D(\idu.io_out_bits_rs1_data [5] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [5] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_27 ( .D(\idu.io_out_bits_rs1_data [4] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [4] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_28 ( .D(\idu.io_out_bits_rs1_data [3] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [3] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_29 ( .D(\idu.io_out_bits_rs1_data [2] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [2] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_3 ( .D(\idu.io_out_bits_rs1_data [28] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [28] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_30 ( .D(\idu.io_out_bits_rs1_data [1] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [1] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_31 ( .D(\idu.io_out_bits_rs1_data [0] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [0] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_4 ( .D(\idu.io_out_bits_rs1_data [27] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [27] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_5 ( .D(\idu.io_out_bits_rs1_data [26] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [26] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_6 ( .D(\idu.io_out_bits_rs1_data [25] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [25] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_7 ( .D(\idu.io_out_bits_rs1_data [24] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [24] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_8 ( .D(\idu.io_out_bits_rs1_data [23] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [23] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs1_data_$_DFFE_PP__Q_9 ( .D(\idu.io_out_bits_rs1_data [22] ), .CK(_13984_ ), .Q(\exu.add.io_rs1_data [22] ), .QN(\exu.addi._io_rd_T_4_$_XNOR__Y_A_$_ANDNOT__A_Y_$_MUX__B_A_$_MUX__Y_B_$_NOR__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q ( .D(\idu.io_out_bits_rs2_data [31] ), .CK(_13984_ ), .Q(\exu._GEN_0 [31] ), .QN(_14651_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_1 ( .D(\idu.io_out_bits_rs2_data [30] ), .CK(_13984_ ), .Q(\exu._GEN_0 [30] ), .QN(_14652_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_10 ( .D(\idu.io_out_bits_rs2_data [21] ), .CK(_13984_ ), .Q(\exu._GEN_0 [21] ), .QN(_14653_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_11 ( .D(\idu.io_out_bits_rs2_data [20] ), .CK(_13984_ ), .Q(\exu._GEN_0 [20] ), .QN(_14654_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_12 ( .D(\idu.io_out_bits_rs2_data [19] ), .CK(_13984_ ), .Q(\exu._GEN_0 [19] ), .QN(_14655_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_13 ( .D(\idu.io_out_bits_rs2_data [18] ), .CK(_13984_ ), .Q(\exu._GEN_0 [18] ), .QN(_14656_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_14 ( .D(\idu.io_out_bits_rs2_data [17] ), .CK(_13984_ ), .Q(\exu._GEN_0 [17] ), .QN(_14657_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_15 ( .D(\idu.io_out_bits_rs2_data [16] ), .CK(_13984_ ), .Q(\exu._GEN_0 [16] ), .QN(_14658_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_16 ( .D(\idu.io_out_bits_rs2_data [15] ), .CK(_13984_ ), .Q(\exu._GEN_0 [15] ), .QN(_14659_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_17 ( .D(\idu.io_out_bits_rs2_data [14] ), .CK(_13984_ ), .Q(\exu._GEN_0 [14] ), .QN(_14660_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_18 ( .D(\idu.io_out_bits_rs2_data [13] ), .CK(_13984_ ), .Q(\exu._GEN_0 [13] ), .QN(_14661_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_19 ( .D(\idu.io_out_bits_rs2_data [12] ), .CK(_13984_ ), .Q(\exu._GEN_0 [12] ), .QN(_14662_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_2 ( .D(\idu.io_out_bits_rs2_data [29] ), .CK(_13984_ ), .Q(\exu._GEN_0 [29] ), .QN(_14663_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_20 ( .D(\idu.io_out_bits_rs2_data [11] ), .CK(_13984_ ), .Q(\exu._GEN_0 [11] ), .QN(_14664_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_21 ( .D(\idu.io_out_bits_rs2_data [10] ), .CK(_13984_ ), .Q(\exu._GEN_0 [10] ), .QN(_14665_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_22 ( .D(\idu.io_out_bits_rs2_data [9] ), .CK(_13984_ ), .Q(\exu._GEN_0 [9] ), .QN(_14666_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_23 ( .D(\idu.io_out_bits_rs2_data [8] ), .CK(_13984_ ), .Q(\exu._GEN_0 [8] ), .QN(_14667_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_24 ( .D(\idu.io_out_bits_rs2_data [7] ), .CK(_13984_ ), .Q(\exu._GEN_0 [7] ), .QN(_14668_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_25 ( .D(\idu.io_out_bits_rs2_data [6] ), .CK(_13984_ ), .Q(\exu._GEN_0 [6] ), .QN(_14669_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_26 ( .D(\idu.io_out_bits_rs2_data [5] ), .CK(_13984_ ), .Q(\exu._GEN_0 [5] ), .QN(_14670_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_27 ( .D(\idu.io_out_bits_rs2_data [4] ), .CK(_13984_ ), .Q(\exu._GEN_0 [4] ), .QN(\exu.io_out_bits_wdata_$_MUX__Y_11_B_$_ANDNOT__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_28 ( .D(\idu.io_out_bits_rs2_data [3] ), .CK(_13984_ ), .Q(\exu._GEN_0 [3] ), .QN(\exu.io_out_bits_wdata_$_MUX__Y_12_B_$_ANDNOT__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_29 ( .D(\idu.io_out_bits_rs2_data [2] ), .CK(_13984_ ), .Q(\exu._GEN_0 [2] ), .QN(\exu.io_out_bits_wdata_$_MUX__Y_13_B_$_ANDNOT__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_3 ( .D(\idu.io_out_bits_rs2_data [28] ), .CK(_13984_ ), .Q(\exu._GEN_0 [28] ), .QN(_14671_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_30 ( .D(\idu.io_out_bits_rs2_data [1] ), .CK(_13984_ ), .Q(\exu._GEN_0 [1] ), .QN(\exu.io_out_bits_wdata_$_MUX__Y_14_B_$_ANDNOT__Y_B ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_31 ( .D(\idu.io_out_bits_rs2_data [0] ), .CK(_13984_ ), .Q(\exu._GEN_0 [0] ), .QN(_14672_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_4 ( .D(\idu.io_out_bits_rs2_data [27] ), .CK(_13984_ ), .Q(\exu._GEN_0 [27] ), .QN(_14673_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_5 ( .D(\idu.io_out_bits_rs2_data [26] ), .CK(_13984_ ), .Q(\exu._GEN_0 [26] ), .QN(_14674_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_6 ( .D(\idu.io_out_bits_rs2_data [25] ), .CK(_13984_ ), .Q(\exu._GEN_0 [25] ), .QN(_14675_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_7 ( .D(\idu.io_out_bits_rs2_data [24] ), .CK(_13984_ ), .Q(\exu._GEN_0 [24] ), .QN(_14676_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_8 ( .D(\idu.io_out_bits_rs2_data [23] ), .CK(_13984_ ), .Q(\exu._GEN_0 [23] ), .QN(_14677_ ) );
DFF_X1 exu_io_in_bits_r_rs2_data_$_DFFE_PP__Q_9 ( .D(\idu.io_out_bits_rs2_data [22] ), .CK(_13984_ ), .Q(\exu._GEN_0 [22] ), .QN(_14678_ ) );
DFF_X1 exu_io_in_bits_r_sb_$_DFFE_PP__Q ( .D(\idu.io_out_bits_sb ), .CK(_13984_ ), .Q(\exu.io_in_bits_sb ), .QN(_14679_ ) );
DFF_X1 exu_io_in_bits_r_sh_$_DFFE_PP__Q ( .D(\idu.io_out_bits_sh ), .CK(_13984_ ), .Q(\exu.io_in_bits_sh ), .QN(_14680_ ) );
DFF_X1 exu_io_in_bits_r_shamt_$_DFFE_PP__Q ( .D(\idu.funct7 [0] ), .CK(_13984_ ), .Q(\exu.io_in_bits_shamt [5] ), .QN(_14681_ ) );
DFF_X1 exu_io_in_bits_r_shamt_$_DFFE_PP__Q_1 ( .D(\idu.immI [4] ), .CK(_13984_ ), .Q(\exu.io_in_bits_shamt [4] ), .QN(\exu.io_out_bits_wdata_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_shamt_$_DFFE_PP__Q_2 ( .D(\idu.immI [3] ), .CK(_13984_ ), .Q(\exu.io_in_bits_shamt [3] ), .QN(\exu.io_out_bits_wdata_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_shamt_$_DFFE_PP__Q_3 ( .D(\idu.immI [2] ), .CK(_13984_ ), .Q(\exu.io_in_bits_shamt [2] ), .QN(\exu.io_out_bits_wdata_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_shamt_$_DFFE_PP__Q_4 ( .D(\idu.immI [1] ), .CK(_13984_ ), .Q(\exu.io_in_bits_shamt [1] ), .QN(\exu.io_out_bits_wdata_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__A_B ) );
DFF_X1 exu_io_in_bits_r_shamt_$_DFFE_PP__Q_5 ( .D(\idu.immI [0] ), .CK(_13984_ ), .Q(\exu.io_in_bits_shamt [0] ), .QN(_14682_ ) );
DFF_X1 exu_io_in_bits_r_sll_$_DFFE_PP__Q ( .D(\idu.io_out_bits_sll ), .CK(_13984_ ), .Q(\exu.io_in_bits_sll ), .QN(_14683_ ) );
DFF_X1 exu_io_in_bits_r_slli_$_DFFE_PP__Q ( .D(\idu.io_out_bits_slli ), .CK(_13984_ ), .Q(\exu.io_in_bits_slli ), .QN(_14684_ ) );
DFF_X1 exu_io_in_bits_r_slt_$_DFFE_PP__Q ( .D(\idu.io_out_bits_slt ), .CK(_13984_ ), .Q(\exu.io_in_bits_slt ), .QN(_14685_ ) );
DFF_X1 exu_io_in_bits_r_slti_$_DFFE_PP__Q ( .D(\idu.io_out_bits_slti ), .CK(_13984_ ), .Q(\exu.io_in_bits_slti ), .QN(exu_io_in_bits_r_slti_$_NOT__A_Y ) );
DFF_X1 exu_io_in_bits_r_sltiu_$_DFFE_PP__Q ( .D(\idu.io_out_bits_sltiu ), .CK(_13984_ ), .Q(\exu.io_in_bits_sltiu ), .QN(_14686_ ) );
DFF_X1 exu_io_in_bits_r_sltu_$_DFFE_PP__Q ( .D(\idu.io_out_bits_sltu ), .CK(_13984_ ), .Q(\exu.io_in_bits_sltu ), .QN(_14687_ ) );
DFF_X1 exu_io_in_bits_r_sra_$_DFFE_PP__Q ( .D(\idu.io_out_bits_sra ), .CK(_13984_ ), .Q(\exu.io_in_bits_sra ), .QN(_14688_ ) );
DFF_X1 exu_io_in_bits_r_srai_$_DFFE_PP__Q ( .D(\idu.io_out_bits_srai ), .CK(_13984_ ), .Q(\exu.io_in_bits_srai ), .QN(_14689_ ) );
DFF_X1 exu_io_in_bits_r_srl_$_DFFE_PP__Q ( .D(\idu.io_out_bits_srl ), .CK(_13984_ ), .Q(\exu.io_in_bits_srl ), .QN(_14690_ ) );
DFF_X1 exu_io_in_bits_r_srli_$_DFFE_PP__Q ( .D(\idu.io_out_bits_srli ), .CK(_13984_ ), .Q(\exu.io_in_bits_srli ), .QN(_14691_ ) );
DFF_X1 exu_io_in_bits_r_sub_$_DFFE_PP__Q ( .D(\idu.io_out_bits_sub ), .CK(_13984_ ), .Q(\exu.io_in_bits_sub ), .QN(_14692_ ) );
DFF_X1 exu_io_in_bits_r_sw_$_DFFE_PP__Q ( .D(\idu.io_out_bits_sw ), .CK(_13984_ ), .Q(\exu.io_in_bits_sw ), .QN(_14693_ ) );
DFF_X1 exu_io_in_bits_r_wen_csr_$_DFFE_PP__Q ( .D(\idu.io_out_bits_wen_csr ), .CK(_13984_ ), .Q(\exu.io_in_bits_wen_csr ), .QN(_14694_ ) );
DFF_X1 exu_io_in_bits_r_wen_rd_$_DFFE_PP__Q ( .D(\idu.io_out_bits_wen_rd ), .CK(_13984_ ), .Q(\exu.io_in_bits_wen_rd ), .QN(_14695_ ) );
DFF_X1 exu_io_in_bits_r_xor_$_DFFE_PP__Q ( .D(\idu.io_out_bits_xor ), .CK(_13984_ ), .Q(\exu.io_in_bits_xor ), .QN(_14696_ ) );
DFF_X1 exu_io_in_bits_r_xori_$_DFFE_PP__Q ( .D(\idu.io_out_bits_xori ), .CK(_13984_ ), .Q(\exu.io_in_bits_xori ), .QN(_14495_ ) );
DFF_X1 exu_io_in_valid_REG_$_SDFF_PP0__Q ( .D(_00134_ ), .CK(clock ), .Q(\exu.io_in_valid ), .QN(exu_io_in_valid_REG_$_NOT__A_Y ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q ( .D(_00133_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [31] ), .QN(_14494_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_1 ( .D(_00135_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [30] ), .QN(_14493_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_10 ( .D(_00136_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [21] ), .QN(_14492_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_11 ( .D(_00137_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [20] ), .QN(_14491_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_12 ( .D(_00138_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [19] ), .QN(_14490_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_13 ( .D(_00139_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [18] ), .QN(_14489_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_14 ( .D(_00140_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [17] ), .QN(_14488_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_15 ( .D(_00141_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [16] ), .QN(_14487_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_16 ( .D(_00142_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [15] ), .QN(_14486_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_17 ( .D(_00143_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [14] ), .QN(_14485_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_18 ( .D(_00144_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [13] ), .QN(_14484_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_19 ( .D(_00145_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [12] ), .QN(_14483_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_2 ( .D(_00146_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [29] ), .QN(_14482_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_20 ( .D(_00147_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [11] ), .QN(_14481_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_21 ( .D(_00148_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [10] ), .QN(_14480_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_22 ( .D(_00149_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [9] ), .QN(_14479_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_23 ( .D(_00150_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [8] ), .QN(_14478_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_24 ( .D(_00151_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [7] ), .QN(_14477_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_25 ( .D(_00152_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [6] ), .QN(_14476_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_26 ( .D(_00153_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [5] ), .QN(_14475_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_27 ( .D(_00154_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [4] ), .QN(_14474_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_28 ( .D(_00155_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [3] ), .QN(_14473_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_29 ( .D(_00156_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [2] ), .QN(_14472_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_3 ( .D(_00157_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [28] ), .QN(_14471_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_30 ( .D(_00158_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [1] ), .QN(_14470_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_31 ( .D(_00159_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [0] ), .QN(_14469_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_4 ( .D(_00160_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [27] ), .QN(_14468_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_5 ( .D(_00161_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [26] ), .QN(_14467_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_6 ( .D(_00162_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [25] ), .QN(_14466_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_7 ( .D(_00163_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [24] ), .QN(_14465_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_8 ( .D(_00164_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [23] ), .QN(_14464_ ) );
DFF_X1 \icache.icache_reg_0_0_$_SDFFE_PP0P__Q_9 ( .D(_00165_ ), .CK(_13983_ ), .Q(\icache.icache_reg_0_0 [22] ), .QN(_14463_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q ( .D(_00133_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [31] ), .QN(_14462_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_1 ( .D(_00135_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [30] ), .QN(_14461_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_10 ( .D(_00136_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [21] ), .QN(_14460_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_11 ( .D(_00137_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [20] ), .QN(_14459_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_12 ( .D(_00138_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [19] ), .QN(_14458_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_13 ( .D(_00139_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [18] ), .QN(_14457_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_14 ( .D(_00140_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [17] ), .QN(_14456_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_15 ( .D(_00141_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [16] ), .QN(_14455_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_16 ( .D(_00142_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [15] ), .QN(_14454_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_17 ( .D(_00143_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [14] ), .QN(_14453_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_18 ( .D(_00144_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [13] ), .QN(_14452_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_19 ( .D(_00145_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [12] ), .QN(_14451_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_2 ( .D(_00146_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [29] ), .QN(_14450_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_20 ( .D(_00147_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [11] ), .QN(_14449_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_21 ( .D(_00148_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [10] ), .QN(_14448_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_22 ( .D(_00149_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [9] ), .QN(_14447_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_23 ( .D(_00150_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [8] ), .QN(_14446_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_24 ( .D(_00151_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [7] ), .QN(_14445_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_25 ( .D(_00152_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [6] ), .QN(_14444_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_26 ( .D(_00153_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [5] ), .QN(_14443_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_27 ( .D(_00154_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [4] ), .QN(_14442_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_28 ( .D(_00155_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [3] ), .QN(_14441_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_29 ( .D(_00156_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [2] ), .QN(_14440_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_3 ( .D(_00157_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [28] ), .QN(_14439_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_30 ( .D(_00158_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [1] ), .QN(_14438_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_31 ( .D(_00159_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [0] ), .QN(_14437_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_4 ( .D(_00160_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [27] ), .QN(_14436_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_5 ( .D(_00161_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [26] ), .QN(_14435_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_6 ( .D(_00162_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [25] ), .QN(_14434_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_7 ( .D(_00163_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [24] ), .QN(_14433_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_8 ( .D(_00164_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [23] ), .QN(_14432_ ) );
DFF_X1 \icache.icache_reg_0_1_$_SDFFE_PP0P__Q_9 ( .D(_00165_ ), .CK(_13982_ ), .Q(\icache.icache_reg_0_1 [22] ), .QN(_14431_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q ( .D(_00133_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [31] ), .QN(_14430_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_1 ( .D(_00135_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [30] ), .QN(_14429_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_10 ( .D(_00136_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [21] ), .QN(_14428_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_11 ( .D(_00137_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [20] ), .QN(_14427_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_12 ( .D(_00138_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [19] ), .QN(_14426_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_13 ( .D(_00139_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [18] ), .QN(_14425_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_14 ( .D(_00140_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [17] ), .QN(_14424_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_15 ( .D(_00141_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [16] ), .QN(_14423_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_16 ( .D(_00142_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [15] ), .QN(_14422_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_17 ( .D(_00143_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [14] ), .QN(_14421_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_18 ( .D(_00144_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [13] ), .QN(_14420_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_19 ( .D(_00145_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [12] ), .QN(_14419_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_2 ( .D(_00146_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [29] ), .QN(_14418_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_20 ( .D(_00147_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [11] ), .QN(_14417_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_21 ( .D(_00148_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [10] ), .QN(_14416_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_22 ( .D(_00149_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [9] ), .QN(_14415_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_23 ( .D(_00150_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [8] ), .QN(_14414_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_24 ( .D(_00151_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [7] ), .QN(_14413_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_25 ( .D(_00152_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [6] ), .QN(_14412_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_26 ( .D(_00153_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [5] ), .QN(_14411_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_27 ( .D(_00154_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [4] ), .QN(_14410_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_28 ( .D(_00155_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [3] ), .QN(_14409_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_29 ( .D(_00156_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [2] ), .QN(_14408_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_3 ( .D(_00157_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [28] ), .QN(_14407_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_30 ( .D(_00158_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [1] ), .QN(_14406_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_31 ( .D(_00159_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [0] ), .QN(_14405_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_4 ( .D(_00160_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [27] ), .QN(_14404_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_5 ( .D(_00161_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [26] ), .QN(_14403_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_6 ( .D(_00162_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [25] ), .QN(_14402_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_7 ( .D(_00163_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [24] ), .QN(_14401_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_8 ( .D(_00164_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [23] ), .QN(_14400_ ) );
DFF_X1 \icache.icache_reg_0_2_$_SDFFE_PP0P__Q_9 ( .D(_00165_ ), .CK(_13981_ ), .Q(\icache.icache_reg_0_2 [22] ), .QN(_14399_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q ( .D(_00133_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [31] ), .QN(_14398_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_1 ( .D(_00135_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [30] ), .QN(_14397_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_10 ( .D(_00136_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [21] ), .QN(_14396_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_11 ( .D(_00137_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [20] ), .QN(_14395_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_12 ( .D(_00138_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [19] ), .QN(_14394_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_13 ( .D(_00139_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [18] ), .QN(_14393_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_14 ( .D(_00140_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [17] ), .QN(_14392_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_15 ( .D(_00141_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [16] ), .QN(_14391_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_16 ( .D(_00142_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [15] ), .QN(_14390_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_17 ( .D(_00143_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [14] ), .QN(_14389_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_18 ( .D(_00144_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [13] ), .QN(_14388_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_19 ( .D(_00145_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [12] ), .QN(_14387_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_2 ( .D(_00146_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [29] ), .QN(_14386_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_20 ( .D(_00147_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [11] ), .QN(_14385_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_21 ( .D(_00148_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [10] ), .QN(_14384_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_22 ( .D(_00149_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [9] ), .QN(_14383_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_23 ( .D(_00150_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [8] ), .QN(_14382_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_24 ( .D(_00151_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [7] ), .QN(_14381_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_25 ( .D(_00152_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [6] ), .QN(_14380_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_26 ( .D(_00153_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [5] ), .QN(_14379_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_27 ( .D(_00154_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [4] ), .QN(_14378_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_28 ( .D(_00155_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [3] ), .QN(_14377_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_29 ( .D(_00156_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [2] ), .QN(_14376_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_3 ( .D(_00157_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [28] ), .QN(_14375_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_30 ( .D(_00158_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [1] ), .QN(_14374_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_31 ( .D(_00159_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [0] ), .QN(_14373_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_4 ( .D(_00160_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [27] ), .QN(_14372_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_5 ( .D(_00161_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [26] ), .QN(_14371_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_6 ( .D(_00162_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [25] ), .QN(_14370_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_7 ( .D(_00163_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [24] ), .QN(_14369_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_8 ( .D(_00164_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [23] ), .QN(_14368_ ) );
DFF_X1 \icache.icache_reg_0_3_$_SDFFE_PP0P__Q_9 ( .D(_00165_ ), .CK(_13980_ ), .Q(\icache.icache_reg_0_3 [22] ), .QN(_14367_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q ( .D(_00133_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [31] ), .QN(_14366_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_1 ( .D(_00135_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [30] ), .QN(_14365_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_10 ( .D(_00136_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [21] ), .QN(_14364_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_11 ( .D(_00137_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [20] ), .QN(_14363_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_12 ( .D(_00138_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [19] ), .QN(_14362_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_13 ( .D(_00139_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [18] ), .QN(_14361_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_14 ( .D(_00140_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [17] ), .QN(_14360_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_15 ( .D(_00141_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [16] ), .QN(_14359_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_16 ( .D(_00142_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [15] ), .QN(_14358_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_17 ( .D(_00143_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [14] ), .QN(_14357_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_18 ( .D(_00144_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [13] ), .QN(_14356_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_19 ( .D(_00145_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [12] ), .QN(_14355_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_2 ( .D(_00146_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [29] ), .QN(_14354_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_20 ( .D(_00147_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [11] ), .QN(_14353_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_21 ( .D(_00148_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [10] ), .QN(_14352_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_22 ( .D(_00149_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [9] ), .QN(_14351_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_23 ( .D(_00150_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [8] ), .QN(_14350_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_24 ( .D(_00151_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [7] ), .QN(_14349_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_25 ( .D(_00152_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [6] ), .QN(_14348_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_26 ( .D(_00153_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [5] ), .QN(_14347_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_27 ( .D(_00154_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [4] ), .QN(_14346_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_28 ( .D(_00155_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [3] ), .QN(_14345_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_29 ( .D(_00156_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [2] ), .QN(_14344_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_3 ( .D(_00157_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [28] ), .QN(_14343_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_30 ( .D(_00158_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [1] ), .QN(_14342_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_31 ( .D(_00159_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [0] ), .QN(_14341_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_4 ( .D(_00160_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [27] ), .QN(_14340_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_5 ( .D(_00161_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [26] ), .QN(_14339_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_6 ( .D(_00162_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [25] ), .QN(_14338_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_7 ( .D(_00163_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [24] ), .QN(_14337_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_8 ( .D(_00164_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [23] ), .QN(_14336_ ) );
DFF_X1 \icache.icache_reg_1_0_$_SDFFE_PP0P__Q_9 ( .D(_00165_ ), .CK(_13979_ ), .Q(\icache.icache_reg_1_0 [22] ), .QN(_14335_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q ( .D(_00133_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [31] ), .QN(_14334_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_1 ( .D(_00135_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [30] ), .QN(_14333_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_10 ( .D(_00136_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [21] ), .QN(_14332_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_11 ( .D(_00137_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [20] ), .QN(_14331_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_12 ( .D(_00138_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [19] ), .QN(_14330_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_13 ( .D(_00139_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [18] ), .QN(_14329_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_14 ( .D(_00140_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [17] ), .QN(_14328_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_15 ( .D(_00141_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [16] ), .QN(_14327_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_16 ( .D(_00142_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [15] ), .QN(_14326_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_17 ( .D(_00143_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [14] ), .QN(_14325_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_18 ( .D(_00144_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [13] ), .QN(_14324_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_19 ( .D(_00145_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [12] ), .QN(_14323_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_2 ( .D(_00146_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [29] ), .QN(_14322_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_20 ( .D(_00147_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [11] ), .QN(_14321_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_21 ( .D(_00148_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [10] ), .QN(_14320_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_22 ( .D(_00149_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [9] ), .QN(_14319_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_23 ( .D(_00150_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [8] ), .QN(_14318_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_24 ( .D(_00151_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [7] ), .QN(_14317_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_25 ( .D(_00152_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [6] ), .QN(_14316_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_26 ( .D(_00153_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [5] ), .QN(_14315_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_27 ( .D(_00154_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [4] ), .QN(_14314_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_28 ( .D(_00155_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [3] ), .QN(_14313_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_29 ( .D(_00156_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [2] ), .QN(_14312_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_3 ( .D(_00157_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [28] ), .QN(_14311_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_30 ( .D(_00158_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [1] ), .QN(_14310_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_31 ( .D(_00159_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [0] ), .QN(_14309_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_4 ( .D(_00160_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [27] ), .QN(_14308_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_5 ( .D(_00161_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [26] ), .QN(_14307_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_6 ( .D(_00162_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [25] ), .QN(_14306_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_7 ( .D(_00163_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [24] ), .QN(_14305_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_8 ( .D(_00164_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [23] ), .QN(_14304_ ) );
DFF_X1 \icache.icache_reg_1_1_$_SDFFE_PP0P__Q_9 ( .D(_00165_ ), .CK(_13978_ ), .Q(\icache.icache_reg_1_1 [22] ), .QN(_14303_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q ( .D(_00133_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [31] ), .QN(_14302_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_1 ( .D(_00135_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [30] ), .QN(_14301_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_10 ( .D(_00136_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [21] ), .QN(_14300_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_11 ( .D(_00137_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [20] ), .QN(_14299_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_12 ( .D(_00138_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [19] ), .QN(_14298_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_13 ( .D(_00139_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [18] ), .QN(_14297_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_14 ( .D(_00140_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [17] ), .QN(_14296_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_15 ( .D(_00141_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [16] ), .QN(_14295_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_16 ( .D(_00142_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [15] ), .QN(_14294_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_17 ( .D(_00143_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [14] ), .QN(_14293_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_18 ( .D(_00144_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [13] ), .QN(_14292_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_19 ( .D(_00145_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [12] ), .QN(_14291_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_2 ( .D(_00146_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [29] ), .QN(_14290_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_20 ( .D(_00147_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [11] ), .QN(_14289_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_21 ( .D(_00148_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [10] ), .QN(_14288_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_22 ( .D(_00149_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [9] ), .QN(_14287_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_23 ( .D(_00150_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [8] ), .QN(_14286_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_24 ( .D(_00151_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [7] ), .QN(_14285_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_25 ( .D(_00152_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [6] ), .QN(_14284_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_26 ( .D(_00153_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [5] ), .QN(_14283_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_27 ( .D(_00154_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [4] ), .QN(_14282_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_28 ( .D(_00155_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [3] ), .QN(_14281_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_29 ( .D(_00156_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [2] ), .QN(_14280_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_3 ( .D(_00157_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [28] ), .QN(_14279_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_30 ( .D(_00158_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [1] ), .QN(_14278_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_31 ( .D(_00159_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [0] ), .QN(_14277_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_4 ( .D(_00160_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [27] ), .QN(_14276_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_5 ( .D(_00161_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [26] ), .QN(_14275_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_6 ( .D(_00162_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [25] ), .QN(_14274_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_7 ( .D(_00163_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [24] ), .QN(_14273_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_8 ( .D(_00164_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [23] ), .QN(_14272_ ) );
DFF_X1 \icache.icache_reg_1_2_$_SDFFE_PP0P__Q_9 ( .D(_00165_ ), .CK(_13977_ ), .Q(\icache.icache_reg_1_2 [22] ), .QN(_14271_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q ( .D(_00166_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [31] ), .QN(_14270_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_1 ( .D(_00167_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [30] ), .QN(_14269_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_10 ( .D(_00168_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [21] ), .QN(_14268_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_11 ( .D(_00169_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [20] ), .QN(_14267_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_12 ( .D(_00170_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [19] ), .QN(_14266_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_13 ( .D(_00171_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [18] ), .QN(_14265_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_14 ( .D(_00172_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [17] ), .QN(_14264_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_15 ( .D(_00173_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [16] ), .QN(_14263_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_16 ( .D(_00174_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [15] ), .QN(_14262_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_17 ( .D(_00175_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [14] ), .QN(_14261_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_18 ( .D(_00176_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [13] ), .QN(_14260_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_19 ( .D(_00177_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [12] ), .QN(_14259_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_2 ( .D(_00178_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [29] ), .QN(_14258_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_20 ( .D(_00179_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [11] ), .QN(_14257_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_21 ( .D(_00180_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [10] ), .QN(_14256_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_22 ( .D(_00181_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [9] ), .QN(_14255_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_23 ( .D(_00182_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [8] ), .QN(_14254_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_24 ( .D(_00183_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [7] ), .QN(_14253_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_25 ( .D(_00184_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [6] ), .QN(_14252_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_26 ( .D(_00185_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [5] ), .QN(_14251_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_27 ( .D(_00186_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [4] ), .QN(_14250_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_28 ( .D(_00187_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [3] ), .QN(_14249_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_29 ( .D(_00188_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [2] ), .QN(_14248_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_3 ( .D(_00189_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [28] ), .QN(_14247_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_30 ( .D(_00190_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [1] ), .QN(_14246_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_31 ( .D(_00191_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [0] ), .QN(_14245_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_4 ( .D(_00192_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [27] ), .QN(_14244_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_5 ( .D(_00193_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [26] ), .QN(_14243_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_6 ( .D(_00194_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [25] ), .QN(_14242_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_7 ( .D(_00195_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [24] ), .QN(_14241_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_8 ( .D(_00196_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [23] ), .QN(_14240_ ) );
DFF_X1 \icache.icache_reg_1_3_$_SDFFE_PP0P__Q_9 ( .D(_00197_ ), .CK(_13976_ ), .Q(\icache.icache_reg_1_3 [22] ), .QN(_14239_ ) );
DFF_X1 \icache.offset_buf_$_SDFFE_PP0P__Q ( .D(_00198_ ), .CK(_13975_ ), .Q(\icache.offset_buf [1] ), .QN(_14238_ ) );
DFF_X1 \icache.offset_buf_$_SDFFE_PP0P__Q_1 ( .D(_00199_ ), .CK(_13975_ ), .Q(\icache.offset_buf [0] ), .QN(_14237_ ) );
DFF_X1 \icache.state_$_DFF_P__Q ( .D(\icache.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\icache._icache_reg_T ), .QN(_14698_ ) );
DFF_X1 \icache.state_$_DFF_P__Q_1 ( .D(\icache.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\icache._io_out_arvalid_T_2 ), .QN(_14699_ ) );
DFF_X1 \icache.state_$_DFF_P__Q_2 ( .D(\icache.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\icache._io_out_arvalid_T ), .QN(_14236_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q ( .D(_00200_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [26] ), .QN(_14697_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_1 ( .D(_00201_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [25] ), .QN(_14235_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_10 ( .D(_00202_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [16] ), .QN(_14234_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_11 ( .D(_00203_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [15] ), .QN(_14233_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_12 ( .D(_00204_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [14] ), .QN(_14232_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_13 ( .D(_00205_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [13] ), .QN(_14231_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_14 ( .D(_00206_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [12] ), .QN(_14230_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_15 ( .D(_00207_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [11] ), .QN(_14229_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_16 ( .D(_00208_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [10] ), .QN(_14228_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_17 ( .D(_00209_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [9] ), .QN(_14227_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_18 ( .D(_00210_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [8] ), .QN(_14226_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_19 ( .D(_00211_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [7] ), .QN(_14225_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_2 ( .D(_00212_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [24] ), .QN(_14224_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_20 ( .D(_00213_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [6] ), .QN(_14223_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_21 ( .D(_00214_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [5] ), .QN(_14222_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_22 ( .D(_00215_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [4] ), .QN(_14221_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_23 ( .D(_00216_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [3] ), .QN(_14220_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_24 ( .D(_00217_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [2] ), .QN(_14219_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_25 ( .D(_00218_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [1] ), .QN(_14218_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_26 ( .D(_00219_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [0] ), .QN(_14217_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_3 ( .D(_00220_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [23] ), .QN(_14216_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_4 ( .D(_00221_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [22] ), .QN(_14215_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_5 ( .D(_00222_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [21] ), .QN(_14214_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_6 ( .D(_00223_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [20] ), .QN(_14213_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_7 ( .D(_00224_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [19] ), .QN(_14212_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_8 ( .D(_00225_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [18] ), .QN(_14211_ ) );
DFF_X1 \icache.tag_reg_0_$_SDFFE_PP0P__Q_9 ( .D(_00226_ ), .CK(_13974_ ), .Q(\icache.tag_reg_0 [17] ), .QN(_14210_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q ( .D(_00200_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [26] ), .QN(_14209_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_1 ( .D(_00201_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [25] ), .QN(_14208_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_10 ( .D(_00202_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [16] ), .QN(_14207_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_11 ( .D(_00203_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [15] ), .QN(_14206_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_12 ( .D(_00204_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [14] ), .QN(_14205_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_13 ( .D(_00205_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [13] ), .QN(_14204_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_14 ( .D(_00206_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [12] ), .QN(_14203_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_15 ( .D(_00207_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [11] ), .QN(_14202_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_16 ( .D(_00208_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [10] ), .QN(_14201_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_17 ( .D(_00209_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [9] ), .QN(_14200_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_18 ( .D(_00210_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [8] ), .QN(_14199_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_19 ( .D(_00211_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [7] ), .QN(_14198_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_2 ( .D(_00212_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [24] ), .QN(_14197_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_20 ( .D(_00213_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [6] ), .QN(_14196_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_21 ( .D(_00214_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [5] ), .QN(_14195_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_22 ( .D(_00215_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [4] ), .QN(_14194_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_23 ( .D(_00216_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [3] ), .QN(_14193_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_24 ( .D(_00217_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [2] ), .QN(_14192_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_25 ( .D(_00218_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [1] ), .QN(_14191_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_26 ( .D(_00219_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [0] ), .QN(_14190_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_3 ( .D(_00220_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [23] ), .QN(_14189_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_4 ( .D(_00221_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [22] ), .QN(_14188_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_5 ( .D(_00222_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [21] ), .QN(_14187_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_6 ( .D(_00223_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [20] ), .QN(_14186_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_7 ( .D(_00224_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [19] ), .QN(_14185_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_8 ( .D(_00225_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [18] ), .QN(_14184_ ) );
DFF_X1 \icache.tag_reg_1_$_SDFFE_PP0P__Q_9 ( .D(_00226_ ), .CK(_13973_ ), .Q(\icache.tag_reg_1 [17] ), .QN(_14183_ ) );
DFF_X1 \icache.valid_reg_0_$_SDFFE_PP0P__Q ( .D(_00227_ ), .CK(_13972_ ), .Q(\icache.valid_reg_0 ), .QN(_14182_ ) );
DFF_X1 \icache.valid_reg_1_$_SDFFE_PP0N__Q ( .D(_00227_ ), .CK(_13971_ ), .Q(\icache.valid_reg_1 ), .QN(_14700_ ) );
DFF_X1 \idu.io_out_valid_REG_$_DFF_P__Q ( .D(\idu.io_raw ), .CK(clock ), .Q(\idu.io_out_valid_REG ), .QN(_14702_ ) );
DFF_X1 \idu.rs_reg_$_DFF_P__Q ( .D(\idu.rs_reg_$_DFF_P__Q_D ), .CK(clock ), .Q(\idu.rs_reg ), .QN(_14181_ ) );
DFF_X1 \idu.state_$_SDFF_PP0__Q ( .D(_00228_ ), .CK(clock ), .Q(\idu.state ), .QN(_14703_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q ( .D(\ifu.io_out_bits_inst [31] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [31] ), .QN(_14701_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_1 ( .D(\ifu.io_out_bits_inst [30] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [30] ), .QN(_14704_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_10 ( .D(\ifu.io_out_bits_inst [21] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [21] ), .QN(_14705_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_11 ( .D(\ifu.io_out_bits_inst [20] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [20] ), .QN(_14706_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_12 ( .D(\ifu.io_out_bits_inst [19] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [19] ), .QN(_14707_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_13 ( .D(\ifu.io_out_bits_inst [18] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [18] ), .QN(_14708_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_14 ( .D(\ifu.io_out_bits_inst [17] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [17] ), .QN(_14709_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_15 ( .D(\ifu.io_out_bits_inst [16] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [16] ), .QN(_14710_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_16 ( .D(\ifu.io_out_bits_inst [15] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [15] ), .QN(_14711_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_17 ( .D(\ifu.io_out_bits_inst [14] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [14] ), .QN(_14712_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_18 ( .D(\ifu.io_out_bits_inst [13] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [13] ), .QN(_14713_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_19 ( .D(\ifu.io_out_bits_inst [12] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [12] ), .QN(_14714_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_2 ( .D(\ifu.io_out_bits_inst [29] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [29] ), .QN(_14715_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_20 ( .D(\ifu.io_out_bits_inst [11] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [11] ), .QN(_14716_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_21 ( .D(\ifu.io_out_bits_inst [10] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [10] ), .QN(_14717_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_22 ( .D(\ifu.io_out_bits_inst [9] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [9] ), .QN(_14718_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_23 ( .D(\ifu.io_out_bits_inst [8] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [8] ), .QN(_14719_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_24 ( .D(\ifu.io_out_bits_inst [7] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [7] ), .QN(_14720_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_25 ( .D(\ifu.io_out_bits_inst [6] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [6] ), .QN(_14721_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_26 ( .D(\ifu.io_out_bits_inst [5] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [5] ), .QN(_14722_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_27 ( .D(\ifu.io_out_bits_inst [4] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [4] ), .QN(_14723_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_28 ( .D(\ifu.io_out_bits_inst [3] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [3] ), .QN(_14724_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_29 ( .D(\ifu.io_out_bits_inst [2] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [2] ), .QN(_14725_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_3 ( .D(\ifu.io_out_bits_inst [28] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [28] ), .QN(_14726_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_30 ( .D(\ifu.io_out_bits_inst [1] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [1] ), .QN(_14727_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_31 ( .D(\ifu.io_out_bits_inst [0] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [0] ), .QN(_14728_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_4 ( .D(\ifu.io_out_bits_inst [27] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [27] ), .QN(_14729_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_5 ( .D(\ifu.io_out_bits_inst [26] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [26] ), .QN(_14730_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_6 ( .D(\ifu.io_out_bits_inst [25] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [25] ), .QN(_14731_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_7 ( .D(\ifu.io_out_bits_inst [24] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [24] ), .QN(_14732_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_8 ( .D(\ifu.io_out_bits_inst [23] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [23] ), .QN(_14733_ ) );
DFF_X1 idu_io_in_bits_r_inst_$_DFFE_PN__Q_9 ( .D(\ifu.io_out_bits_inst [22] ), .CK(_13970_ ), .Q(\idu.io_in_bits_inst [22] ), .QN(_14734_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q ( .D(\ifu.io_out_bits_pc [31] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [31] ), .QN(_14735_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_1 ( .D(\ifu.io_out_bits_pc [30] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [30] ), .QN(_14736_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_10 ( .D(\ifu.io_out_bits_pc [21] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [21] ), .QN(_14737_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_11 ( .D(\ifu.io_out_bits_pc [20] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [20] ), .QN(_14738_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_12 ( .D(\ifu.io_out_bits_pc [19] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [19] ), .QN(_14739_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_13 ( .D(\ifu.io_out_bits_pc [18] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [18] ), .QN(_14740_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_14 ( .D(\ifu.io_out_bits_pc [17] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [17] ), .QN(_14741_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_15 ( .D(\ifu.io_out_bits_pc [16] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [16] ), .QN(_14742_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_16 ( .D(\ifu.io_out_bits_pc [15] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [15] ), .QN(_14743_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_17 ( .D(\ifu.io_out_bits_pc [14] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [14] ), .QN(_14744_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_18 ( .D(\ifu.io_out_bits_pc [13] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [13] ), .QN(_14745_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_19 ( .D(\ifu.io_out_bits_pc [12] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [12] ), .QN(_14746_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_2 ( .D(\ifu.io_out_bits_pc [29] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [29] ), .QN(_14747_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_20 ( .D(\ifu.io_out_bits_pc [11] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [11] ), .QN(_14748_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_21 ( .D(\ifu.io_out_bits_pc [10] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [10] ), .QN(_14749_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_22 ( .D(\ifu.io_out_bits_pc [9] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [9] ), .QN(_14750_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_23 ( .D(\ifu.io_out_bits_pc [8] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [8] ), .QN(_14751_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_24 ( .D(\ifu.io_out_bits_pc [7] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [7] ), .QN(_14752_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_25 ( .D(\ifu.io_out_bits_pc [6] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [6] ), .QN(_14753_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_26 ( .D(\ifu.io_out_bits_pc [5] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [5] ), .QN(_14754_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_27 ( .D(\ifu.io_out_bits_pc [4] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [4] ), .QN(_14755_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_28 ( .D(\ifu.io_out_bits_pc [3] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [3] ), .QN(_14756_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_29 ( .D(\ifu.io_out_bits_pc [2] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [2] ), .QN(_14757_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_3 ( .D(\ifu.io_out_bits_pc [28] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [28] ), .QN(_14758_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_30 ( .D(\ifu.io_out_bits_pc [1] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [1] ), .QN(_14759_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_31 ( .D(\ifu.io_out_bits_pc [0] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [0] ), .QN(_14760_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_4 ( .D(\ifu.io_out_bits_pc [27] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [27] ), .QN(_14761_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_5 ( .D(\ifu.io_out_bits_pc [26] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [26] ), .QN(_14762_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_6 ( .D(\ifu.io_out_bits_pc [25] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [25] ), .QN(_14763_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_7 ( .D(\ifu.io_out_bits_pc [24] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [24] ), .QN(_14764_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_8 ( .D(\ifu.io_out_bits_pc [23] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [23] ), .QN(_14765_ ) );
DFF_X1 idu_io_in_bits_r_pc_$_DFFE_PN__Q_9 ( .D(\ifu.io_out_bits_pc [22] ), .CK(_13970_ ), .Q(\idu.io_in_bits_pc [22] ), .QN(_14180_ ) );
DFF_X1 idu_io_in_valid_REG_$_SDFF_PP0__Q ( .D(_00230_ ), .CK(clock ), .Q(\idu.io_in_valid ), .QN(_14178_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q ( .D(_00231_ ), .CK(clock ), .Q(\ifu.inst [31] ), .QN(_14177_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_1 ( .D(_00232_ ), .CK(clock ), .Q(\ifu.inst [30] ), .QN(_14176_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_10 ( .D(_00233_ ), .CK(clock ), .Q(\ifu.inst [21] ), .QN(_14175_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_11 ( .D(_00234_ ), .CK(clock ), .Q(\ifu.inst [20] ), .QN(_14174_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_12 ( .D(_00235_ ), .CK(clock ), .Q(\ifu.inst [19] ), .QN(_14173_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_13 ( .D(_00236_ ), .CK(clock ), .Q(\ifu.inst [18] ), .QN(_14172_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_14 ( .D(_00237_ ), .CK(clock ), .Q(\ifu.inst [17] ), .QN(_14171_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_15 ( .D(_00238_ ), .CK(clock ), .Q(\ifu.inst [16] ), .QN(_14170_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_16 ( .D(_00239_ ), .CK(clock ), .Q(\ifu.inst [15] ), .QN(_14169_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_17 ( .D(_00240_ ), .CK(clock ), .Q(\ifu.inst [14] ), .QN(_14168_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_18 ( .D(_00241_ ), .CK(clock ), .Q(\ifu.inst [13] ), .QN(_14167_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_19 ( .D(_00242_ ), .CK(clock ), .Q(\ifu.inst [12] ), .QN(_14166_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_2 ( .D(_00243_ ), .CK(clock ), .Q(\ifu.inst [29] ), .QN(_14165_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_20 ( .D(_00244_ ), .CK(clock ), .Q(\ifu.inst [11] ), .QN(_14164_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_21 ( .D(_00245_ ), .CK(clock ), .Q(\ifu.inst [10] ), .QN(_14163_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_22 ( .D(_00246_ ), .CK(clock ), .Q(\ifu.inst [9] ), .QN(_14162_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_23 ( .D(_00247_ ), .CK(clock ), .Q(\ifu.inst [8] ), .QN(_14161_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_24 ( .D(_00248_ ), .CK(clock ), .Q(\ifu.inst [7] ), .QN(_14160_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_25 ( .D(_00249_ ), .CK(clock ), .Q(\ifu.inst [6] ), .QN(_14159_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_26 ( .D(_00250_ ), .CK(clock ), .Q(\ifu.inst [5] ), .QN(_14158_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_27 ( .D(_00251_ ), .CK(clock ), .Q(\ifu.inst [4] ), .QN(_14157_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_28 ( .D(_00252_ ), .CK(clock ), .Q(\ifu.inst [3] ), .QN(_14156_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_29 ( .D(_00253_ ), .CK(clock ), .Q(\ifu.inst [2] ), .QN(_14155_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_3 ( .D(_00254_ ), .CK(clock ), .Q(\ifu.inst [28] ), .QN(_14154_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_30 ( .D(_00255_ ), .CK(clock ), .Q(\ifu.inst [1] ), .QN(_14153_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_31 ( .D(_00256_ ), .CK(clock ), .Q(\ifu.inst [0] ), .QN(_14152_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_4 ( .D(_00257_ ), .CK(clock ), .Q(\ifu.inst [27] ), .QN(_14151_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_5 ( .D(_00258_ ), .CK(clock ), .Q(\ifu.inst [26] ), .QN(_14150_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_6 ( .D(_00259_ ), .CK(clock ), .Q(\ifu.inst [25] ), .QN(_14149_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_7 ( .D(_00260_ ), .CK(clock ), .Q(\ifu.inst [24] ), .QN(_14148_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_8 ( .D(_00261_ ), .CK(clock ), .Q(\ifu.inst [23] ), .QN(_14147_ ) );
DFF_X1 \ifu.inst_$_SDFF_PP0__Q_9 ( .D(_00262_ ), .CK(clock ), .Q(\ifu.inst [22] ), .QN(_14146_ ) );
DFF_X1 \ifu.pc_$_SDFFE_PP0P__Q ( .D(_00229_ ), .CK(_13969_ ), .Q(\ifu._pc_T_8 [1] ), .QN(_14179_ ) );
DFF_X1 \ifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00263_ ), .CK(_13969_ ), .Q(\ifu._pc_T_8 [0] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_16_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q ( .D(_00265_ ), .CK(clock ), .Q(\ifu.pc [31] ), .QN(_14145_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_1 ( .D(_00266_ ), .CK(clock ), .Q(\ifu.pc [30] ), .QN(_14144_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_10 ( .D(_00267_ ), .CK(clock ), .Q(\ifu.pc [19] ), .QN(_14143_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_11 ( .D(_00268_ ), .CK(clock ), .Q(\ifu.pc [18] ), .QN(_14142_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_12 ( .D(_00269_ ), .CK(clock ), .Q(\ifu.pc [17] ), .QN(_14141_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_13 ( .D(_00270_ ), .CK(clock ), .Q(\ifu.pc [16] ), .QN(_14140_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_14 ( .D(_00271_ ), .CK(clock ), .Q(\ifu.pc [15] ), .QN(_14139_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_15 ( .D(_00272_ ), .CK(clock ), .Q(\ifu.pc [14] ), .QN(_14138_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_16 ( .D(_00273_ ), .CK(clock ), .Q(\ifu.pc [13] ), .QN(_14137_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_17 ( .D(_00274_ ), .CK(clock ), .Q(\ifu.pc [12] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_5_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_18 ( .D(_00275_ ), .CK(clock ), .Q(\ifu.pc [11] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_6_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_19 ( .D(_00276_ ), .CK(clock ), .Q(\ifu.pc [10] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_7_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_2 ( .D(_00277_ ), .CK(clock ), .Q(\ifu.pc [27] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_20 ( .D(_00278_ ), .CK(clock ), .Q(\ifu.pc [9] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_8_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_21 ( .D(_00279_ ), .CK(clock ), .Q(\ifu.pc [8] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_9_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_22 ( .D(_00280_ ), .CK(clock ), .Q(\ifu.pc [7] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_10_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_23 ( .D(_00281_ ), .CK(clock ), .Q(\ifu.pc [6] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_11_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_24 ( .D(_00282_ ), .CK(clock ), .Q(\ifu.pc [5] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_12_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_25 ( .D(_00283_ ), .CK(clock ), .Q(\ifu.pc [4] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_13_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_26 ( .D(_00284_ ), .CK(clock ), .Q(\ifu.pc [3] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_14_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_27 ( .D(_00285_ ), .CK(clock ), .Q(\ifu.pc [2] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_15_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_3 ( .D(_00286_ ), .CK(clock ), .Q(\ifu.pc [26] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_1_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_4 ( .D(_00287_ ), .CK(clock ), .Q(\ifu.pc [25] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_2_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_5 ( .D(_00288_ ), .CK(clock ), .Q(\ifu.pc [24] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_3_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_6 ( .D(_00289_ ), .CK(clock ), .Q(\ifu.pc [23] ), .QN(\ifu.io_out_bits_pc_$_NOT__Y_4_A_$_MUX__Y_B ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_7 ( .D(_00290_ ), .CK(clock ), .Q(\ifu.pc [22] ), .QN(_14136_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_8 ( .D(_00291_ ), .CK(clock ), .Q(\ifu.pc [21] ), .QN(_14135_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP0__Q_9 ( .D(_00292_ ), .CK(clock ), .Q(\ifu.pc [20] ), .QN(_14134_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP1__Q ( .D(_00293_ ), .CK(clock ), .Q(\ifu.pc [29] ), .QN(_14133_ ) );
DFF_X1 \ifu.pc_$_SDFF_PP1__Q_1 ( .D(_00294_ ), .CK(clock ), .Q(\ifu.pc [28] ), .QN(_14766_ ) );
DFF_X1 \ifu.ren_REG_$_DFF_P__Q ( .D(\ifu.ren_REG_$_DFF_P__Q_D ), .CK(clock ), .Q(\ifu.ren_REG ), .QN(_14132_ ) );
DFF_X1 \ifu.start_$_SDFFE_PP0P__Q ( .D(_00264_ ), .CK(_13968_ ), .Q(\ifu.start [0] ), .QN(\ifu._start_T_2 [0] ) );
DFF_X1 \ifu.start_$_SDFFE_PP1P__Q ( .D(_00295_ ), .CK(_13968_ ), .Q(\ifu.start [1] ), .QN(_14767_ ) );
DFF_X1 \ifu.state_$_DFF_P__Q ( .D(\ifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\ifu.state [2] ), .QN(_14769_ ) );
DFF_X1 \ifu.state_$_DFF_P__Q_1 ( .D(\ifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\ifu.state [1] ), .QN(_14770_ ) );
DFF_X1 \ifu.state_$_DFF_P__Q_2 ( .D(\ifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\ifu.state [0] ), .QN(_14771_ ) );
DFF_X1 \lsu.state_$_DFF_P__Q ( .D(\lsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(io_master_bready ), .QN(_14772_ ) );
DFF_X1 \lsu.state_$_DFF_P__Q_1 ( .D(\lsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\lsu._io_axi_awvalid_T_1 ), .QN(_14773_ ) );
DFF_X1 \lsu.state_$_DFF_P__Q_2 ( .D(\lsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\lsu.state [1] ), .QN(_14774_ ) );
DFF_X1 \lsu.state_$_DFF_P__Q_3 ( .D(\lsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\lsu._io_in_ready_T ), .QN(_14775_ ) );
DFF_X1 lsu_io_in_bits_csr_waddr_$_DFFE_PP__Q ( .D(\exu.io_in_bits_csr_waddr [1] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_waddr [1] ), .QN(_14768_ ) );
DFF_X1 lsu_io_in_bits_csr_waddr_$_DFFE_PP__Q_1 ( .D(\exu.io_in_bits_csr_waddr [0] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_waddr [0] ), .QN(_14776_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q ( .D(\exu.addi._io_rd_T_4 [31] ), .CK(_13967_ ), .Q(\io_master_awaddr [31] ), .QN(_14777_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_1 ( .D(\exu.addi._io_rd_T_4 [30] ), .CK(_13967_ ), .Q(\io_master_awaddr [30] ), .QN(_14778_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_10 ( .D(\exu.addi._io_rd_T_4 [21] ), .CK(_13967_ ), .Q(\io_master_awaddr [21] ), .QN(_14779_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_11 ( .D(\exu.addi._io_rd_T_4 [20] ), .CK(_13967_ ), .Q(\io_master_awaddr [20] ), .QN(_14780_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_12 ( .D(\exu.addi._io_rd_T_4 [19] ), .CK(_13967_ ), .Q(\io_master_awaddr [19] ), .QN(_14781_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_13 ( .D(\exu.addi._io_rd_T_4 [18] ), .CK(_13967_ ), .Q(\io_master_awaddr [18] ), .QN(_14782_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_14 ( .D(\exu.addi._io_rd_T_4 [17] ), .CK(_13967_ ), .Q(\io_master_awaddr [17] ), .QN(_14783_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_15 ( .D(\exu.addi._io_rd_T_4 [16] ), .CK(_13967_ ), .Q(\io_master_awaddr [16] ), .QN(_14784_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_16 ( .D(\exu.addi._io_rd_T_4 [15] ), .CK(_13967_ ), .Q(\io_master_awaddr [15] ), .QN(_14785_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_17 ( .D(\exu.addi._io_rd_T_4 [14] ), .CK(_13967_ ), .Q(\io_master_awaddr [14] ), .QN(_14786_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_18 ( .D(\exu.addi._io_rd_T_4 [13] ), .CK(_13967_ ), .Q(\io_master_awaddr [13] ), .QN(_14787_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_19 ( .D(\exu.addi._io_rd_T_4 [12] ), .CK(_13967_ ), .Q(\io_master_awaddr [12] ), .QN(_14788_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_2 ( .D(\exu.addi._io_rd_T_4 [29] ), .CK(_13967_ ), .Q(\io_master_awaddr [29] ), .QN(_14789_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_20 ( .D(\exu.addi._io_rd_T_4 [11] ), .CK(_13967_ ), .Q(\io_master_awaddr [11] ), .QN(_14790_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_21 ( .D(\exu.addi._io_rd_T_4 [10] ), .CK(_13967_ ), .Q(\io_master_awaddr [10] ), .QN(_14791_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_22 ( .D(\exu.addi._io_rd_T_4 [9] ), .CK(_13967_ ), .Q(\io_master_awaddr [9] ), .QN(_14792_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_23 ( .D(\exu.addi._io_rd_T_4 [8] ), .CK(_13967_ ), .Q(\io_master_awaddr [8] ), .QN(_14793_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_24 ( .D(\exu.addi._io_rd_T_4 [7] ), .CK(_13967_ ), .Q(\io_master_awaddr [7] ), .QN(_14794_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_25 ( .D(\exu.addi._io_rd_T_4 [6] ), .CK(_13967_ ), .Q(\io_master_awaddr [6] ), .QN(_14795_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_26 ( .D(\exu.addi._io_rd_T_4 [5] ), .CK(_13967_ ), .Q(\io_master_awaddr [5] ), .QN(_14796_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_27 ( .D(\exu.addi._io_rd_T_4 [4] ), .CK(_13967_ ), .Q(\io_master_awaddr [4] ), .QN(_14797_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_28 ( .D(\exu.addi._io_rd_T_4 [3] ), .CK(_13967_ ), .Q(\io_master_awaddr [3] ), .QN(_14798_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_29 ( .D(\exu.addi._io_rd_T_4 [2] ), .CK(_13967_ ), .Q(fanout_net_16 ), .QN(_14799_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_3 ( .D(\exu.addi._io_rd_T_4 [28] ), .CK(_13967_ ), .Q(\io_master_awaddr [28] ), .QN(_14800_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_30 ( .D(\exu._io_out_bits_wdata_T_1 [4] ), .CK(_13967_ ), .Q(\io_master_awaddr [1] ), .QN(io_master_wstrb_$_ANDNOT__Y_A ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_31 ( .D(\exu._io_out_bits_wdata_T_1 [3] ), .CK(_13967_ ), .Q(\io_master_awaddr [0] ), .QN(lsu_io_in_bits_r_sb_$_ANDNOT__B_Y_$_ANDNOT__B_A ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_4 ( .D(\exu.addi._io_rd_T_4 [27] ), .CK(_13967_ ), .Q(\io_master_awaddr [27] ), .QN(_14801_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_5 ( .D(\exu.addi._io_rd_T_4 [26] ), .CK(_13967_ ), .Q(\io_master_awaddr [26] ), .QN(_14802_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_6 ( .D(\exu.addi._io_rd_T_4 [25] ), .CK(_13967_ ), .Q(\io_master_awaddr [25] ), .QN(_14803_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_7 ( .D(\exu.addi._io_rd_T_4 [24] ), .CK(_13967_ ), .Q(\io_master_awaddr [24] ), .QN(_14804_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_8 ( .D(\exu.addi._io_rd_T_4 [23] ), .CK(_13967_ ), .Q(\io_master_awaddr [23] ), .QN(_14805_ ) );
DFF_X1 lsu_io_in_bits_r_addr_$_DFFE_PP__Q_9 ( .D(\exu.addi._io_rd_T_4 [22] ), .CK(_13967_ ), .Q(\io_master_awaddr [22] ), .QN(_14806_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q ( .D(\exu.io_out_bits_csr_wdata [31] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [31] ), .QN(_14807_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_1 ( .D(\exu.io_out_bits_csr_wdata [30] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [30] ), .QN(_14808_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_10 ( .D(\exu.io_out_bits_csr_wdata [21] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [21] ), .QN(_14809_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_11 ( .D(\exu.io_out_bits_csr_wdata [20] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [20] ), .QN(_14810_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_12 ( .D(\exu.io_out_bits_csr_wdata [19] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [19] ), .QN(_14811_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_13 ( .D(\exu.io_out_bits_csr_wdata [18] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [18] ), .QN(_14812_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_14 ( .D(\exu.io_out_bits_csr_wdata [17] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [17] ), .QN(_14813_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_15 ( .D(\exu.io_out_bits_csr_wdata [16] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [16] ), .QN(_14814_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_16 ( .D(\exu.io_out_bits_csr_wdata [15] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [15] ), .QN(_14815_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_17 ( .D(\exu.io_out_bits_csr_wdata [14] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [14] ), .QN(_14816_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_18 ( .D(\exu.io_out_bits_csr_wdata [13] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [13] ), .QN(_14817_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_19 ( .D(\exu.io_out_bits_csr_wdata [12] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [12] ), .QN(_14818_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_2 ( .D(\exu.io_out_bits_csr_wdata [29] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [29] ), .QN(_14819_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_20 ( .D(\exu.io_out_bits_csr_wdata [11] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [11] ), .QN(_14820_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_21 ( .D(\exu.io_out_bits_csr_wdata [10] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [10] ), .QN(_14821_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_22 ( .D(\exu.io_out_bits_csr_wdata [9] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [9] ), .QN(_14822_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_23 ( .D(\exu.io_out_bits_csr_wdata [8] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [8] ), .QN(_14823_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_24 ( .D(\exu.io_out_bits_csr_wdata [7] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [7] ), .QN(_14824_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_25 ( .D(\exu.io_out_bits_csr_wdata [6] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [6] ), .QN(_14825_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_26 ( .D(\exu.io_out_bits_csr_wdata [5] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [5] ), .QN(_14826_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_27 ( .D(\exu.io_out_bits_csr_wdata [4] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [4] ), .QN(_14827_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_28 ( .D(\exu.io_out_bits_csr_wdata [3] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [3] ), .QN(_14828_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_29 ( .D(\exu.io_out_bits_csr_wdata [2] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [2] ), .QN(_14829_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_3 ( .D(\exu.io_out_bits_csr_wdata [28] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [28] ), .QN(_14830_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_30 ( .D(\exu.io_out_bits_csr_wdata [1] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [1] ), .QN(_14831_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_31 ( .D(\exu.io_out_bits_csr_wdata [0] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [0] ), .QN(_14832_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_4 ( .D(\exu.io_out_bits_csr_wdata [27] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [27] ), .QN(_14833_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_5 ( .D(\exu.io_out_bits_csr_wdata [26] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [26] ), .QN(_14834_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_6 ( .D(\exu.io_out_bits_csr_wdata [25] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [25] ), .QN(_14835_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_7 ( .D(\exu.io_out_bits_csr_wdata [24] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [24] ), .QN(_14836_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_8 ( .D(\exu.io_out_bits_csr_wdata [23] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [23] ), .QN(_14837_ ) );
DFF_X1 lsu_io_in_bits_r_csr_wdata_$_DFFE_PP__Q_9 ( .D(\exu.io_out_bits_csr_wdata [22] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_csr_wdata [22] ), .QN(_14838_ ) );
DFF_X1 lsu_io_in_bits_r_ecall_$_DFFE_PP__Q ( .D(\exu.ecall.io_is ), .CK(_13967_ ), .Q(\lsu.io_in_bits_ecall ), .QN(_14839_ ) );
DFF_X1 lsu_io_in_bits_r_lb_$_DFFE_PP__Q ( .D(\exu.io_in_bits_lb ), .CK(_13967_ ), .Q(\lsu.io_in_bits_lb ), .QN(_14840_ ) );
DFF_X1 lsu_io_in_bits_r_lbu_$_DFFE_PP__Q ( .D(\exu.io_in_bits_lbu ), .CK(_13967_ ), .Q(\lsu.io_in_bits_lbu ), .QN(_14841_ ) );
DFF_X1 lsu_io_in_bits_r_lh_$_DFFE_PP__Q ( .D(\exu.io_in_bits_lh ), .CK(_13967_ ), .Q(\lsu.io_in_bits_lh ), .QN(_14842_ ) );
DFF_X1 lsu_io_in_bits_r_lhu_$_DFFE_PP__Q ( .D(\exu.io_in_bits_lhu ), .CK(_13967_ ), .Q(\lsu.io_in_bits_lhu ), .QN(_14843_ ) );
DFF_X1 lsu_io_in_bits_r_lw_$_DFFE_PP__Q ( .D(\exu.io_in_bits_lw ), .CK(_13967_ ), .Q(\arbiter.io_lsu_arsize [1] ), .QN(_14844_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q ( .D(\exu.auipc.io_rs1_data [31] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [31] ), .QN(_14845_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_1 ( .D(\exu.auipc.io_rs1_data [30] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [30] ), .QN(_14846_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_10 ( .D(\exu.auipc.io_rs1_data [21] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [21] ), .QN(_14847_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_11 ( .D(\exu.auipc.io_rs1_data [20] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [20] ), .QN(_14848_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_12 ( .D(\exu.auipc.io_rs1_data [19] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [19] ), .QN(_14849_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_13 ( .D(\exu.auipc.io_rs1_data [18] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [18] ), .QN(_14850_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_14 ( .D(\exu.auipc.io_rs1_data [17] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [17] ), .QN(_14851_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_15 ( .D(\exu.auipc.io_rs1_data [16] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [16] ), .QN(_14852_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_16 ( .D(\exu.auipc.io_rs1_data [15] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [15] ), .QN(_14853_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_17 ( .D(\exu.auipc.io_rs1_data [14] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [14] ), .QN(_14854_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_18 ( .D(\exu.auipc.io_rs1_data [13] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [13] ), .QN(_14855_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_19 ( .D(\exu.auipc.io_rs1_data [12] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [12] ), .QN(_14856_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_2 ( .D(\exu.auipc.io_rs1_data [29] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [29] ), .QN(_14857_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_20 ( .D(\exu.auipc.io_rs1_data [11] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [11] ), .QN(_14858_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_21 ( .D(\exu.auipc.io_rs1_data [10] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [10] ), .QN(_14859_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_22 ( .D(\exu.auipc.io_rs1_data [9] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [9] ), .QN(_14860_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_23 ( .D(\exu.auipc.io_rs1_data [8] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [8] ), .QN(_14861_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_24 ( .D(\exu.auipc.io_rs1_data [7] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [7] ), .QN(_14862_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_25 ( .D(\exu.auipc.io_rs1_data [6] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [6] ), .QN(_14863_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_26 ( .D(\exu.auipc.io_rs1_data [5] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [5] ), .QN(_14864_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_27 ( .D(\exu.auipc.io_rs1_data [4] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [4] ), .QN(_14865_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_28 ( .D(\exu.auipc.io_rs1_data [3] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [3] ), .QN(_14866_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_29 ( .D(\exu.auipc.io_rs1_data [2] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [2] ), .QN(_14867_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_3 ( .D(\exu.auipc.io_rs1_data [28] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [28] ), .QN(_14868_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_30 ( .D(\exu.auipc.io_rs1_data [1] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [1] ), .QN(_14869_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_31 ( .D(\exu.auipc.io_rs1_data [0] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [0] ), .QN(_14870_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_4 ( .D(\exu.auipc.io_rs1_data [27] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [27] ), .QN(_14871_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_5 ( .D(\exu.auipc.io_rs1_data [26] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [26] ), .QN(_14872_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_6 ( .D(\exu.auipc.io_rs1_data [25] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [25] ), .QN(_14873_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_7 ( .D(\exu.auipc.io_rs1_data [24] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [24] ), .QN(_14874_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_8 ( .D(\exu.auipc.io_rs1_data [23] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [23] ), .QN(_14875_ ) );
DFF_X1 lsu_io_in_bits_r_pc_$_DFFE_PP__Q_9 ( .D(\exu.auipc.io_rs1_data [22] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_pc [22] ), .QN(_14876_ ) );
DFF_X1 lsu_io_in_bits_r_rd_$_DFFE_PP__Q ( .D(\exu.io_in_bits_rd [4] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd [4] ), .QN(_14877_ ) );
DFF_X1 lsu_io_in_bits_r_rd_$_DFFE_PP__Q_1 ( .D(\exu.io_in_bits_rd [3] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd [3] ), .QN(_14878_ ) );
DFF_X1 lsu_io_in_bits_r_rd_$_DFFE_PP__Q_2 ( .D(\exu.io_in_bits_rd [2] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd [2] ), .QN(_14879_ ) );
DFF_X1 lsu_io_in_bits_r_rd_$_DFFE_PP__Q_3 ( .D(\exu.io_in_bits_rd [1] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd [1] ), .QN(_14880_ ) );
DFF_X1 lsu_io_in_bits_r_rd_$_DFFE_PP__Q_4 ( .D(\exu.io_in_bits_rd [0] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd [0] ), .QN(_14881_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q ( .D(\exu.io_out_bits_rd_wdata [31] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [31] ), .QN(_14882_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_1 ( .D(\exu.io_out_bits_rd_wdata [30] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [30] ), .QN(_14883_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_10 ( .D(\exu.io_out_bits_rd_wdata [21] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [21] ), .QN(_14884_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_11 ( .D(\exu.io_out_bits_rd_wdata [20] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [20] ), .QN(_14885_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_12 ( .D(\exu.io_out_bits_rd_wdata [19] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [19] ), .QN(_14886_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_13 ( .D(\exu.io_out_bits_rd_wdata [18] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [18] ), .QN(_14887_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_14 ( .D(\exu.io_out_bits_rd_wdata [17] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [17] ), .QN(_14888_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_15 ( .D(\exu.io_out_bits_rd_wdata [16] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [16] ), .QN(_14889_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_16 ( .D(\exu.io_out_bits_rd_wdata [15] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [15] ), .QN(_14890_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_17 ( .D(\exu.io_out_bits_rd_wdata [14] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [14] ), .QN(_14891_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_18 ( .D(\exu.io_out_bits_rd_wdata [13] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [13] ), .QN(_14892_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_19 ( .D(\exu.io_out_bits_rd_wdata [12] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [12] ), .QN(_14893_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_2 ( .D(\exu.io_out_bits_rd_wdata [29] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [29] ), .QN(_14894_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_20 ( .D(\exu.io_out_bits_rd_wdata [11] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [11] ), .QN(_14895_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_21 ( .D(\exu.io_out_bits_rd_wdata [10] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [10] ), .QN(_14896_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_22 ( .D(\exu.io_out_bits_rd_wdata [9] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [9] ), .QN(_14897_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_23 ( .D(\exu.io_out_bits_rd_wdata [8] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [8] ), .QN(_14898_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_24 ( .D(\exu.io_out_bits_rd_wdata [7] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [7] ), .QN(_14899_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_25 ( .D(\exu.io_out_bits_rd_wdata [6] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [6] ), .QN(_14900_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_26 ( .D(\exu.io_out_bits_rd_wdata [5] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [5] ), .QN(_14901_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_27 ( .D(\exu.io_out_bits_rd_wdata [4] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [4] ), .QN(_14902_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_28 ( .D(\exu.io_out_bits_rd_wdata [3] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [3] ), .QN(_14903_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_29 ( .D(\exu.io_out_bits_rd_wdata [2] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [2] ), .QN(_14904_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_3 ( .D(\exu.io_out_bits_rd_wdata [28] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [28] ), .QN(_14905_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_30 ( .D(\exu.io_out_bits_rd_wdata [1] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [1] ), .QN(_14906_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_31 ( .D(\exu.io_out_bits_rd_wdata [0] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [0] ), .QN(_14907_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_4 ( .D(\exu.io_out_bits_rd_wdata [27] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [27] ), .QN(_14908_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_5 ( .D(\exu.io_out_bits_rd_wdata [26] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [26] ), .QN(_14909_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_6 ( .D(\exu.io_out_bits_rd_wdata [25] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [25] ), .QN(_14910_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_7 ( .D(\exu.io_out_bits_rd_wdata [24] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [24] ), .QN(_14911_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_8 ( .D(\exu.io_out_bits_rd_wdata [23] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [23] ), .QN(_14912_ ) );
DFF_X1 lsu_io_in_bits_r_rd_wdata_$_DFFE_PP__Q_9 ( .D(\exu.io_out_bits_rd_wdata [22] ), .CK(_13967_ ), .Q(\lsu.io_in_bits_rd_wdata [22] ), .QN(_14913_ ) );
DFF_X1 lsu_io_in_bits_r_ren_$_DFFE_PP__Q ( .D(\exu.io_out_bits_ren ), .CK(_13967_ ), .Q(\lsu.io_in_bits_ren ), .QN(\idu.io_raw_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 lsu_io_in_bits_r_sb_$_DFFE_PP__Q ( .D(\exu.io_in_bits_sb ), .CK(_13967_ ), .Q(\lsu._GEN_1 [0] ), .QN(_14914_ ) );
DFF_X1 lsu_io_in_bits_r_sh_$_DFFE_PP__Q ( .D(\exu.io_in_bits_sh ), .CK(_13967_ ), .Q(\io_master_awsize [0] ), .QN(_14915_ ) );
DFF_X1 lsu_io_in_bits_r_sw_$_DFFE_PP__Q ( .D(\exu.io_in_bits_sw ), .CK(_13967_ ), .Q(\io_master_awsize [1] ), .QN(_14916_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q ( .D(\exu._io_out_bits_wdata_T_2 [31] ), .CK(_13967_ ), .Q(\io_master_wdata [31] ), .QN(_14917_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_1 ( .D(\exu._io_out_bits_wdata_T_2 [30] ), .CK(_13967_ ), .Q(\io_master_wdata [30] ), .QN(_14918_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_10 ( .D(\exu._io_out_bits_wdata_T_2 [21] ), .CK(_13967_ ), .Q(\io_master_wdata [21] ), .QN(_14919_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_11 ( .D(\exu._io_out_bits_wdata_T_2 [20] ), .CK(_13967_ ), .Q(\io_master_wdata [20] ), .QN(_14920_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_12 ( .D(\exu._io_out_bits_wdata_T_2 [19] ), .CK(_13967_ ), .Q(\io_master_wdata [19] ), .QN(_14921_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_13 ( .D(\exu._io_out_bits_wdata_T_2 [18] ), .CK(_13967_ ), .Q(\io_master_wdata [18] ), .QN(_14922_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_14 ( .D(\exu._io_out_bits_wdata_T_2 [17] ), .CK(_13967_ ), .Q(\io_master_wdata [17] ), .QN(_14923_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_15 ( .D(\exu._io_out_bits_wdata_T_2 [16] ), .CK(_13967_ ), .Q(\io_master_wdata [16] ), .QN(_14924_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_2 ( .D(\exu._io_out_bits_wdata_T_2 [29] ), .CK(_13967_ ), .Q(\io_master_wdata [29] ), .QN(_14925_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_3 ( .D(\exu._io_out_bits_wdata_T_2 [28] ), .CK(_13967_ ), .Q(\io_master_wdata [28] ), .QN(_14926_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_4 ( .D(\exu._io_out_bits_wdata_T_2 [27] ), .CK(_13967_ ), .Q(\io_master_wdata [27] ), .QN(_14927_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_5 ( .D(\exu._io_out_bits_wdata_T_2 [26] ), .CK(_13967_ ), .Q(\io_master_wdata [26] ), .QN(_14928_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_6 ( .D(\exu._io_out_bits_wdata_T_2 [25] ), .CK(_13967_ ), .Q(\io_master_wdata [25] ), .QN(_14929_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_7 ( .D(\exu._io_out_bits_wdata_T_2 [24] ), .CK(_13967_ ), .Q(\io_master_wdata [24] ), .QN(_14930_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_8 ( .D(\exu._io_out_bits_wdata_T_2 [23] ), .CK(_13967_ ), .Q(\io_master_wdata [23] ), .QN(_14931_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_DFFE_PP__Q_9 ( .D(\exu._io_out_bits_wdata_T_2 [22] ), .CK(_13967_ ), .Q(\io_master_wdata [22] ), .QN(_14131_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q ( .D(_00296_ ), .CK(_13967_ ), .Q(\io_master_wdata [15] ), .QN(_14130_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_1 ( .D(_00297_ ), .CK(_13967_ ), .Q(\io_master_wdata [14] ), .QN(_14129_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_10 ( .D(_00298_ ), .CK(_13967_ ), .Q(\io_master_wdata [5] ), .QN(_14128_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_11 ( .D(_00299_ ), .CK(_13967_ ), .Q(\io_master_wdata [4] ), .QN(_14127_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_12 ( .D(_00300_ ), .CK(_13967_ ), .Q(\io_master_wdata [3] ), .QN(_14126_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_13 ( .D(_00301_ ), .CK(_13967_ ), .Q(\io_master_wdata [2] ), .QN(_14125_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_14 ( .D(_00302_ ), .CK(_13967_ ), .Q(\io_master_wdata [1] ), .QN(_14124_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_15 ( .D(_00303_ ), .CK(_13967_ ), .Q(\io_master_wdata [0] ), .QN(_14123_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_2 ( .D(_00304_ ), .CK(_13967_ ), .Q(\io_master_wdata [13] ), .QN(_14122_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_3 ( .D(_00305_ ), .CK(_13967_ ), .Q(\io_master_wdata [12] ), .QN(_14121_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_4 ( .D(_00306_ ), .CK(_13967_ ), .Q(\io_master_wdata [11] ), .QN(_14120_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_5 ( .D(_00307_ ), .CK(_13967_ ), .Q(\io_master_wdata [10] ), .QN(_14119_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_6 ( .D(_00308_ ), .CK(_13967_ ), .Q(\io_master_wdata [9] ), .QN(_14118_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_7 ( .D(_00309_ ), .CK(_13967_ ), .Q(\io_master_wdata [8] ), .QN(_14117_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_8 ( .D(_00310_ ), .CK(_13967_ ), .Q(\io_master_wdata [7] ), .QN(_14116_ ) );
DFF_X1 lsu_io_in_bits_r_wdata_$_SDFFCE_PP0P__Q_9 ( .D(_00311_ ), .CK(_13967_ ), .Q(\io_master_wdata [6] ), .QN(_14932_ ) );
DFF_X1 lsu_io_in_bits_r_wen_$_DFFE_PP__Q ( .D(\exu.io_out_bits_wen ), .CK(_13967_ ), .Q(\lsu.io_in_bits_wen ), .QN(_14933_ ) );
DFF_X1 lsu_io_in_bits_r_wen_csr_$_DFFE_PP__Q ( .D(\exu.io_in_bits_wen_csr ), .CK(_13967_ ), .Q(\lsu.io_in_bits_wen_csr ), .QN(_14934_ ) );
DFF_X1 lsu_io_in_bits_r_wen_rd_$_DFFE_PP__Q ( .D(\exu.io_in_bits_wen_rd ), .CK(_13967_ ), .Q(\lsu.io_in_bits_wen_rd ), .QN(_14115_ ) );
DFF_X1 lsu_io_in_valid_REG_$_SDFF_PP0__Q ( .D(_00312_ ), .CK(clock ), .Q(\lsu.io_in_valid ), .QN(_14113_ ) );
DFF_X1 \wbu.csr_0_$_SDFFE_PP0P__Q ( .D(\ifu.ren_REG_$_DFF_P__Q_D_$_NAND__Y_B ), .CK(_13966_ ), .Q(\wbu.csr_0 [0] ), .QN(_14114_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q ( .D(_00313_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [31] ), .QN(_14112_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_1 ( .D(_00314_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [30] ), .QN(_14111_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_10 ( .D(_00315_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [21] ), .QN(_14110_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_11 ( .D(_00316_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [20] ), .QN(_14109_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_12 ( .D(_00317_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [19] ), .QN(_14108_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_13 ( .D(_00318_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [18] ), .QN(_14107_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_14 ( .D(_00319_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [17] ), .QN(_14106_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_15 ( .D(_00320_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [16] ), .QN(_14105_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_16 ( .D(_00321_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [15] ), .QN(_14104_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_17 ( .D(_00322_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [14] ), .QN(_14103_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_18 ( .D(_00323_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [13] ), .QN(_14102_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_19 ( .D(_00324_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [12] ), .QN(_14101_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_2 ( .D(_00325_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [29] ), .QN(_14100_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_20 ( .D(_00326_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [11] ), .QN(_14099_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_21 ( .D(_00327_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [10] ), .QN(_14098_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_22 ( .D(_00328_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [9] ), .QN(_14097_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_23 ( .D(_00329_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [8] ), .QN(_14096_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_24 ( .D(_00330_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [7] ), .QN(_14095_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_25 ( .D(_00331_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [6] ), .QN(_14094_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_26 ( .D(_00332_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [5] ), .QN(_14093_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_27 ( .D(_00333_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [4] ), .QN(_14092_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_28 ( .D(_00334_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [3] ), .QN(_14091_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_29 ( .D(_00335_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [2] ), .QN(_14090_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_3 ( .D(_00336_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [28] ), .QN(_14089_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_30 ( .D(_00337_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [1] ), .QN(_14088_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_31 ( .D(_00338_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [0] ), .QN(_14087_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_4 ( .D(_00339_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [27] ), .QN(_14086_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_5 ( .D(_00340_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [26] ), .QN(_14085_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_6 ( .D(_00341_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [25] ), .QN(_14084_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_7 ( .D(_00342_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [24] ), .QN(_14083_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_8 ( .D(_00343_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [23] ), .QN(_14082_ ) );
DFF_X1 \wbu.csr_1_$_SDFFE_PP0N__Q_9 ( .D(_00344_ ), .CK(_13965_ ), .Q(\wbu._GEN_135 [22] ), .QN(_14081_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q ( .D(_00313_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [31] ), .QN(_14080_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_1 ( .D(_00314_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [30] ), .QN(_14079_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_10 ( .D(_00315_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [21] ), .QN(_14078_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_11 ( .D(_00316_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [20] ), .QN(_14077_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_12 ( .D(_00317_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [19] ), .QN(_14076_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_13 ( .D(_00318_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [18] ), .QN(_14075_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_14 ( .D(_00319_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [17] ), .QN(_14074_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_15 ( .D(_00320_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [16] ), .QN(_14073_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_16 ( .D(_00321_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [15] ), .QN(_14072_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_17 ( .D(_00322_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [14] ), .QN(_14071_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_18 ( .D(_00323_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [13] ), .QN(_14070_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_19 ( .D(_00324_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [12] ), .QN(_14069_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_2 ( .D(_00325_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [29] ), .QN(_14068_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_20 ( .D(_00326_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [11] ), .QN(_14067_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_21 ( .D(_00327_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [10] ), .QN(_14066_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_22 ( .D(_00328_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [9] ), .QN(_14065_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_23 ( .D(_00329_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [8] ), .QN(_14064_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_24 ( .D(_00330_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [7] ), .QN(_14063_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_25 ( .D(_00331_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [6] ), .QN(_14062_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_26 ( .D(_00332_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [5] ), .QN(_14061_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_27 ( .D(_00333_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [4] ), .QN(_14060_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_28 ( .D(_00334_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [3] ), .QN(_14059_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_29 ( .D(_00335_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [2] ), .QN(_14058_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_3 ( .D(_00336_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [28] ), .QN(_14057_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_30 ( .D(_00337_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [1] ), .QN(_14056_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_31 ( .D(_00338_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [0] ), .QN(_14055_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_4 ( .D(_00339_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [27] ), .QN(_14054_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_5 ( .D(_00340_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [26] ), .QN(_14053_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_6 ( .D(_00341_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [25] ), .QN(_14052_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_7 ( .D(_00342_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [24] ), .QN(_14051_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_8 ( .D(_00343_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [23] ), .QN(_14050_ ) );
DFF_X1 \wbu.csr_2_$_SDFFE_PP0P__Q_9 ( .D(_00344_ ), .CK(_13964_ ), .Q(\wbu.csr_2 [22] ), .QN(_14049_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q ( .D(_00314_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [30] ), .QN(_14048_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_1 ( .D(_00325_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [29] ), .QN(_14047_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_10 ( .D(_00316_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [20] ), .QN(_14046_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_11 ( .D(_00317_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [19] ), .QN(_14045_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_12 ( .D(_00318_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [18] ), .QN(_14044_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_13 ( .D(_00319_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [17] ), .QN(_14043_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_14 ( .D(_00320_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [16] ), .QN(_14042_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_15 ( .D(_00321_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [15] ), .QN(_14041_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_16 ( .D(_00322_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [14] ), .QN(_14040_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_17 ( .D(_00323_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [13] ), .QN(_14039_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_18 ( .D(_00324_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [12] ), .QN(_14038_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_19 ( .D(_00326_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [11] ), .QN(_14037_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_2 ( .D(_00336_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [28] ), .QN(_14036_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_20 ( .D(_00327_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [10] ), .QN(_14035_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_21 ( .D(_00328_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [9] ), .QN(_14034_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_22 ( .D(_00329_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [8] ), .QN(_14033_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_23 ( .D(_00330_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [7] ), .QN(_14032_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_24 ( .D(_00331_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [6] ), .QN(_14031_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_25 ( .D(_00332_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [5] ), .QN(_14030_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_26 ( .D(_00333_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [4] ), .QN(_14029_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_27 ( .D(_00334_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [3] ), .QN(_14028_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_28 ( .D(_00335_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [2] ), .QN(_14027_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_29 ( .D(_00337_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [1] ), .QN(_14026_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_3 ( .D(_00339_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [27] ), .QN(_14025_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_30 ( .D(_00338_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [0] ), .QN(_14024_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_4 ( .D(_00340_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [26] ), .QN(_14023_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_5 ( .D(_00341_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [25] ), .QN(_14022_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_6 ( .D(_00342_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [24] ), .QN(_14021_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_7 ( .D(_00343_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [23] ), .QN(_14020_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_8 ( .D(_00344_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [22] ), .QN(_14019_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP0P__Q_9 ( .D(_00315_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [21] ), .QN(_14018_ ) );
DFF_X1 \wbu.csr_3_$_SDFFE_PP1P__Q ( .D(_00345_ ), .CK(_13963_ ), .Q(\wbu.csr_3 [31] ), .QN(_14017_ ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [0] ), .QN(_14016_ ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_10_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13962_ ), .Q(\wbu.rf_10 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [0] ), .QN(_14015_ ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_11_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13961_ ), .Q(\wbu.rf_11 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [0] ), .QN(_14014_ ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_12_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13960_ ), .Q(\wbu.rf_12 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [0] ), .QN(_14013_ ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_13_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13959_ ), .Q(\wbu.rf_13 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [0] ), .QN(_14012_ ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_14_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13958_ ), .Q(\wbu.rf_14 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [0] ), .QN(_14011_ ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_15_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13957_ ), .Q(\wbu.rf_15 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [0] ), .QN(_14010_ ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_16_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13956_ ), .Q(\wbu.rf_16 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [0] ), .QN(_14009_ ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_17_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13955_ ), .Q(\wbu.rf_17 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [0] ), .QN(_14008_ ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_18_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13954_ ), .Q(\wbu.rf_18 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [0] ), .QN(_14007_ ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_19_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13953_ ), .Q(\wbu.rf_19 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q ( .D(_00346_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_1 ( .D(_00347_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_10 ( .D(_00348_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_11 ( .D(_00349_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_12 ( .D(_00350_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_13 ( .D(_00351_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_14 ( .D(_00352_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_15 ( .D(_00353_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_16 ( .D(_00354_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_17 ( .D(_00355_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_18 ( .D(_00356_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_19 ( .D(_00357_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_2 ( .D(_00358_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_20 ( .D(_00359_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_21 ( .D(_00360_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_22 ( .D(_00361_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_23 ( .D(_00362_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_24 ( .D(_00363_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_25 ( .D(_00364_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_26 ( .D(_00365_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_27 ( .D(_00366_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_28 ( .D(_00367_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_29 ( .D(_00368_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_3 ( .D(_00369_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_30 ( .D(_00370_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_31 ( .D(_00371_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [0] ), .QN(_14006_ ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_4 ( .D(_00372_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_5 ( .D(_00373_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_6 ( .D(_00374_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_7 ( .D(_00375_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_8 ( .D(_00376_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_1_$_SDFFE_PP0N__Q_9 ( .D(_00377_ ), .CK(_13952_ ), .Q(\wbu._GEN_71 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [0] ), .QN(_14005_ ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_20_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13951_ ), .Q(\wbu.rf_20 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [0] ), .QN(_14004_ ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_21_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13950_ ), .Q(\wbu.rf_21 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [0] ), .QN(_14003_ ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_22_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13949_ ), .Q(\wbu.rf_22 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [0] ), .QN(_14002_ ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_23_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13948_ ), .Q(\wbu.rf_23 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [0] ), .QN(_14001_ ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_24_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13947_ ), .Q(\wbu.rf_24 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [0] ), .QN(_14000_ ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_25_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13946_ ), .Q(\wbu.rf_25 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [0] ), .QN(_13999_ ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_26_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13945_ ), .Q(\wbu.rf_26 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [0] ), .QN(_13998_ ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_27_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13944_ ), .Q(\wbu.rf_27 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [0] ), .QN(_13997_ ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_28_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13943_ ), .Q(\wbu.rf_28 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [0] ), .QN(_13996_ ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_29_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13942_ ), .Q(\wbu.rf_29 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [0] ), .QN(_13995_ ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_2_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13941_ ), .Q(\wbu.rf_2 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [0] ), .QN(_13994_ ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_30_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13940_ ), .Q(\wbu.rf_30 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q ( .D(_00378_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_1 ( .D(_00379_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_10 ( .D(_00380_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_11 ( .D(_00381_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_12 ( .D(_00382_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_13 ( .D(_00383_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_14 ( .D(_00384_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_15 ( .D(_00385_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_16 ( .D(_00386_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_17 ( .D(_00387_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_18 ( .D(_00388_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_19 ( .D(_00389_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_2 ( .D(_00390_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_20 ( .D(_00391_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_21 ( .D(_00392_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_22 ( .D(_00393_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_23 ( .D(_00394_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_24 ( .D(_00395_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_25 ( .D(_00396_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_26 ( .D(_00397_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_27 ( .D(_00398_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_28 ( .D(_00399_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_29 ( .D(_00400_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_3 ( .D(_00401_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_30 ( .D(_00402_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_31 ( .D(_00403_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [0] ), .QN(_13993_ ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_4 ( .D(_00404_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_5 ( .D(_00405_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_6 ( .D(_00406_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_7 ( .D(_00407_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_8 ( .D(_00408_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_31_$_SDFFE_PP0P__Q_9 ( .D(_00409_ ), .CK(_13939_ ), .Q(\wbu.rf_31 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [0] ), .QN(_13992_ ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_3_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13938_ ), .Q(\wbu.rf_3 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [0] ), .QN(_13991_ ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_4_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13937_ ), .Q(\wbu.rf_4 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [0] ), .QN(_13990_ ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_5_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13936_ ), .Q(\wbu.rf_5 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [0] ), .QN(_13989_ ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_6_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13935_ ), .Q(\wbu.rf_6 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [0] ), .QN(_13988_ ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_7_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13934_ ), .Q(\wbu.rf_7 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [0] ), .QN(_13987_ ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_8_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13933_ ), .Q(\wbu.rf_8 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q ( .D(_00346_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [31] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_1 ( .D(_00347_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [30] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_1_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_10 ( .D(_00348_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [21] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_10_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_11 ( .D(_00349_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [20] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_11_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_12 ( .D(_00350_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [19] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_12_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_13 ( .D(_00351_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [18] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_13_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_14 ( .D(_00352_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [17] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_14_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_15 ( .D(_00353_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [16] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_15_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_16 ( .D(_00354_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [15] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_16_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_17 ( .D(_00355_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [14] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_17_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_18 ( .D(_00356_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [13] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_18_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_19 ( .D(_00357_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [12] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_19_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_2 ( .D(_00358_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [29] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_2_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_20 ( .D(_00359_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [11] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_20_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_21 ( .D(_00360_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [10] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_21_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_22 ( .D(_00361_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [9] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_22_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_23 ( .D(_00362_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [8] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_23_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_24 ( .D(_00363_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [7] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_24_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_25 ( .D(_00364_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [6] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_25_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_26 ( .D(_00365_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [5] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_26_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_27 ( .D(_00366_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [4] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_27_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_28 ( .D(_00367_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [3] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_28_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_29 ( .D(_00368_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [2] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_29_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_3 ( .D(_00369_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [28] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_3_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_30 ( .D(_00370_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [1] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_30_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_31 ( .D(_00371_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [0] ), .QN(_13986_ ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_4 ( .D(_00372_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [27] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_4_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_5 ( .D(_00373_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [26] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_5_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_6 ( .D(_00374_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [25] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_6_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_7 ( .D(_00375_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [24] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_7_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_8 ( .D(_00376_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [23] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_8_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \wbu.rf_9_$_SDFFE_PP0P__Q_9 ( .D(_00377_ ), .CK(_13932_ ), .Q(\wbu.rf_9 [22] ), .QN(idu_io_out_bits_rs2_data_$_MUX__Y_9_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 wbu_io_in_bits_csr_waddr_$_DFFE_PN__Q ( .D(\lsu.io_in_bits_csr_waddr [1] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_waddr [1] ), .QN(_14935_ ) );
DFF_X1 wbu_io_in_bits_csr_waddr_$_DFFE_PN__Q_1 ( .D(\lsu.io_in_bits_csr_waddr [0] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_waddr [0] ), .QN(_14936_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q ( .D(\lsu.io_in_bits_csr_wdata [31] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [31] ), .QN(_14937_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_1 ( .D(\lsu.io_in_bits_csr_wdata [30] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [30] ), .QN(_14938_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_10 ( .D(\lsu.io_in_bits_csr_wdata [21] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [21] ), .QN(_14939_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_11 ( .D(\lsu.io_in_bits_csr_wdata [20] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [20] ), .QN(_14940_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_12 ( .D(\lsu.io_in_bits_csr_wdata [19] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [19] ), .QN(_14941_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_13 ( .D(\lsu.io_in_bits_csr_wdata [18] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [18] ), .QN(_14942_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_14 ( .D(\lsu.io_in_bits_csr_wdata [17] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [17] ), .QN(_14943_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_15 ( .D(\lsu.io_in_bits_csr_wdata [16] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [16] ), .QN(_14944_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_16 ( .D(\lsu.io_in_bits_csr_wdata [15] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [15] ), .QN(_14945_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_17 ( .D(\lsu.io_in_bits_csr_wdata [14] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [14] ), .QN(_14946_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_18 ( .D(\lsu.io_in_bits_csr_wdata [13] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [13] ), .QN(_14947_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_19 ( .D(\lsu.io_in_bits_csr_wdata [12] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [12] ), .QN(_14948_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_2 ( .D(\lsu.io_in_bits_csr_wdata [29] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [29] ), .QN(_14949_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_20 ( .D(\lsu.io_in_bits_csr_wdata [11] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [11] ), .QN(_14950_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_21 ( .D(\lsu.io_in_bits_csr_wdata [10] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [10] ), .QN(_14951_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_22 ( .D(\lsu.io_in_bits_csr_wdata [9] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [9] ), .QN(_14952_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_23 ( .D(\lsu.io_in_bits_csr_wdata [8] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [8] ), .QN(_14953_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_24 ( .D(\lsu.io_in_bits_csr_wdata [7] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [7] ), .QN(_14954_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_25 ( .D(\lsu.io_in_bits_csr_wdata [6] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [6] ), .QN(_14955_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_26 ( .D(\lsu.io_in_bits_csr_wdata [5] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [5] ), .QN(_14956_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_27 ( .D(\lsu.io_in_bits_csr_wdata [4] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [4] ), .QN(_14957_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_28 ( .D(\lsu.io_in_bits_csr_wdata [3] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [3] ), .QN(_14958_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_29 ( .D(\lsu.io_in_bits_csr_wdata [2] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [2] ), .QN(_14959_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_3 ( .D(\lsu.io_in_bits_csr_wdata [28] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [28] ), .QN(_14960_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_30 ( .D(\lsu.io_in_bits_csr_wdata [1] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [1] ), .QN(_14961_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_31 ( .D(\lsu.io_in_bits_csr_wdata [0] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [0] ), .QN(_14962_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_4 ( .D(\lsu.io_in_bits_csr_wdata [27] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [27] ), .QN(_14963_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_5 ( .D(\lsu.io_in_bits_csr_wdata [26] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [26] ), .QN(_14964_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_6 ( .D(\lsu.io_in_bits_csr_wdata [25] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [25] ), .QN(_14965_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_7 ( .D(\lsu.io_in_bits_csr_wdata [24] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [24] ), .QN(_14966_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_8 ( .D(\lsu.io_in_bits_csr_wdata [23] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [23] ), .QN(_14967_ ) );
DFF_X1 wbu_io_in_bits_r_csr_wdata_$_DFFE_PN__Q_9 ( .D(\lsu.io_in_bits_csr_wdata [22] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_csr_wdata [22] ), .QN(_14968_ ) );
DFF_X1 wbu_io_in_bits_r_ecall_$_DFFE_PN__Q ( .D(\lsu.io_in_bits_ecall ), .CK(_13931_ ), .Q(\wbu.io_in_bits_ecall ), .QN(_14969_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q ( .D(\lsu.io_in_bits_pc [31] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [31] ), .QN(_14970_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_1 ( .D(\lsu.io_in_bits_pc [30] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [30] ), .QN(_14971_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_10 ( .D(\lsu.io_in_bits_pc [21] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [21] ), .QN(_14972_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_11 ( .D(\lsu.io_in_bits_pc [20] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [20] ), .QN(_14973_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_12 ( .D(\lsu.io_in_bits_pc [19] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [19] ), .QN(_14974_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_13 ( .D(\lsu.io_in_bits_pc [18] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [18] ), .QN(_14975_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_14 ( .D(\lsu.io_in_bits_pc [17] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [17] ), .QN(_14976_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_15 ( .D(\lsu.io_in_bits_pc [16] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [16] ), .QN(_14977_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_16 ( .D(\lsu.io_in_bits_pc [15] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [15] ), .QN(_14978_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_17 ( .D(\lsu.io_in_bits_pc [14] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [14] ), .QN(_14979_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_18 ( .D(\lsu.io_in_bits_pc [13] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [13] ), .QN(_14980_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_19 ( .D(\lsu.io_in_bits_pc [12] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [12] ), .QN(_14981_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_2 ( .D(\lsu.io_in_bits_pc [29] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [29] ), .QN(_14982_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_20 ( .D(\lsu.io_in_bits_pc [11] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [11] ), .QN(_14983_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_21 ( .D(\lsu.io_in_bits_pc [10] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [10] ), .QN(_14984_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_22 ( .D(\lsu.io_in_bits_pc [9] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [9] ), .QN(_14985_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_23 ( .D(\lsu.io_in_bits_pc [8] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [8] ), .QN(_14986_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_24 ( .D(\lsu.io_in_bits_pc [7] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [7] ), .QN(_14987_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_25 ( .D(\lsu.io_in_bits_pc [6] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [6] ), .QN(_14988_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_26 ( .D(\lsu.io_in_bits_pc [5] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [5] ), .QN(_14989_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_27 ( .D(\lsu.io_in_bits_pc [4] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [4] ), .QN(_14990_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_28 ( .D(\lsu.io_in_bits_pc [3] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [3] ), .QN(_14991_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_29 ( .D(\lsu.io_in_bits_pc [2] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [2] ), .QN(_14992_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_3 ( .D(\lsu.io_in_bits_pc [28] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [28] ), .QN(_14993_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_30 ( .D(\lsu.io_in_bits_pc [1] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [1] ), .QN(_14994_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_31 ( .D(\lsu.io_in_bits_pc [0] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [0] ), .QN(_14995_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_4 ( .D(\lsu.io_in_bits_pc [27] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [27] ), .QN(_14996_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_5 ( .D(\lsu.io_in_bits_pc [26] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [26] ), .QN(_14997_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_6 ( .D(\lsu.io_in_bits_pc [25] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [25] ), .QN(_14998_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_7 ( .D(\lsu.io_in_bits_pc [24] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [24] ), .QN(_14999_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_8 ( .D(\lsu.io_in_bits_pc [23] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [23] ), .QN(_15000_ ) );
DFF_X1 wbu_io_in_bits_r_pc_$_DFFE_PN__Q_9 ( .D(\lsu.io_in_bits_pc [22] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_pc [22] ), .QN(_15001_ ) );
DFF_X1 wbu_io_in_bits_r_rd_$_DFFE_PN__Q ( .D(\lsu.io_in_bits_rd [4] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd [4] ), .QN(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ) );
DFF_X1 wbu_io_in_bits_r_rd_$_DFFE_PN__Q_1 ( .D(\lsu.io_in_bits_rd [3] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd [3] ), .QN(_15002_ ) );
DFF_X1 wbu_io_in_bits_r_rd_$_DFFE_PN__Q_2 ( .D(\lsu.io_in_bits_rd [2] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd [2] ), .QN(_15003_ ) );
DFF_X1 wbu_io_in_bits_r_rd_$_DFFE_PN__Q_3 ( .D(\lsu.io_in_bits_rd [1] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd [1] ), .QN(_15004_ ) );
DFF_X1 wbu_io_in_bits_r_rd_$_DFFE_PN__Q_4 ( .D(\lsu.io_in_bits_rd [0] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd [0] ), .QN(_15005_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q ( .D(\lsu.io_out_bits_rd_wdata [31] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [31] ), .QN(_15006_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_1 ( .D(\lsu.io_out_bits_rd_wdata [30] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [30] ), .QN(_15007_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_10 ( .D(\lsu.io_out_bits_rd_wdata [21] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [21] ), .QN(_15008_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_11 ( .D(\lsu.io_out_bits_rd_wdata [20] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [20] ), .QN(_15009_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_12 ( .D(\lsu.io_out_bits_rd_wdata [19] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [19] ), .QN(_15010_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_13 ( .D(\lsu.io_out_bits_rd_wdata [18] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [18] ), .QN(_15011_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_14 ( .D(\lsu.io_out_bits_rd_wdata [17] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [17] ), .QN(_15012_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_15 ( .D(\lsu.io_out_bits_rd_wdata [16] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [16] ), .QN(_15013_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_16 ( .D(\lsu.io_out_bits_rd_wdata [15] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [15] ), .QN(_15014_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_17 ( .D(\lsu.io_out_bits_rd_wdata [14] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [14] ), .QN(_15015_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_18 ( .D(\lsu.io_out_bits_rd_wdata [13] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [13] ), .QN(_15016_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_19 ( .D(\lsu.io_out_bits_rd_wdata [12] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [12] ), .QN(_15017_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_2 ( .D(\lsu.io_out_bits_rd_wdata [29] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [29] ), .QN(_15018_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_20 ( .D(\lsu.io_out_bits_rd_wdata [11] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [11] ), .QN(_15019_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_21 ( .D(\lsu.io_out_bits_rd_wdata [10] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [10] ), .QN(_15020_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_22 ( .D(\lsu.io_out_bits_rd_wdata [9] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [9] ), .QN(_15021_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_23 ( .D(\lsu.io_out_bits_rd_wdata [8] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [8] ), .QN(_15022_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_24 ( .D(\lsu.io_out_bits_rd_wdata [7] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [7] ), .QN(_15023_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_25 ( .D(\lsu.io_out_bits_rd_wdata [6] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [6] ), .QN(_15024_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_26 ( .D(\lsu.io_out_bits_rd_wdata [5] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [5] ), .QN(_15025_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_27 ( .D(\lsu.io_out_bits_rd_wdata [4] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [4] ), .QN(_15026_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_28 ( .D(\lsu.io_out_bits_rd_wdata [3] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [3] ), .QN(_15027_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_29 ( .D(\lsu.io_out_bits_rd_wdata [2] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [2] ), .QN(_15028_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_3 ( .D(\lsu.io_out_bits_rd_wdata [28] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [28] ), .QN(_15029_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_30 ( .D(\lsu.io_out_bits_rd_wdata [1] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [1] ), .QN(_15030_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_31 ( .D(\lsu.io_out_bits_rd_wdata [0] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [0] ), .QN(_15031_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_4 ( .D(\lsu.io_out_bits_rd_wdata [27] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [27] ), .QN(_15032_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_5 ( .D(\lsu.io_out_bits_rd_wdata [26] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [26] ), .QN(_15033_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_6 ( .D(\lsu.io_out_bits_rd_wdata [25] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [25] ), .QN(_15034_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_7 ( .D(\lsu.io_out_bits_rd_wdata [24] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [24] ), .QN(_15035_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_8 ( .D(\lsu.io_out_bits_rd_wdata [23] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [23] ), .QN(_15036_ ) );
DFF_X1 wbu_io_in_bits_r_rd_wdata_$_DFFE_PN__Q_9 ( .D(\lsu.io_out_bits_rd_wdata [22] ), .CK(_13931_ ), .Q(\wbu.io_in_bits_rd_wdata [22] ), .QN(_15037_ ) );
DFF_X1 wbu_io_in_bits_r_wen_csr_$_DFFE_PN__Q ( .D(\lsu.io_in_bits_wen_csr ), .CK(_13931_ ), .Q(\wbu.io_in_bits_wen_csr ), .QN(_15038_ ) );
DFF_X1 wbu_io_in_bits_r_wen_rd_$_DFFE_PN__Q ( .D(\lsu.io_in_bits_wen_rd ), .CK(_13931_ ), .Q(\wbu.io_in_bits_wen_rd ), .QN(_13985_ ) );
DFF_X1 wbu_io_in_valid_REG_$_SDFF_PP0__Q ( .D(_00410_ ), .CK(clock ), .Q(\ifu.io_valid ), .QN(wbu_io_in_valid_REG_$_NOT__A_Y ) );
BUF_X8 fanout_buf_1 ( .A(\arbiter._io_axi_araddr_T ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(\arbiter._io_axi_araddr_T_6 ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(\arbiter._io_axi_araddr_T_6 ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(\exu.and_.io_is ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\exu.andi.io_is ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\exu.blt.io_is ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\exu.bltu.io_is ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\exu.ecall.io_is ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\exu.io_in_bits_jal ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\exu.io_in_bits_jalr ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\exu.io_in_bits_mret ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\exu.io_in_bits_sll ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\icache._io_out_arvalid_T ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\ifu.start [0] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\ifu.start [1] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(fanout_net_16 ), .Z(\io_master_awaddr [2] ) );
BUF_X8 fanout_buf_17 ( .A(fanout_net_27 ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(fanout_net_27 ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(fanout_net_27 ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(fanout_net_27 ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(fanout_net_27 ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(fanout_net_27 ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(reset ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(reset ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(reset ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(reset ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(reset ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\wbu.io_in_bits_csr_waddr [1] ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(fanout_net_36 ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(fanout_net_36 ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(fanout_net_36 ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(fanout_net_36 ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\wbu.io_in_bits_rd [4] ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\wbu.io_in_bits_rd [4] ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\wbu.io_in_bits_rd [4] ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\wbu.io_in_bits_rd [4] ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(wbu_io_in_bits_r_wen_rd_$_NAND__A_Y_$_NOR__B_A_$_ANDNOT__Y_A ), .Z(fanout_net_38 ) );

endmodule
