module state(
    
);
endmodule