//Generate the verilog at 2025-09-28T20:37:09 by iSTA.
module foo (
clock,
reset,
check_quest,
stall_quest_fencei,
check_assert,
stall_quest_exception_IFU,
readyFromIDU,
validToIDU,
arvalid,
arready,
rvalid,
rready,
rlast,
rmem_quest,
pc_jump,
mtvec,
pc,
inst,
araddr,
arid,
arlen,
arsize,
arburst,
rdata,
rresp,
rid
);

input clock ;
input reset ;
input check_quest ;
input stall_quest_fencei ;
output check_assert ;
input stall_quest_exception_IFU ;
input readyFromIDU ;
output validToIDU ;
output arvalid ;
input arready ;
input rvalid ;
output rready ;
input rlast ;
output rmem_quest ;
input [31:0] pc_jump ;
input [31:0] mtvec ;
output [31:0] pc ;
output [31:0] inst ;
output [31:0] araddr ;
output [3:0] arid ;
output [7:0] arlen ;
output [2:0] arsize ;
output [1:0] arburst ;
input [31:0] rdata ;
input [1:0] rresp ;
input [3:0] rid ;

wire clock ;
wire reset ;
wire check_quest ;
wire stall_quest_fencei ;
wire check_assert ;
wire stall_quest_exception_IFU ;
wire readyFromIDU ;
wire validToIDU ;
wire fanout_net_2 ;
wire fanout_net_6 ;
wire arvalid ;
wire arready ;
wire rvalid ;
wire rready ;
wire rlast ;
wire rmem_quest ;
wire _0000_ ;
wire _0001_ ;
wire _0002_ ;
wire _0003_ ;
wire _0004_ ;
wire _0005_ ;
wire _0006_ ;
wire _0007_ ;
wire _0008_ ;
wire _0009_ ;
wire _0010_ ;
wire _0011_ ;
wire _0012_ ;
wire _0013_ ;
wire _0014_ ;
wire _0015_ ;
wire _0016_ ;
wire _0017_ ;
wire _0018_ ;
wire _0019_ ;
wire _0020_ ;
wire _0021_ ;
wire _0022_ ;
wire _0023_ ;
wire _0024_ ;
wire _0025_ ;
wire _0026_ ;
wire _0027_ ;
wire _0028_ ;
wire _0029_ ;
wire _0030_ ;
wire _0031_ ;
wire _0032_ ;
wire _0033_ ;
wire _0034_ ;
wire _0035_ ;
wire _0036_ ;
wire _0037_ ;
wire _0038_ ;
wire _0039_ ;
wire _0040_ ;
wire _0041_ ;
wire _0042_ ;
wire _0043_ ;
wire _0044_ ;
wire _0045_ ;
wire _0046_ ;
wire _0047_ ;
wire _0048_ ;
wire _0049_ ;
wire _0050_ ;
wire _0051_ ;
wire _0052_ ;
wire _0053_ ;
wire _0054_ ;
wire _0055_ ;
wire _0056_ ;
wire _0057_ ;
wire _0058_ ;
wire _0059_ ;
wire _0060_ ;
wire _0061_ ;
wire _0062_ ;
wire _0063_ ;
wire _0064_ ;
wire _0065_ ;
wire _0066_ ;
wire _0067_ ;
wire _0068_ ;
wire _0069_ ;
wire _0070_ ;
wire _0071_ ;
wire _0072_ ;
wire _0073_ ;
wire _0074_ ;
wire _0075_ ;
wire _0076_ ;
wire _0077_ ;
wire _0078_ ;
wire _0079_ ;
wire _0080_ ;
wire _0081_ ;
wire _0082_ ;
wire _0083_ ;
wire _0084_ ;
wire _0085_ ;
wire _0086_ ;
wire _0087_ ;
wire _0088_ ;
wire _0089_ ;
wire _0090_ ;
wire _0091_ ;
wire _0092_ ;
wire _0093_ ;
wire _0094_ ;
wire _0095_ ;
wire _0096_ ;
wire _0097_ ;
wire _0098_ ;
wire _0099_ ;
wire _0100_ ;
wire _0101_ ;
wire _0102_ ;
wire _0103_ ;
wire _0104_ ;
wire _0105_ ;
wire _0106_ ;
wire _0107_ ;
wire _0108_ ;
wire _0109_ ;
wire _0110_ ;
wire _0111_ ;
wire _0112_ ;
wire _0113_ ;
wire _0114_ ;
wire _0115_ ;
wire _0116_ ;
wire _0117_ ;
wire _0118_ ;
wire _0119_ ;
wire _0120_ ;
wire _0121_ ;
wire _0122_ ;
wire _0123_ ;
wire _0124_ ;
wire _0125_ ;
wire _0126_ ;
wire _0127_ ;
wire _0128_ ;
wire _0129_ ;
wire _0130_ ;
wire _0131_ ;
wire _0132_ ;
wire _0133_ ;
wire _0134_ ;
wire _0135_ ;
wire _0136_ ;
wire _0137_ ;
wire _0138_ ;
wire _0139_ ;
wire _0140_ ;
wire _0141_ ;
wire _0142_ ;
wire _0143_ ;
wire _0144_ ;
wire _0145_ ;
wire _0146_ ;
wire _0147_ ;
wire _0148_ ;
wire _0149_ ;
wire _0150_ ;
wire _0151_ ;
wire _0152_ ;
wire _0153_ ;
wire _0154_ ;
wire _0155_ ;
wire _0156_ ;
wire _0157_ ;
wire _0158_ ;
wire _0159_ ;
wire _0160_ ;
wire _0161_ ;
wire _0162_ ;
wire _0163_ ;
wire _0164_ ;
wire _0165_ ;
wire _0166_ ;
wire _0167_ ;
wire _0168_ ;
wire _0169_ ;
wire _0170_ ;
wire _0171_ ;
wire _0172_ ;
wire _0173_ ;
wire _0174_ ;
wire _0175_ ;
wire _0176_ ;
wire _0177_ ;
wire _0178_ ;
wire _0179_ ;
wire _0180_ ;
wire _0181_ ;
wire _0182_ ;
wire _0183_ ;
wire _0184_ ;
wire _0185_ ;
wire _0186_ ;
wire _0187_ ;
wire _0188_ ;
wire _0189_ ;
wire _0190_ ;
wire _0191_ ;
wire _0192_ ;
wire _0193_ ;
wire _0194_ ;
wire _0195_ ;
wire _0196_ ;
wire _0197_ ;
wire _0198_ ;
wire _0199_ ;
wire _0200_ ;
wire _0201_ ;
wire _0202_ ;
wire _0203_ ;
wire _0204_ ;
wire _0205_ ;
wire _0206_ ;
wire _0207_ ;
wire _0208_ ;
wire _0209_ ;
wire _0210_ ;
wire _0211_ ;
wire _0212_ ;
wire _0213_ ;
wire _0214_ ;
wire _0215_ ;
wire _0216_ ;
wire _0217_ ;
wire _0218_ ;
wire _0219_ ;
wire _0220_ ;
wire _0221_ ;
wire _0222_ ;
wire _0223_ ;
wire _0224_ ;
wire _0225_ ;
wire _0226_ ;
wire _0227_ ;
wire _0228_ ;
wire _0229_ ;
wire _0230_ ;
wire _0231_ ;
wire _0232_ ;
wire _0233_ ;
wire _0234_ ;
wire _0235_ ;
wire _0236_ ;
wire _0237_ ;
wire _0238_ ;
wire _0239_ ;
wire _0240_ ;
wire _0241_ ;
wire _0242_ ;
wire _0243_ ;
wire _0244_ ;
wire _0245_ ;
wire _0246_ ;
wire _0247_ ;
wire _0248_ ;
wire _0249_ ;
wire _0250_ ;
wire _0251_ ;
wire _0252_ ;
wire _0253_ ;
wire _0254_ ;
wire _0255_ ;
wire _0256_ ;
wire _0257_ ;
wire _0258_ ;
wire _0259_ ;
wire _0260_ ;
wire _0261_ ;
wire _0262_ ;
wire _0263_ ;
wire _0264_ ;
wire _0265_ ;
wire _0266_ ;
wire _0267_ ;
wire _0268_ ;
wire _0269_ ;
wire _0270_ ;
wire _0271_ ;
wire _0272_ ;
wire _0273_ ;
wire _0274_ ;
wire _0275_ ;
wire _0276_ ;
wire _0277_ ;
wire _0278_ ;
wire _0279_ ;
wire _0280_ ;
wire _0281_ ;
wire _0282_ ;
wire _0283_ ;
wire _0284_ ;
wire _0285_ ;
wire _0286_ ;
wire _0287_ ;
wire _0288_ ;
wire _0289_ ;
wire _0290_ ;
wire _0291_ ;
wire _0292_ ;
wire _0293_ ;
wire _0294_ ;
wire _0295_ ;
wire _0296_ ;
wire _0297_ ;
wire _0298_ ;
wire _0299_ ;
wire _0300_ ;
wire _0301_ ;
wire _0302_ ;
wire _0303_ ;
wire _0304_ ;
wire _0305_ ;
wire _0306_ ;
wire _0307_ ;
wire _0308_ ;
wire _0309_ ;
wire _0310_ ;
wire _0311_ ;
wire _0312_ ;
wire _0313_ ;
wire _0314_ ;
wire _0315_ ;
wire _0316_ ;
wire _0317_ ;
wire _0318_ ;
wire _0319_ ;
wire _0320_ ;
wire _0321_ ;
wire _0322_ ;
wire _0323_ ;
wire _0324_ ;
wire _0325_ ;
wire _0326_ ;
wire _0327_ ;
wire _0328_ ;
wire _0329_ ;
wire _0330_ ;
wire _0331_ ;
wire _0332_ ;
wire _0333_ ;
wire _0334_ ;
wire _0335_ ;
wire _0336_ ;
wire _0337_ ;
wire _0338_ ;
wire _0339_ ;
wire _0340_ ;
wire _0341_ ;
wire _0342_ ;
wire _0343_ ;
wire _0344_ ;
wire _0345_ ;
wire _0346_ ;
wire _0347_ ;
wire _0348_ ;
wire _0349_ ;
wire _0350_ ;
wire _0351_ ;
wire _0352_ ;
wire _0353_ ;
wire _0354_ ;
wire _0355_ ;
wire _0356_ ;
wire _0357_ ;
wire _0358_ ;
wire _0359_ ;
wire _0360_ ;
wire _0361_ ;
wire _0362_ ;
wire _0363_ ;
wire _0364_ ;
wire _0365_ ;
wire _0366_ ;
wire _0367_ ;
wire _0368_ ;
wire _0369_ ;
wire _0370_ ;
wire _0371_ ;
wire _0372_ ;
wire _0373_ ;
wire _0374_ ;
wire _0375_ ;
wire _0376_ ;
wire _0377_ ;
wire _0378_ ;
wire _0379_ ;
wire _0380_ ;
wire _0381_ ;
wire _0382_ ;
wire _0383_ ;
wire _0384_ ;
wire _0385_ ;
wire _0386_ ;
wire _0387_ ;
wire _0388_ ;
wire _0389_ ;
wire _0390_ ;
wire _0391_ ;
wire _0392_ ;
wire _0393_ ;
wire _0394_ ;
wire _0395_ ;
wire _0396_ ;
wire _0397_ ;
wire _0398_ ;
wire _0399_ ;
wire _0400_ ;
wire _0401_ ;
wire _0402_ ;
wire _0403_ ;
wire _0404_ ;
wire _0405_ ;
wire _0406_ ;
wire _0407_ ;
wire _0408_ ;
wire _0409_ ;
wire _0410_ ;
wire _0411_ ;
wire _0412_ ;
wire _0413_ ;
wire _0414_ ;
wire _0415_ ;
wire _0416_ ;
wire _0417_ ;
wire _0418_ ;
wire _0419_ ;
wire _0420_ ;
wire _0421_ ;
wire _0422_ ;
wire _0423_ ;
wire _0424_ ;
wire _0425_ ;
wire _0426_ ;
wire _0427_ ;
wire _0428_ ;
wire _0429_ ;
wire _0430_ ;
wire _0431_ ;
wire _0432_ ;
wire _0433_ ;
wire _0434_ ;
wire _0435_ ;
wire _0436_ ;
wire _0437_ ;
wire _0438_ ;
wire _0439_ ;
wire _0440_ ;
wire _0441_ ;
wire _0442_ ;
wire _0443_ ;
wire _0444_ ;
wire _0445_ ;
wire _0446_ ;
wire _0447_ ;
wire _0448_ ;
wire _0449_ ;
wire _0450_ ;
wire _0451_ ;
wire _0452_ ;
wire _0453_ ;
wire _0454_ ;
wire _0455_ ;
wire _0456_ ;
wire _0457_ ;
wire _0458_ ;
wire _0459_ ;
wire _0460_ ;
wire _0461_ ;
wire _0462_ ;
wire _0463_ ;
wire _0464_ ;
wire _0465_ ;
wire _0466_ ;
wire _0467_ ;
wire _0468_ ;
wire _0469_ ;
wire _0470_ ;
wire _0471_ ;
wire _0472_ ;
wire _0473_ ;
wire _0474_ ;
wire _0475_ ;
wire _0476_ ;
wire _0477_ ;
wire _0478_ ;
wire _0479_ ;
wire _0480_ ;
wire _0481_ ;
wire _0482_ ;
wire _0483_ ;
wire _0484_ ;
wire _0485_ ;
wire _0486_ ;
wire _0487_ ;
wire _0488_ ;
wire _0489_ ;
wire _0490_ ;
wire _0491_ ;
wire _0492_ ;
wire _0493_ ;
wire _0494_ ;
wire _0495_ ;
wire _0496_ ;
wire _0497_ ;
wire _0498_ ;
wire _0499_ ;
wire _0500_ ;
wire _0501_ ;
wire _0502_ ;
wire _0503_ ;
wire _0504_ ;
wire _0505_ ;
wire _0506_ ;
wire _0507_ ;
wire _0508_ ;
wire _0509_ ;
wire _0510_ ;
wire _0511_ ;
wire _0512_ ;
wire _0513_ ;
wire _0514_ ;
wire _0515_ ;
wire _0516_ ;
wire _0517_ ;
wire _0518_ ;
wire _0519_ ;
wire _0520_ ;
wire _0521_ ;
wire _0522_ ;
wire _0523_ ;
wire _0524_ ;
wire _0525_ ;
wire _0526_ ;
wire _0527_ ;
wire _0528_ ;
wire _0529_ ;
wire _0530_ ;
wire _0531_ ;
wire _0532_ ;
wire _0533_ ;
wire _0534_ ;
wire _0535_ ;
wire _0536_ ;
wire _0537_ ;
wire _0538_ ;
wire _0539_ ;
wire _0540_ ;
wire _0541_ ;
wire _0542_ ;
wire _0543_ ;
wire _0544_ ;
wire _0545_ ;
wire _0546_ ;
wire _0547_ ;
wire _0548_ ;
wire _0549_ ;
wire _0550_ ;
wire _0551_ ;
wire _0552_ ;
wire _0553_ ;
wire _0554_ ;
wire _0555_ ;
wire _0556_ ;
wire _0557_ ;
wire _0558_ ;
wire _0559_ ;
wire _0560_ ;
wire _0561_ ;
wire _0562_ ;
wire _0563_ ;
wire _0564_ ;
wire _0565_ ;
wire _0566_ ;
wire _0567_ ;
wire _0568_ ;
wire _0569_ ;
wire _0570_ ;
wire _0571_ ;
wire _0572_ ;
wire _0573_ ;
wire _0574_ ;
wire _0575_ ;
wire _0576_ ;
wire _0577_ ;
wire _0578_ ;
wire _0579_ ;
wire _0580_ ;
wire _0581_ ;
wire _0582_ ;
wire _0583_ ;
wire _0584_ ;
wire _0585_ ;
wire _0586_ ;
wire _0587_ ;
wire _0588_ ;
wire _0589_ ;
wire _0590_ ;
wire _0591_ ;
wire _0592_ ;
wire _0593_ ;
wire _0594_ ;
wire _0595_ ;
wire _0596_ ;
wire _0597_ ;
wire _0598_ ;
wire _0599_ ;
wire _0600_ ;
wire _0601_ ;
wire _0602_ ;
wire _0603_ ;
wire _0604_ ;
wire _0605_ ;
wire _0606_ ;
wire _0607_ ;
wire _0608_ ;
wire _0609_ ;
wire _0610_ ;
wire _0611_ ;
wire _0612_ ;
wire _0613_ ;
wire _0614_ ;
wire _0615_ ;
wire _0616_ ;
wire _0617_ ;
wire _0618_ ;
wire _0619_ ;
wire _0620_ ;
wire _0621_ ;
wire _0622_ ;
wire _0623_ ;
wire _0624_ ;
wire _0625_ ;
wire _0626_ ;
wire _0627_ ;
wire _0628_ ;
wire _0629_ ;
wire _0630_ ;
wire _0631_ ;
wire _0632_ ;
wire _0633_ ;
wire _0634_ ;
wire _0635_ ;
wire _0636_ ;
wire _0637_ ;
wire _0638_ ;
wire _0639_ ;
wire _0640_ ;
wire _0641_ ;
wire _0642_ ;
wire _0643_ ;
wire _0644_ ;
wire _0645_ ;
wire _0646_ ;
wire _0647_ ;
wire _0648_ ;
wire _0649_ ;
wire _0650_ ;
wire _0651_ ;
wire _0652_ ;
wire _0653_ ;
wire _0654_ ;
wire _0655_ ;
wire _0656_ ;
wire _0657_ ;
wire _0658_ ;
wire _0659_ ;
wire _0660_ ;
wire _0661_ ;
wire _0662_ ;
wire _0663_ ;
wire _0664_ ;
wire _0665_ ;
wire _0666_ ;
wire _0667_ ;
wire _0668_ ;
wire _0669_ ;
wire _0670_ ;
wire _0671_ ;
wire _0672_ ;
wire _0673_ ;
wire _0674_ ;
wire _0675_ ;
wire _0676_ ;
wire _0677_ ;
wire _0678_ ;
wire _0679_ ;
wire _0680_ ;
wire _0681_ ;
wire _0682_ ;
wire _0683_ ;
wire _0684_ ;
wire _0685_ ;
wire _0686_ ;
wire _0687_ ;
wire _0688_ ;
wire _0689_ ;
wire _0690_ ;
wire _0691_ ;
wire _0692_ ;
wire _0693_ ;
wire _0694_ ;
wire _0695_ ;
wire _0696_ ;
wire _0697_ ;
wire _0698_ ;
wire _0699_ ;
wire _0700_ ;
wire _0701_ ;
wire _0702_ ;
wire _0703_ ;
wire _0704_ ;
wire _0705_ ;
wire _0706_ ;
wire _0707_ ;
wire _0708_ ;
wire _0709_ ;
wire _0710_ ;
wire _0711_ ;
wire _0712_ ;
wire _0713_ ;
wire _0714_ ;
wire _0715_ ;
wire _0716_ ;
wire _0717_ ;
wire _0718_ ;
wire _0719_ ;
wire _0720_ ;
wire _0721_ ;
wire _0722_ ;
wire _0723_ ;
wire _0724_ ;
wire _0725_ ;
wire _0726_ ;
wire _0727_ ;
wire _0728_ ;
wire _0729_ ;
wire _0730_ ;
wire _0731_ ;
wire _0732_ ;
wire _0733_ ;
wire _0734_ ;
wire _0735_ ;
wire _0736_ ;
wire _0737_ ;
wire _0738_ ;
wire _0739_ ;
wire _0740_ ;
wire _0741_ ;
wire _0742_ ;
wire _0743_ ;
wire _0744_ ;
wire _0745_ ;
wire _0746_ ;
wire _0747_ ;
wire _0748_ ;
wire _0749_ ;
wire _0750_ ;
wire _0751_ ;
wire _0752_ ;
wire _0753_ ;
wire _0754_ ;
wire _0755_ ;
wire _0756_ ;
wire _0757_ ;
wire _0758_ ;
wire _0759_ ;
wire _0760_ ;
wire _0761_ ;
wire _0762_ ;
wire _0763_ ;
wire _0764_ ;
wire _0765_ ;
wire _0766_ ;
wire _0767_ ;
wire _0768_ ;
wire _0769_ ;
wire _0770_ ;
wire _0771_ ;
wire _0772_ ;
wire _0773_ ;
wire _0774_ ;
wire _0775_ ;
wire _0776_ ;
wire _0777_ ;
wire _0778_ ;
wire _0779_ ;
wire _0780_ ;
wire _0781_ ;
wire _0782_ ;
wire _0783_ ;
wire _0784_ ;
wire _0785_ ;
wire _0786_ ;
wire _0787_ ;
wire _0788_ ;
wire _0789_ ;
wire _0790_ ;
wire _0791_ ;
wire _0792_ ;
wire _0793_ ;
wire _0794_ ;
wire _0795_ ;
wire _0796_ ;
wire _0797_ ;
wire _0798_ ;
wire _0799_ ;
wire _0800_ ;
wire _0801_ ;
wire _0802_ ;
wire _0803_ ;
wire _0804_ ;
wire _0805_ ;
wire _0806_ ;
wire _0807_ ;
wire _0808_ ;
wire _0809_ ;
wire _0810_ ;
wire _0811_ ;
wire _0812_ ;
wire _0813_ ;
wire _0814_ ;
wire _0815_ ;
wire _0816_ ;
wire _0817_ ;
wire _0818_ ;
wire _0819_ ;
wire _0820_ ;
wire _0821_ ;
wire _0822_ ;
wire _0823_ ;
wire _0824_ ;
wire _0825_ ;
wire _0826_ ;
wire _0827_ ;
wire _0828_ ;
wire _0829_ ;
wire _0830_ ;
wire _0831_ ;
wire _0832_ ;
wire _0833_ ;
wire _0834_ ;
wire _0835_ ;
wire _0836_ ;
wire _0837_ ;
wire _0838_ ;
wire _0839_ ;
wire _0840_ ;
wire _0841_ ;
wire _0842_ ;
wire _0843_ ;
wire _0844_ ;
wire _0845_ ;
wire _0846_ ;
wire _0847_ ;
wire _0848_ ;
wire _0849_ ;
wire _0850_ ;
wire _0851_ ;
wire _0852_ ;
wire _0853_ ;
wire _0854_ ;
wire _0855_ ;
wire _0856_ ;
wire _0857_ ;
wire _0858_ ;
wire _0859_ ;
wire _0860_ ;
wire _0861_ ;
wire _0862_ ;
wire _0863_ ;
wire _0864_ ;
wire _0865_ ;
wire _0866_ ;
wire _0867_ ;
wire _0868_ ;
wire _0869_ ;
wire _0870_ ;
wire _0871_ ;
wire _0872_ ;
wire _0873_ ;
wire _0874_ ;
wire _0875_ ;
wire _0876_ ;
wire _0877_ ;
wire _0878_ ;
wire _0879_ ;
wire _0880_ ;
wire _0881_ ;
wire _0882_ ;
wire _0883_ ;
wire _0884_ ;
wire _0885_ ;
wire _0886_ ;
wire _0887_ ;
wire _0888_ ;
wire _0889_ ;
wire _0890_ ;
wire _0891_ ;
wire _0892_ ;
wire _0893_ ;
wire _0894_ ;
wire _0895_ ;
wire _0896_ ;
wire _0897_ ;
wire _0898_ ;
wire _0899_ ;
wire _0900_ ;
wire _0901_ ;
wire _0902_ ;
wire _0903_ ;
wire _0904_ ;
wire _0905_ ;
wire _0906_ ;
wire _0907_ ;
wire _0908_ ;
wire _0909_ ;
wire _0910_ ;
wire _0911_ ;
wire _0912_ ;
wire _0913_ ;
wire _0914_ ;
wire _0915_ ;
wire _0916_ ;
wire _0917_ ;
wire _0918_ ;
wire _0919_ ;
wire _0920_ ;
wire _0921_ ;
wire _0922_ ;
wire _0923_ ;
wire _0924_ ;
wire _0925_ ;
wire _0926_ ;
wire _0927_ ;
wire _0928_ ;
wire _0929_ ;
wire _0930_ ;
wire _0931_ ;
wire _0932_ ;
wire _0933_ ;
wire _0934_ ;
wire _0935_ ;
wire _0936_ ;
wire _0937_ ;
wire _0938_ ;
wire _0939_ ;
wire _0940_ ;
wire _0941_ ;
wire _0942_ ;
wire _0943_ ;
wire _0944_ ;
wire _0945_ ;
wire _0946_ ;
wire _0947_ ;
wire _0948_ ;
wire _0949_ ;
wire _0950_ ;
wire _0951_ ;
wire _0952_ ;
wire _0953_ ;
wire _0954_ ;
wire _0955_ ;
wire _0956_ ;
wire _0957_ ;
wire _0958_ ;
wire _0959_ ;
wire _0960_ ;
wire _0961_ ;
wire _0962_ ;
wire _0963_ ;
wire _0964_ ;
wire _0965_ ;
wire _0966_ ;
wire _0967_ ;
wire _0968_ ;
wire _0969_ ;
wire _0970_ ;
wire _0971_ ;
wire _0972_ ;
wire _0973_ ;
wire _0974_ ;
wire _0975_ ;
wire _0976_ ;
wire _0977_ ;
wire _0978_ ;
wire _0979_ ;
wire _0980_ ;
wire _0981_ ;
wire _0982_ ;
wire _0983_ ;
wire _0984_ ;
wire _0985_ ;
wire _0986_ ;
wire _0987_ ;
wire _0988_ ;
wire _0989_ ;
wire _0990_ ;
wire _0991_ ;
wire _0992_ ;
wire _0993_ ;
wire _0994_ ;
wire _0995_ ;
wire _0996_ ;
wire _0997_ ;
wire _0998_ ;
wire _0999_ ;
wire _1000_ ;
wire _1001_ ;
wire _1002_ ;
wire _1003_ ;
wire _1004_ ;
wire _1005_ ;
wire _1006_ ;
wire _1007_ ;
wire _1008_ ;
wire _1009_ ;
wire _1010_ ;
wire _1011_ ;
wire _1012_ ;
wire _1013_ ;
wire _1014_ ;
wire _1015_ ;
wire _1016_ ;
wire _1017_ ;
wire _1018_ ;
wire _1019_ ;
wire _1020_ ;
wire _1021_ ;
wire _1022_ ;
wire _1023_ ;
wire _1024_ ;
wire _1025_ ;
wire _1026_ ;
wire _1027_ ;
wire _1028_ ;
wire _1029_ ;
wire _1030_ ;
wire _1031_ ;
wire _1032_ ;
wire _1033_ ;
wire _1034_ ;
wire _1035_ ;
wire _1036_ ;
wire _1037_ ;
wire _1038_ ;
wire _1039_ ;
wire _1040_ ;
wire _1041_ ;
wire _1042_ ;
wire _1043_ ;
wire _1044_ ;
wire _1045_ ;
wire _1046_ ;
wire _1047_ ;
wire _1048_ ;
wire _1049_ ;
wire _1050_ ;
wire _1051_ ;
wire _1052_ ;
wire _1053_ ;
wire _1054_ ;
wire _1055_ ;
wire _1056_ ;
wire _1057_ ;
wire _1058_ ;
wire _1059_ ;
wire _1060_ ;
wire _1061_ ;
wire _1062_ ;
wire _1063_ ;
wire _1064_ ;
wire _1065_ ;
wire _1066_ ;
wire _1067_ ;
wire _1068_ ;
wire _1069_ ;
wire _1070_ ;
wire _1071_ ;
wire _1072_ ;
wire _1073_ ;
wire _1074_ ;
wire _1075_ ;
wire _1076_ ;
wire _1077_ ;
wire _1078_ ;
wire _1079_ ;
wire _1080_ ;
wire _1081_ ;
wire _1082_ ;
wire _1083_ ;
wire _1084_ ;
wire _1085_ ;
wire _1086_ ;
wire _1087_ ;
wire _1088_ ;
wire _1089_ ;
wire _1090_ ;
wire _1091_ ;
wire _1092_ ;
wire _1093_ ;
wire _1094_ ;
wire _1095_ ;
wire _1096_ ;
wire _1097_ ;
wire _1098_ ;
wire _1099_ ;
wire _1100_ ;
wire _1101_ ;
wire _1102_ ;
wire _1103_ ;
wire _1104_ ;
wire _1105_ ;
wire _1106_ ;
wire _1107_ ;
wire _1108_ ;
wire _1109_ ;
wire _1110_ ;
wire _1111_ ;
wire _1112_ ;
wire _1113_ ;
wire _1114_ ;
wire _1115_ ;
wire _1116_ ;
wire _1117_ ;
wire _1118_ ;
wire _1119_ ;
wire _1120_ ;
wire _1121_ ;
wire _1122_ ;
wire _1123_ ;
wire _1124_ ;
wire _1125_ ;
wire _1126_ ;
wire _1127_ ;
wire _1128_ ;
wire _1129_ ;
wire _1130_ ;
wire _1131_ ;
wire _1132_ ;
wire _1133_ ;
wire _1134_ ;
wire _1135_ ;
wire _1136_ ;
wire _1137_ ;
wire _1138_ ;
wire _1139_ ;
wire _1140_ ;
wire _1141_ ;
wire _1142_ ;
wire _1143_ ;
wire _1144_ ;
wire _1145_ ;
wire _1146_ ;
wire _1147_ ;
wire _1148_ ;
wire _1149_ ;
wire _1150_ ;
wire _1151_ ;
wire _1152_ ;
wire _1153_ ;
wire _1154_ ;
wire _1155_ ;
wire _1156_ ;
wire _1157_ ;
wire _1158_ ;
wire _1159_ ;
wire _1160_ ;
wire _1161_ ;
wire _1162_ ;
wire _1163_ ;
wire _1164_ ;
wire _1165_ ;
wire _1166_ ;
wire _1167_ ;
wire _1168_ ;
wire _1169_ ;
wire _1170_ ;
wire _1171_ ;
wire _1172_ ;
wire _1173_ ;
wire _1174_ ;
wire _1175_ ;
wire _1176_ ;
wire _1177_ ;
wire _1178_ ;
wire _1179_ ;
wire _1180_ ;
wire _1181_ ;
wire _1182_ ;
wire _1183_ ;
wire _1184_ ;
wire _1185_ ;
wire _1186_ ;
wire _1187_ ;
wire _1188_ ;
wire _1189_ ;
wire _1190_ ;
wire _1191_ ;
wire _1192_ ;
wire _1193_ ;
wire _1194_ ;
wire _1195_ ;
wire _1196_ ;
wire _1197_ ;
wire _1198_ ;
wire _1199_ ;
wire _1200_ ;
wire _1201_ ;
wire _1202_ ;
wire _1203_ ;
wire _1204_ ;
wire _1205_ ;
wire _1206_ ;
wire _1207_ ;
wire _1208_ ;
wire _1209_ ;
wire _1210_ ;
wire _1211_ ;
wire _1212_ ;
wire _1213_ ;
wire _1214_ ;
wire _1215_ ;
wire _1216_ ;
wire _1217_ ;
wire _1218_ ;
wire _1219_ ;
wire _1220_ ;
wire _1221_ ;
wire _1222_ ;
wire _1223_ ;
wire _1224_ ;
wire _1225_ ;
wire _1226_ ;
wire _1227_ ;
wire _1228_ ;
wire _1229_ ;
wire _1230_ ;
wire _1231_ ;
wire _1232_ ;
wire _1233_ ;
wire _1234_ ;
wire _1235_ ;
wire _1236_ ;
wire _1237_ ;
wire _1238_ ;
wire _1239_ ;
wire _1240_ ;
wire _1241_ ;
wire _1242_ ;
wire _1243_ ;
wire _1244_ ;
wire _1245_ ;
wire _1246_ ;
wire _1247_ ;
wire _1248_ ;
wire _1249_ ;
wire _1250_ ;
wire _1251_ ;
wire _1252_ ;
wire _1253_ ;
wire _1254_ ;
wire _1255_ ;
wire _1256_ ;
wire _1257_ ;
wire _1258_ ;
wire _1259_ ;
wire _1260_ ;
wire _1261_ ;
wire _1262_ ;
wire _1263_ ;
wire _1264_ ;
wire _1265_ ;
wire _1266_ ;
wire _1267_ ;
wire _1268_ ;
wire _1269_ ;
wire _1270_ ;
wire _1271_ ;
wire _1272_ ;
wire _1273_ ;
wire _1274_ ;
wire _1275_ ;
wire _1276_ ;
wire _1277_ ;
wire _1278_ ;
wire _1279_ ;
wire _1280_ ;
wire _1281_ ;
wire _1282_ ;
wire _1283_ ;
wire _1284_ ;
wire _1285_ ;
wire _1286_ ;
wire _1287_ ;
wire _1288_ ;
wire _1289_ ;
wire _1290_ ;
wire _1291_ ;
wire _1292_ ;
wire _1293_ ;
wire _1294_ ;
wire _1295_ ;
wire _1296_ ;
wire _1297_ ;
wire _1298_ ;
wire _1299_ ;
wire _1300_ ;
wire _1301_ ;
wire _1302_ ;
wire _1303_ ;
wire _1304_ ;
wire _1305_ ;
wire _1306_ ;
wire _1307_ ;
wire _1308_ ;
wire _1309_ ;
wire _1310_ ;
wire _1311_ ;
wire _1312_ ;
wire _1313_ ;
wire _1314_ ;
wire _1315_ ;
wire _1316_ ;
wire _1317_ ;
wire _1318_ ;
wire _1319_ ;
wire _1320_ ;
wire _1321_ ;
wire _1322_ ;
wire _1323_ ;
wire _1324_ ;
wire _1325_ ;
wire _1326_ ;
wire _1327_ ;
wire _1328_ ;
wire _1329_ ;
wire _1330_ ;
wire _1331_ ;
wire _1332_ ;
wire _1333_ ;
wire _1334_ ;
wire _1335_ ;
wire _1336_ ;
wire _1337_ ;
wire _1338_ ;
wire _1339_ ;
wire _1340_ ;
wire _1341_ ;
wire _1342_ ;
wire _1343_ ;
wire _1344_ ;
wire _1345_ ;
wire _1346_ ;
wire _1347_ ;
wire _1348_ ;
wire _1349_ ;
wire _1350_ ;
wire _1351_ ;
wire _1352_ ;
wire _1353_ ;
wire _1354_ ;
wire _1355_ ;
wire _1356_ ;
wire _1357_ ;
wire _1358_ ;
wire _1359_ ;
wire _1360_ ;
wire _1361_ ;
wire _1362_ ;
wire _1363_ ;
wire _1364_ ;
wire _1365_ ;
wire _1366_ ;
wire _1367_ ;
wire _1368_ ;
wire _1369_ ;
wire _1370_ ;
wire _1371_ ;
wire _1372_ ;
wire _1373_ ;
wire _1374_ ;
wire _1375_ ;
wire _1376_ ;
wire _1377_ ;
wire _1378_ ;
wire _1379_ ;
wire _1380_ ;
wire _1381_ ;
wire _1382_ ;
wire _1383_ ;
wire _1384_ ;
wire _1385_ ;
wire _1386_ ;
wire _1387_ ;
wire _1388_ ;
wire _1389_ ;
wire _1390_ ;
wire _1391_ ;
wire _1392_ ;
wire _1393_ ;
wire _1394_ ;
wire _1395_ ;
wire _1396_ ;
wire _1397_ ;
wire _1398_ ;
wire _1399_ ;
wire _1400_ ;
wire _1401_ ;
wire _1402_ ;
wire _1403_ ;
wire _1404_ ;
wire _1405_ ;
wire _1406_ ;
wire _1407_ ;
wire _1408_ ;
wire _1409_ ;
wire _1410_ ;
wire _1411_ ;
wire _1412_ ;
wire _1413_ ;
wire _1414_ ;
wire _1415_ ;
wire _1416_ ;
wire _1417_ ;
wire _1418_ ;
wire _1419_ ;
wire _1420_ ;
wire _1421_ ;
wire _1422_ ;
wire _1423_ ;
wire _1424_ ;
wire _1425_ ;
wire _1426_ ;
wire _1427_ ;
wire _1428_ ;
wire _1429_ ;
wire _1430_ ;
wire _1431_ ;
wire _1432_ ;
wire _1433_ ;
wire _1434_ ;
wire _1435_ ;
wire _1436_ ;
wire _1437_ ;
wire _1438_ ;
wire _1439_ ;
wire _1440_ ;
wire _1441_ ;
wire _1442_ ;
wire _1443_ ;
wire _1444_ ;
wire _1445_ ;
wire _1446_ ;
wire _1447_ ;
wire _1448_ ;
wire _1449_ ;
wire _1450_ ;
wire _1451_ ;
wire _1452_ ;
wire _1453_ ;
wire _1454_ ;
wire _1455_ ;
wire _1456_ ;
wire _1457_ ;
wire _1458_ ;
wire _1459_ ;
wire _1460_ ;
wire _1461_ ;
wire _1462_ ;
wire _1463_ ;
wire _1464_ ;
wire _1465_ ;
wire _1466_ ;
wire _1467_ ;
wire _1468_ ;
wire _1469_ ;
wire _1470_ ;
wire _1471_ ;
wire _1472_ ;
wire _1473_ ;
wire _1474_ ;
wire _1475_ ;
wire _1476_ ;
wire _1477_ ;
wire _1478_ ;
wire _1479_ ;
wire _1480_ ;
wire _1481_ ;
wire _1482_ ;
wire _1483_ ;
wire _1484_ ;
wire _1485_ ;
wire _1486_ ;
wire _1487_ ;
wire _1488_ ;
wire _1489_ ;
wire _1490_ ;
wire _1491_ ;
wire _1492_ ;
wire _1493_ ;
wire _1494_ ;
wire _1495_ ;
wire _1496_ ;
wire _1497_ ;
wire _1498_ ;
wire _1499_ ;
wire _1500_ ;
wire _1501_ ;
wire _1502_ ;
wire _1503_ ;
wire _1504_ ;
wire _1505_ ;
wire _1506_ ;
wire _1507_ ;
wire _1508_ ;
wire _1509_ ;
wire _1510_ ;
wire _1511_ ;
wire _1512_ ;
wire _1513_ ;
wire _1514_ ;
wire _1515_ ;
wire _1516_ ;
wire _1517_ ;
wire _1518_ ;
wire _1519_ ;
wire _1520_ ;
wire _1521_ ;
wire _1522_ ;
wire _1523_ ;
wire _1524_ ;
wire _1525_ ;
wire _1526_ ;
wire _1527_ ;
wire _1528_ ;
wire _1529_ ;
wire _1530_ ;
wire _1531_ ;
wire _1532_ ;
wire _1533_ ;
wire _1534_ ;
wire _1535_ ;
wire _1536_ ;
wire _1537_ ;
wire _1538_ ;
wire _1539_ ;
wire _1540_ ;
wire _1541_ ;
wire _1542_ ;
wire _1543_ ;
wire _1544_ ;
wire _1545_ ;
wire _1546_ ;
wire _1547_ ;
wire _1548_ ;
wire _1549_ ;
wire _1550_ ;
wire _1551_ ;
wire _1552_ ;
wire _1553_ ;
wire _1554_ ;
wire _1555_ ;
wire _1556_ ;
wire _1557_ ;
wire _1558_ ;
wire _1559_ ;
wire _1560_ ;
wire _1561_ ;
wire _1562_ ;
wire _1563_ ;
wire _1564_ ;
wire _1565_ ;
wire _1566_ ;
wire _1567_ ;
wire _1568_ ;
wire _1569_ ;
wire _1570_ ;
wire _1571_ ;
wire _1572_ ;
wire _1573_ ;
wire _1574_ ;
wire _1575_ ;
wire _1576_ ;
wire _1577_ ;
wire _1578_ ;
wire _1579_ ;
wire _1580_ ;
wire _1581_ ;
wire _1582_ ;
wire _1583_ ;
wire _1584_ ;
wire _1585_ ;
wire _1586_ ;
wire _1587_ ;
wire _1588_ ;
wire _1589_ ;
wire _1590_ ;
wire _1591_ ;
wire _1592_ ;
wire _1593_ ;
wire _1594_ ;
wire _1595_ ;
wire _1596_ ;
wire _1597_ ;
wire _1598_ ;
wire _1599_ ;
wire _1600_ ;
wire _1601_ ;
wire _1602_ ;
wire _1603_ ;
wire _1604_ ;
wire _1605_ ;
wire _1606_ ;
wire _1607_ ;
wire _1608_ ;
wire _1609_ ;
wire _1610_ ;
wire _1611_ ;
wire _1612_ ;
wire _1613_ ;
wire _1614_ ;
wire _1615_ ;
wire _1616_ ;
wire _1617_ ;
wire _1618_ ;
wire _1619_ ;
wire _1620_ ;
wire _1621_ ;
wire _1622_ ;
wire _1623_ ;
wire _1624_ ;
wire _1625_ ;
wire _1626_ ;
wire _1627_ ;
wire _1628_ ;
wire _1629_ ;
wire _1630_ ;
wire _1631_ ;
wire check_assert_$_DFFE_PP__Q_E ;
wire check_assert_$_DFFE_PP__Q_E_$_ANDNOT__Y_B_$_MUX__Y_A ;
wire \myicache.data[0][0] ;
wire \myicache.data[0][10] ;
wire \myicache.data[0][11] ;
wire \myicache.data[0][12] ;
wire \myicache.data[0][13] ;
wire \myicache.data[0][14] ;
wire \myicache.data[0][15] ;
wire \myicache.data[0][16] ;
wire \myicache.data[0][17] ;
wire \myicache.data[0][18] ;
wire \myicache.data[0][19] ;
wire \myicache.data[0][1] ;
wire \myicache.data[0][20] ;
wire \myicache.data[0][21] ;
wire \myicache.data[0][22] ;
wire \myicache.data[0][23] ;
wire \myicache.data[0][24] ;
wire \myicache.data[0][25] ;
wire \myicache.data[0][26] ;
wire \myicache.data[0][27] ;
wire \myicache.data[0][28] ;
wire \myicache.data[0][29] ;
wire \myicache.data[0][2] ;
wire \myicache.data[0][30] ;
wire \myicache.data[0][31] ;
wire \myicache.data[0][3] ;
wire \myicache.data[0][4] ;
wire \myicache.data[0][5] ;
wire \myicache.data[0][6] ;
wire \myicache.data[0][7] ;
wire \myicache.data[0][8] ;
wire \myicache.data[0][9] ;
wire \myicache.data[1][0] ;
wire \myicache.data[1][10] ;
wire \myicache.data[1][11] ;
wire \myicache.data[1][12] ;
wire \myicache.data[1][13] ;
wire \myicache.data[1][14] ;
wire \myicache.data[1][15] ;
wire \myicache.data[1][16] ;
wire \myicache.data[1][17] ;
wire \myicache.data[1][18] ;
wire \myicache.data[1][19] ;
wire \myicache.data[1][1] ;
wire \myicache.data[1][20] ;
wire \myicache.data[1][21] ;
wire \myicache.data[1][22] ;
wire \myicache.data[1][23] ;
wire \myicache.data[1][24] ;
wire \myicache.data[1][25] ;
wire \myicache.data[1][26] ;
wire \myicache.data[1][27] ;
wire \myicache.data[1][28] ;
wire \myicache.data[1][29] ;
wire \myicache.data[1][2] ;
wire \myicache.data[1][30] ;
wire \myicache.data[1][31] ;
wire \myicache.data[1][3] ;
wire \myicache.data[1][4] ;
wire \myicache.data[1][5] ;
wire \myicache.data[1][6] ;
wire \myicache.data[1][7] ;
wire \myicache.data[1][8] ;
wire \myicache.data[1][9] ;
wire \myicache.data[2][0] ;
wire \myicache.data[2][10] ;
wire \myicache.data[2][11] ;
wire \myicache.data[2][12] ;
wire \myicache.data[2][13] ;
wire \myicache.data[2][14] ;
wire \myicache.data[2][15] ;
wire \myicache.data[2][16] ;
wire \myicache.data[2][17] ;
wire \myicache.data[2][18] ;
wire \myicache.data[2][19] ;
wire \myicache.data[2][1] ;
wire \myicache.data[2][20] ;
wire \myicache.data[2][21] ;
wire \myicache.data[2][22] ;
wire \myicache.data[2][23] ;
wire \myicache.data[2][24] ;
wire \myicache.data[2][25] ;
wire \myicache.data[2][26] ;
wire \myicache.data[2][27] ;
wire \myicache.data[2][28] ;
wire \myicache.data[2][29] ;
wire \myicache.data[2][2] ;
wire \myicache.data[2][30] ;
wire \myicache.data[2][31] ;
wire \myicache.data[2][3] ;
wire \myicache.data[2][4] ;
wire \myicache.data[2][5] ;
wire \myicache.data[2][6] ;
wire \myicache.data[2][7] ;
wire \myicache.data[2][8] ;
wire \myicache.data[2][9] ;
wire \myicache.data[3][0] ;
wire \myicache.data[3][10] ;
wire \myicache.data[3][11] ;
wire \myicache.data[3][12] ;
wire \myicache.data[3][13] ;
wire \myicache.data[3][14] ;
wire \myicache.data[3][15] ;
wire \myicache.data[3][16] ;
wire \myicache.data[3][17] ;
wire \myicache.data[3][18] ;
wire \myicache.data[3][19] ;
wire \myicache.data[3][1] ;
wire \myicache.data[3][20] ;
wire \myicache.data[3][21] ;
wire \myicache.data[3][22] ;
wire \myicache.data[3][23] ;
wire \myicache.data[3][24] ;
wire \myicache.data[3][25] ;
wire \myicache.data[3][26] ;
wire \myicache.data[3][27] ;
wire \myicache.data[3][28] ;
wire \myicache.data[3][29] ;
wire \myicache.data[3][2] ;
wire \myicache.data[3][30] ;
wire \myicache.data[3][31] ;
wire \myicache.data[3][3] ;
wire \myicache.data[3][4] ;
wire \myicache.data[3][5] ;
wire \myicache.data[3][6] ;
wire \myicache.data[3][7] ;
wire \myicache.data[3][8] ;
wire \myicache.data[3][9] ;
wire \myicache.data[4][0] ;
wire \myicache.data[4][10] ;
wire \myicache.data[4][11] ;
wire \myicache.data[4][12] ;
wire \myicache.data[4][13] ;
wire \myicache.data[4][14] ;
wire \myicache.data[4][15] ;
wire \myicache.data[4][16] ;
wire \myicache.data[4][17] ;
wire \myicache.data[4][18] ;
wire \myicache.data[4][19] ;
wire \myicache.data[4][1] ;
wire \myicache.data[4][20] ;
wire \myicache.data[4][21] ;
wire \myicache.data[4][22] ;
wire \myicache.data[4][23] ;
wire \myicache.data[4][24] ;
wire \myicache.data[4][25] ;
wire \myicache.data[4][26] ;
wire \myicache.data[4][27] ;
wire \myicache.data[4][28] ;
wire \myicache.data[4][29] ;
wire \myicache.data[4][2] ;
wire \myicache.data[4][30] ;
wire \myicache.data[4][31] ;
wire \myicache.data[4][3] ;
wire \myicache.data[4][4] ;
wire \myicache.data[4][5] ;
wire \myicache.data[4][6] ;
wire \myicache.data[4][7] ;
wire \myicache.data[4][8] ;
wire \myicache.data[4][9] ;
wire \myicache.data[5][0] ;
wire \myicache.data[5][10] ;
wire \myicache.data[5][11] ;
wire \myicache.data[5][12] ;
wire \myicache.data[5][13] ;
wire \myicache.data[5][14] ;
wire \myicache.data[5][15] ;
wire \myicache.data[5][16] ;
wire \myicache.data[5][17] ;
wire \myicache.data[5][18] ;
wire \myicache.data[5][19] ;
wire \myicache.data[5][1] ;
wire \myicache.data[5][20] ;
wire \myicache.data[5][21] ;
wire \myicache.data[5][22] ;
wire \myicache.data[5][23] ;
wire \myicache.data[5][24] ;
wire \myicache.data[5][25] ;
wire \myicache.data[5][26] ;
wire \myicache.data[5][27] ;
wire \myicache.data[5][28] ;
wire \myicache.data[5][29] ;
wire \myicache.data[5][2] ;
wire \myicache.data[5][30] ;
wire \myicache.data[5][31] ;
wire \myicache.data[5][3] ;
wire \myicache.data[5][4] ;
wire \myicache.data[5][5] ;
wire \myicache.data[5][6] ;
wire \myicache.data[5][7] ;
wire \myicache.data[5][8] ;
wire \myicache.data[5][9] ;
wire \myicache.data[6][0] ;
wire \myicache.data[6][10] ;
wire \myicache.data[6][11] ;
wire \myicache.data[6][12] ;
wire \myicache.data[6][13] ;
wire \myicache.data[6][14] ;
wire \myicache.data[6][15] ;
wire \myicache.data[6][16] ;
wire \myicache.data[6][17] ;
wire \myicache.data[6][18] ;
wire \myicache.data[6][19] ;
wire \myicache.data[6][1] ;
wire \myicache.data[6][20] ;
wire \myicache.data[6][21] ;
wire \myicache.data[6][22] ;
wire \myicache.data[6][23] ;
wire \myicache.data[6][24] ;
wire \myicache.data[6][25] ;
wire \myicache.data[6][26] ;
wire \myicache.data[6][27] ;
wire \myicache.data[6][28] ;
wire \myicache.data[6][29] ;
wire \myicache.data[6][2] ;
wire \myicache.data[6][30] ;
wire \myicache.data[6][31] ;
wire \myicache.data[6][3] ;
wire \myicache.data[6][4] ;
wire \myicache.data[6][5] ;
wire \myicache.data[6][6] ;
wire \myicache.data[6][7] ;
wire \myicache.data[6][8] ;
wire \myicache.data[6][9] ;
wire \myicache.data[7][0] ;
wire \myicache.data[7][10] ;
wire \myicache.data[7][11] ;
wire \myicache.data[7][12] ;
wire \myicache.data[7][13] ;
wire \myicache.data[7][14] ;
wire \myicache.data[7][15] ;
wire \myicache.data[7][16] ;
wire \myicache.data[7][17] ;
wire \myicache.data[7][18] ;
wire \myicache.data[7][19] ;
wire \myicache.data[7][1] ;
wire \myicache.data[7][20] ;
wire \myicache.data[7][21] ;
wire \myicache.data[7][22] ;
wire \myicache.data[7][23] ;
wire \myicache.data[7][24] ;
wire \myicache.data[7][25] ;
wire \myicache.data[7][26] ;
wire \myicache.data[7][27] ;
wire \myicache.data[7][28] ;
wire \myicache.data[7][29] ;
wire \myicache.data[7][2] ;
wire \myicache.data[7][30] ;
wire \myicache.data[7][31] ;
wire \myicache.data[7][3] ;
wire \myicache.data[7][4] ;
wire \myicache.data[7][5] ;
wire \myicache.data[7][6] ;
wire \myicache.data[7][7] ;
wire \myicache.data[7][8] ;
wire \myicache.data[7][9] ;
wire \myicache.tag[0][0] ;
wire \myicache.tag[0][10] ;
wire \myicache.tag[0][11] ;
wire \myicache.tag[0][12] ;
wire \myicache.tag[0][13] ;
wire \myicache.tag[0][14] ;
wire \myicache.tag[0][15] ;
wire \myicache.tag[0][16] ;
wire \myicache.tag[0][17] ;
wire \myicache.tag[0][18] ;
wire \myicache.tag[0][19] ;
wire \myicache.tag[0][1] ;
wire \myicache.tag[0][20] ;
wire \myicache.tag[0][21] ;
wire \myicache.tag[0][22] ;
wire \myicache.tag[0][23] ;
wire \myicache.tag[0][24] ;
wire \myicache.tag[0][25] ;
wire \myicache.tag[0][26] ;
wire \myicache.tag[0][2] ;
wire \myicache.tag[0][3] ;
wire \myicache.tag[0][4] ;
wire \myicache.tag[0][5] ;
wire \myicache.tag[0][6] ;
wire \myicache.tag[0][7] ;
wire \myicache.tag[0][8] ;
wire \myicache.tag[0][9] ;
wire \myicache.tag[1][0] ;
wire \myicache.tag[1][10] ;
wire \myicache.tag[1][11] ;
wire \myicache.tag[1][12] ;
wire \myicache.tag[1][13] ;
wire \myicache.tag[1][14] ;
wire \myicache.tag[1][15] ;
wire \myicache.tag[1][16] ;
wire \myicache.tag[1][17] ;
wire \myicache.tag[1][18] ;
wire \myicache.tag[1][19] ;
wire \myicache.tag[1][1] ;
wire \myicache.tag[1][20] ;
wire \myicache.tag[1][21] ;
wire \myicache.tag[1][22] ;
wire \myicache.tag[1][23] ;
wire \myicache.tag[1][24] ;
wire \myicache.tag[1][25] ;
wire \myicache.tag[1][26] ;
wire \myicache.tag[1][2] ;
wire \myicache.tag[1][3] ;
wire \myicache.tag[1][4] ;
wire \myicache.tag[1][5] ;
wire \myicache.tag[1][6] ;
wire \myicache.tag[1][7] ;
wire \myicache.tag[1][8] ;
wire \myicache.tag[1][9] ;
wire \myicache.tag[2][0] ;
wire \myicache.tag[2][10] ;
wire \myicache.tag[2][11] ;
wire \myicache.tag[2][12] ;
wire \myicache.tag[2][13] ;
wire \myicache.tag[2][14] ;
wire \myicache.tag[2][15] ;
wire \myicache.tag[2][16] ;
wire \myicache.tag[2][17] ;
wire \myicache.tag[2][18] ;
wire \myicache.tag[2][19] ;
wire \myicache.tag[2][1] ;
wire \myicache.tag[2][20] ;
wire \myicache.tag[2][21] ;
wire \myicache.tag[2][22] ;
wire \myicache.tag[2][23] ;
wire \myicache.tag[2][24] ;
wire \myicache.tag[2][25] ;
wire \myicache.tag[2][26] ;
wire \myicache.tag[2][2] ;
wire \myicache.tag[2][3] ;
wire \myicache.tag[2][4] ;
wire \myicache.tag[2][5] ;
wire \myicache.tag[2][6] ;
wire \myicache.tag[2][7] ;
wire \myicache.tag[2][8] ;
wire \myicache.tag[2][9] ;
wire \myicache.tag[3][0] ;
wire \myicache.tag[3][10] ;
wire \myicache.tag[3][11] ;
wire \myicache.tag[3][12] ;
wire \myicache.tag[3][13] ;
wire \myicache.tag[3][14] ;
wire \myicache.tag[3][15] ;
wire \myicache.tag[3][16] ;
wire \myicache.tag[3][17] ;
wire \myicache.tag[3][18] ;
wire \myicache.tag[3][19] ;
wire \myicache.tag[3][1] ;
wire \myicache.tag[3][20] ;
wire \myicache.tag[3][21] ;
wire \myicache.tag[3][22] ;
wire \myicache.tag[3][23] ;
wire \myicache.tag[3][24] ;
wire \myicache.tag[3][25] ;
wire \myicache.tag[3][26] ;
wire \myicache.tag[3][2] ;
wire \myicache.tag[3][3] ;
wire \myicache.tag[3][4] ;
wire \myicache.tag[3][5] ;
wire \myicache.tag[3][6] ;
wire \myicache.tag[3][7] ;
wire \myicache.tag[3][8] ;
wire \myicache.tag[3][9] ;
wire \myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myicache.wen ;
wire pc_$_SDFFE_PP0P__Q_10_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_12_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ORNOT__Y_B_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_12_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_12_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_14_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_14_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_16_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_16_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ;
wire pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B ;
wire pc_$_SDFFE_PP0P__Q_30_E ;
wire pc_$_SDFFE_PP0P__Q_8_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_B ;
wire readyFromIDU_$_AND__B_Y ;
wire rmem_quest_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y ;
wire state_$_DFF_P__Q_1_D ;
wire state_$_DFF_P__Q_2_D ;
wire state_$_DFF_P__Q_D ;
wire tmp_offset_$_SDFFE_PP0P__Q_E ;
wire tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ;
wire to_reset ;
wire wen_$_ANDNOT__A_Y ;
wire wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ;
wire wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ;
wire wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ;
wire wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ;
wire wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ;
wire wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ;
wire wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ;
wire wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire wen_$_ANDNOT__A_Y_$_AND__B_1_Y ;
wire wen_$_ANDNOT__A_Y_$_AND__B_2_Y ;
wire wen_$_ANDNOT__A_Y_$_AND__B_3_Y ;
wire wen_$_ANDNOT__A_Y_$_AND__B_Y ;
wire wen_$_SDFFE_PP0P__Q_E ;
wire fanout_net_1 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire [31:0] pc_jump ;
wire [31:0] mtvec ;
wire [31:0] pc ;
wire [31:0] inst ;
wire [31:0] araddr ;
wire [3:0] arid ;
wire [7:0] arlen ;
wire [2:0] arsize ;
wire [1:0] arburst ;
wire [31:0] rdata ;
wire [1:0] rresp ;
wire [3:0] rid ;
wire [3:0] \myicache.valid ;
wire [1:0] pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y ;
wire [2:0] state ;
wire [2:0] tmp_offset ;

assign \pc [3] = \araddr [3] ;
assign \pc [4] = \araddr [4] ;
assign \pc [5] = \araddr [5] ;
assign \pc [6] = \araddr [6] ;
assign \pc [7] = \araddr [7] ;
assign \pc [8] = \araddr [8] ;
assign \pc [9] = \araddr [9] ;
assign \pc [10] = \araddr [10] ;
assign \pc [11] = \araddr [11] ;
assign \pc [12] = \araddr [12] ;
assign \pc [13] = \araddr [13] ;
assign \pc [14] = \araddr [14] ;
assign \pc [15] = \araddr [15] ;
assign \pc [16] = \araddr [16] ;
assign \pc [17] = \araddr [17] ;
assign \pc [18] = \araddr [18] ;
assign \pc [19] = \araddr [19] ;
assign \pc [20] = \araddr [20] ;
assign \pc [21] = \araddr [21] ;
assign \pc [22] = \araddr [22] ;
assign \pc [23] = \araddr [23] ;
assign \pc [24] = \araddr [24] ;
assign \pc [25] = \araddr [25] ;
assign \pc [26] = \araddr [26] ;
assign \pc [27] = \araddr [27] ;
assign \pc [28] = \araddr [28] ;
assign \pc [29] = \araddr [29] ;
assign \pc [30] = \araddr [30] ;
assign \pc [31] = \araddr [31] ;
assign \araddr [1] = \araddr [0] ;
assign \araddr [2] = \araddr [0] ;
assign \arid [0] = \arburst [0] ;
assign \arid [1] = \araddr [0] ;
assign \arid [2] = \araddr [0] ;
assign \arid [3] = \araddr [0] ;
assign \arlen [0] = \arburst [0] ;
assign \arlen [1] = \araddr [0] ;
assign \arlen [2] = \araddr [0] ;
assign \arlen [3] = \araddr [0] ;
assign \arlen [4] = \araddr [0] ;
assign \arlen [5] = \araddr [0] ;
assign \arlen [6] = \araddr [0] ;
assign \arlen [7] = \araddr [0] ;
assign \arsize [0] = \araddr [0] ;
assign \arsize [1] = \arburst [0] ;
assign \arsize [2] = \araddr [0] ;
assign \arburst [1] = \araddr [0] ;

NOR2_X4 _1632_ ( .A1(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(\inst [4] ), .ZN(_0888_ ) );
AND2_X4 _1633_ ( .A1(_0888_ ), .A2(\inst [5] ), .ZN(_0889_ ) );
INV_X8 _1634_ ( .A(_0889_ ), .ZN(_0890_ ) );
NOR2_X4 _1635_ ( .A1(\inst [3] ), .A2(\inst [2] ), .ZN(_0891_ ) );
NAND4_X4 _1636_ ( .A1(_0891_ ), .A2(\inst [1] ), .A3(\inst [0] ), .A4(\inst [31] ), .ZN(_0892_ ) );
NOR2_X4 _1637_ ( .A1(_0890_ ), .A2(_0892_ ), .ZN(_0893_ ) );
AND4_X4 _1638_ ( .A1(\inst [3] ), .A2(\inst [2] ), .A3(\inst [1] ), .A4(\inst [0] ), .ZN(_0894_ ) );
AND2_X4 _1639_ ( .A1(_0889_ ), .A2(_0894_ ), .ZN(_0895_ ) );
NOR2_X4 _1640_ ( .A1(_0893_ ), .A2(_0895_ ), .ZN(_0896_ ) );
NOR2_X4 _1641_ ( .A1(_0896_ ), .A2(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_0897_ ) );
BUF_X4 _1642_ ( .A(_0897_ ), .Z(_0898_ ) );
XOR2_X1 _1643_ ( .A(_0898_ ), .B(\araddr [28] ), .Z(_0899_ ) );
INV_X1 _1644_ ( .A(\araddr [27] ), .ZN(_0900_ ) );
XNOR2_X1 _1645_ ( .A(_0898_ ), .B(_0900_ ), .ZN(_0901_ ) );
AND2_X1 _1646_ ( .A1(_0899_ ), .A2(_0901_ ), .ZN(_0902_ ) );
BUF_X4 _1647_ ( .A(_0898_ ), .Z(_0903_ ) );
INV_X1 _1648_ ( .A(\araddr [26] ), .ZN(_0904_ ) );
XNOR2_X1 _1649_ ( .A(_0903_ ), .B(_0904_ ), .ZN(_0905_ ) );
INV_X1 _1650_ ( .A(\araddr [25] ), .ZN(_0906_ ) );
XNOR2_X1 _1651_ ( .A(_0898_ ), .B(_0906_ ), .ZN(_0907_ ) );
AND2_X1 _1652_ ( .A1(_0905_ ), .A2(_0907_ ), .ZN(_0908_ ) );
AND2_X4 _1653_ ( .A1(_0893_ ), .A2(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_0909_ ) );
INV_X8 _1654_ ( .A(_0895_ ), .ZN(_0910_ ) );
BUF_X8 _1655_ ( .A(_0910_ ), .Z(_0911_ ) );
OR2_X1 _1656_ ( .A1(_0911_ ), .A2(pc_$_SDFFE_PP0P__Q_14_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0912_ ) );
INV_X2 _1657_ ( .A(_0893_ ), .ZN(_0913_ ) );
AOI21_X1 _1658_ ( .A(_0909_ ), .B1(_0912_ ), .B2(_0913_ ), .ZN(_0914_ ) );
XOR2_X2 _1659_ ( .A(_0914_ ), .B(\araddr [16] ), .Z(_0915_ ) );
OR2_X4 _1660_ ( .A1(_0911_ ), .A2(pc_$_SDFFE_PP0P__Q_14_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0916_ ) );
AOI21_X2 _1661_ ( .A(_0909_ ), .B1(_0916_ ), .B2(_0913_ ), .ZN(_0917_ ) );
INV_X1 _1662_ ( .A(\araddr [15] ), .ZN(_0918_ ) );
XNOR2_X2 _1663_ ( .A(_0917_ ), .B(_0918_ ), .ZN(_0919_ ) );
NAND2_X1 _1664_ ( .A1(_0915_ ), .A2(_0919_ ), .ZN(_0920_ ) );
NAND2_X4 _1665_ ( .A1(_0893_ ), .A2(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_0921_ ) );
NOR2_X1 _1666_ ( .A1(_0911_ ), .A2(pc_$_SDFFE_PP0P__Q_16_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0922_ ) );
OAI21_X1 _1667_ ( .A(_0921_ ), .B1(_0922_ ), .B2(_0893_ ), .ZN(_0923_ ) );
XNOR2_X1 _1668_ ( .A(_0923_ ), .B(\araddr [13] ), .ZN(_0924_ ) );
OAI22_X1 _1669_ ( .A1(_0910_ ), .A2(pc_$_SDFFE_PP0P__Q_16_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .B1(_0890_ ), .B2(_0892_ ), .ZN(_0925_ ) );
AND2_X1 _1670_ ( .A1(_0925_ ), .A2(_0921_ ), .ZN(_0926_ ) );
OR2_X2 _1671_ ( .A1(_0926_ ), .A2(\araddr [14] ), .ZN(_0927_ ) );
NAND3_X1 _1672_ ( .A1(_0925_ ), .A2(\araddr [14] ), .A3(_0921_ ), .ZN(_0928_ ) );
NAND3_X1 _1673_ ( .A1(_0924_ ), .A2(_0927_ ), .A3(_0928_ ), .ZN(_0929_ ) );
NOR2_X1 _1674_ ( .A1(_0920_ ), .A2(_0929_ ), .ZN(_0930_ ) );
AOI21_X1 _1675_ ( .A(pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B1(_0913_ ), .B2(_0910_ ), .ZN(_0931_ ) );
XOR2_X1 _1676_ ( .A(_0931_ ), .B(\araddr [9] ), .Z(_0932_ ) );
INV_X1 _1677_ ( .A(pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_0933_ ) );
OAI21_X1 _1678_ ( .A(_0933_ ), .B1(_0893_ ), .B2(_0895_ ), .ZN(_0934_ ) );
XNOR2_X1 _1679_ ( .A(_0934_ ), .B(\araddr [10] ), .ZN(_0935_ ) );
AND2_X1 _1680_ ( .A1(_0932_ ), .A2(_0935_ ), .ZN(_0936_ ) );
NOR2_X1 _1681_ ( .A1(_0910_ ), .A2(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0937_ ) );
OAI21_X1 _1682_ ( .A(_0921_ ), .B1(_0937_ ), .B2(_0893_ ), .ZN(_0938_ ) );
XNOR2_X1 _1683_ ( .A(_0938_ ), .B(\araddr [12] ), .ZN(_0939_ ) );
OR3_X1 _1684_ ( .A1(_0890_ ), .A2(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_0892_ ), .ZN(_0940_ ) );
OAI21_X1 _1685_ ( .A(_0940_ ), .B1(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ), .B2(_0911_ ), .ZN(_0941_ ) );
XOR2_X1 _1686_ ( .A(_0941_ ), .B(\araddr [11] ), .Z(_0942_ ) );
AND3_X1 _1687_ ( .A1(_0936_ ), .A2(_0939_ ), .A3(_0942_ ), .ZN(_0943_ ) );
OR3_X4 _1688_ ( .A1(_0890_ ), .A2(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_0892_ ), .ZN(_0944_ ) );
OAI21_X4 _1689_ ( .A(_0944_ ), .B1(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .B2(_0910_ ), .ZN(_0945_ ) );
INV_X1 _1690_ ( .A(\araddr [4] ), .ZN(_0946_ ) );
XNOR2_X2 _1691_ ( .A(_0945_ ), .B(_0946_ ), .ZN(_0947_ ) );
NOR2_X1 _1692_ ( .A1(_0910_ ), .A2(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0948_ ) );
NOR3_X1 _1693_ ( .A1(_0890_ ), .A2(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .A3(_0892_ ), .ZN(_0949_ ) );
NOR2_X1 _1694_ ( .A1(_0948_ ), .A2(_0949_ ), .ZN(_0950_ ) );
NOR2_X1 _1695_ ( .A1(_0950_ ), .A2(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_0951_ ) );
AND2_X1 _1696_ ( .A1(_0947_ ), .A2(_0951_ ), .ZN(_0952_ ) );
AOI21_X1 _1697_ ( .A(_0952_ ), .B1(\araddr [4] ), .B2(_0945_ ), .ZN(_0953_ ) );
INV_X1 _1698_ ( .A(_0953_ ), .ZN(_0954_ ) );
INV_X1 _1699_ ( .A(pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_0955_ ) );
NOR3_X2 _1700_ ( .A1(_0890_ ), .A2(_0955_ ), .A3(_0892_ ), .ZN(_0956_ ) );
AND4_X1 _1701_ ( .A1(pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .A2(_0894_ ), .A3(\inst [5] ), .A4(_0888_ ), .ZN(_0957_ ) );
NOR2_X1 _1702_ ( .A1(_0956_ ), .A2(_0957_ ), .ZN(_0958_ ) );
INV_X1 _1703_ ( .A(\pc [2] ), .ZN(_0959_ ) );
XNOR2_X1 _1704_ ( .A(_0958_ ), .B(_0959_ ), .ZN(_0960_ ) );
NOR2_X1 _1705_ ( .A1(_0910_ ), .A2(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0961_ ) );
NOR3_X1 _1706_ ( .A1(_0890_ ), .A2(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_0892_ ), .ZN(_0962_ ) );
NOR2_X1 _1707_ ( .A1(_0961_ ), .A2(_0962_ ), .ZN(_0963_ ) );
NOR2_X1 _1708_ ( .A1(_0963_ ), .A2(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B ), .ZN(_0964_ ) );
AND2_X2 _1709_ ( .A1(_0960_ ), .A2(_0964_ ), .ZN(_0965_ ) );
NOR3_X1 _1710_ ( .A1(_0956_ ), .A2(_0959_ ), .A3(_0957_ ), .ZN(_0966_ ) );
NOR2_X2 _1711_ ( .A1(_0965_ ), .A2(_0966_ ), .ZN(_0967_ ) );
INV_X1 _1712_ ( .A(_0947_ ), .ZN(_0968_ ) );
INV_X1 _1713_ ( .A(\araddr [3] ), .ZN(_0969_ ) );
XNOR2_X1 _1714_ ( .A(_0950_ ), .B(_0969_ ), .ZN(_0970_ ) );
NOR3_X4 _1715_ ( .A1(_0967_ ), .A2(_0968_ ), .A3(_0970_ ), .ZN(_0971_ ) );
NOR2_X4 _1716_ ( .A1(_0954_ ), .A2(_0971_ ), .ZN(_0972_ ) );
AOI21_X4 _1717_ ( .A(pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B1(_0913_ ), .B2(_0911_ ), .ZN(_0973_ ) );
XOR2_X1 _1718_ ( .A(_0973_ ), .B(\araddr [8] ), .Z(_0974_ ) );
INV_X1 _1719_ ( .A(_0974_ ), .ZN(_0975_ ) );
AOI21_X2 _1720_ ( .A(pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B1(_0913_ ), .B2(_0911_ ), .ZN(_0976_ ) );
XOR2_X2 _1721_ ( .A(_0976_ ), .B(\araddr [7] ), .Z(_0977_ ) );
INV_X1 _1722_ ( .A(_0977_ ), .ZN(_0978_ ) );
NOR2_X4 _1723_ ( .A1(_0896_ ), .A2(pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_0979_ ) );
XNOR2_X2 _1724_ ( .A(_0979_ ), .B(\araddr [5] ), .ZN(_0980_ ) );
INV_X4 _1725_ ( .A(_0896_ ), .ZN(_0981_ ) );
INV_X1 _1726_ ( .A(pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_0982_ ) );
AOI21_X2 _1727_ ( .A(\araddr [6] ), .B1(_0981_ ), .B2(_0982_ ), .ZN(_0983_ ) );
AND3_X4 _1728_ ( .A1(_0981_ ), .A2(\araddr [6] ), .A3(_0982_ ), .ZN(_0984_ ) );
NOR3_X2 _1729_ ( .A1(_0980_ ), .A2(_0983_ ), .A3(_0984_ ), .ZN(_0985_ ) );
INV_X1 _1730_ ( .A(_0985_ ), .ZN(_0986_ ) );
NOR4_X4 _1731_ ( .A1(_0972_ ), .A2(_0975_ ), .A3(_0978_ ), .A4(_0986_ ), .ZN(_0987_ ) );
OR3_X4 _1732_ ( .A1(_0896_ ), .A2(pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .A3(pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_0988_ ) );
NOR3_X2 _1733_ ( .A1(_0984_ ), .A2(_0983_ ), .A3(_0988_ ), .ZN(_0989_ ) );
OR2_X4 _1734_ ( .A1(_0989_ ), .A2(_0984_ ), .ZN(_0990_ ) );
AND3_X4 _1735_ ( .A1(_0990_ ), .A2(_0974_ ), .A3(_0977_ ), .ZN(_0991_ ) );
AND2_X1 _1736_ ( .A1(_0973_ ), .A2(\araddr [8] ), .ZN(_0992_ ) );
AND2_X1 _1737_ ( .A1(_0976_ ), .A2(\araddr [7] ), .ZN(_0993_ ) );
AND2_X1 _1738_ ( .A1(_0974_ ), .A2(_0993_ ), .ZN(_0994_ ) );
OR3_X4 _1739_ ( .A1(_0991_ ), .A2(_0992_ ), .A3(_0994_ ), .ZN(_0995_ ) );
OAI211_X2 _1740_ ( .A(_0930_ ), .B(_0943_ ), .C1(_0987_ ), .C2(_0995_ ), .ZN(_0996_ ) );
AND2_X1 _1741_ ( .A1(_0931_ ), .A2(\araddr [9] ), .ZN(_0997_ ) );
AND2_X1 _1742_ ( .A1(_0935_ ), .A2(_0997_ ), .ZN(_0998_ ) );
AND3_X1 _1743_ ( .A1(_0981_ ), .A2(\araddr [10] ), .A3(_0933_ ), .ZN(_0999_ ) );
OAI211_X1 _1744_ ( .A(_0939_ ), .B(_0942_ ), .C1(_0998_ ), .C2(_0999_ ), .ZN(_1000_ ) );
INV_X1 _1745_ ( .A(\araddr [12] ), .ZN(_1001_ ) );
NOR2_X1 _1746_ ( .A1(_0938_ ), .A2(_1001_ ), .ZN(_1002_ ) );
AND2_X1 _1747_ ( .A1(_0941_ ), .A2(\araddr [11] ), .ZN(_1003_ ) );
AOI21_X1 _1748_ ( .A(_1002_ ), .B1(_0939_ ), .B2(_1003_ ), .ZN(_1004_ ) );
AND2_X1 _1749_ ( .A1(_1000_ ), .A2(_1004_ ), .ZN(_1005_ ) );
NOR3_X1 _1750_ ( .A1(_1005_ ), .A2(_0920_ ), .A3(_0929_ ), .ZN(_1006_ ) );
AND2_X1 _1751_ ( .A1(_0914_ ), .A2(\araddr [16] ), .ZN(_1007_ ) );
INV_X1 _1752_ ( .A(\araddr [13] ), .ZN(_1008_ ) );
OAI21_X1 _1753_ ( .A(_0928_ ), .B1(_0923_ ), .B2(_1008_ ), .ZN(_1009_ ) );
AND2_X1 _1754_ ( .A1(_0927_ ), .A2(_1009_ ), .ZN(_1010_ ) );
AND3_X1 _1755_ ( .A1(_1010_ ), .A2(_0915_ ), .A3(_0919_ ), .ZN(_1011_ ) );
AND2_X1 _1756_ ( .A1(_0917_ ), .A2(\araddr [15] ), .ZN(_1012_ ) );
AND2_X1 _1757_ ( .A1(_0915_ ), .A2(_1012_ ), .ZN(_1013_ ) );
NOR4_X2 _1758_ ( .A1(_1006_ ), .A2(_1007_ ), .A3(_1011_ ), .A4(_1013_ ), .ZN(_1014_ ) );
AND2_X2 _1759_ ( .A1(_0996_ ), .A2(_1014_ ), .ZN(_1015_ ) );
INV_X2 _1760_ ( .A(_1015_ ), .ZN(_1016_ ) );
INV_X1 _1761_ ( .A(\araddr [21] ), .ZN(_1017_ ) );
XNOR2_X1 _1762_ ( .A(_0897_ ), .B(_1017_ ), .ZN(_1018_ ) );
XNOR2_X1 _1763_ ( .A(_0897_ ), .B(pc_$_SDFFE_PP0P__Q_8_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_1019_ ) );
AND2_X1 _1764_ ( .A1(_1018_ ), .A2(_1019_ ), .ZN(_1020_ ) );
INV_X1 _1765_ ( .A(_1020_ ), .ZN(_1021_ ) );
INV_X1 _1766_ ( .A(\araddr [23] ), .ZN(_1022_ ) );
XNOR2_X1 _1767_ ( .A(_0897_ ), .B(_1022_ ), .ZN(_1023_ ) );
INV_X1 _1768_ ( .A(_1023_ ), .ZN(_1024_ ) );
XNOR2_X1 _1769_ ( .A(_0898_ ), .B(\araddr [24] ), .ZN(_1025_ ) );
NOR3_X1 _1770_ ( .A1(_1021_ ), .A2(_1024_ ), .A3(_1025_ ), .ZN(_1026_ ) );
OAI22_X1 _1771_ ( .A1(_0911_ ), .A2(pc_$_SDFFE_PP0P__Q_12_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .B1(_0890_ ), .B2(_0892_ ), .ZN(_1027_ ) );
AND2_X2 _1772_ ( .A1(_1027_ ), .A2(_0921_ ), .ZN(_1028_ ) );
XNOR2_X2 _1773_ ( .A(_1028_ ), .B(pc_$_SDFFE_PP0P__Q_12_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_1029_ ) );
NOR2_X1 _1774_ ( .A1(_0911_ ), .A2(pc_$_SDFFE_PP0P__Q_12_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ORNOT__Y_B_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_1030_ ) );
OAI21_X1 _1775_ ( .A(_0921_ ), .B1(_1030_ ), .B2(_0893_ ), .ZN(_1031_ ) );
XNOR2_X1 _1776_ ( .A(_1031_ ), .B(\araddr [17] ), .ZN(_1032_ ) );
AND2_X1 _1777_ ( .A1(_1029_ ), .A2(_1032_ ), .ZN(_1033_ ) );
INV_X1 _1778_ ( .A(\araddr [20] ), .ZN(_1034_ ) );
XNOR2_X1 _1779_ ( .A(_0897_ ), .B(_1034_ ), .ZN(_1035_ ) );
OR2_X1 _1780_ ( .A1(_0911_ ), .A2(pc_$_SDFFE_PP0P__Q_10_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_1036_ ) );
AOI21_X1 _1781_ ( .A(_0909_ ), .B1(_1036_ ), .B2(_0913_ ), .ZN(_1037_ ) );
XOR2_X1 _1782_ ( .A(_1037_ ), .B(\araddr [19] ), .Z(_1038_ ) );
AND3_X1 _1783_ ( .A1(_1033_ ), .A2(_1035_ ), .A3(_1038_ ), .ZN(_1039_ ) );
AND3_X4 _1784_ ( .A1(_1016_ ), .A2(_1026_ ), .A3(_1039_ ), .ZN(_1040_ ) );
NAND2_X1 _1785_ ( .A1(_0898_ ), .A2(\araddr [23] ), .ZN(_1041_ ) );
OAI22_X1 _1786_ ( .A1(_0911_ ), .A2(pc_$_SDFFE_PP0P__Q_12_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ORNOT__Y_B_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ), .B1(_0890_ ), .B2(_0892_ ), .ZN(_1042_ ) );
AND3_X1 _1787_ ( .A1(_1042_ ), .A2(\araddr [17] ), .A3(_0921_ ), .ZN(_1043_ ) );
AND2_X2 _1788_ ( .A1(_1029_ ), .A2(_1043_ ), .ZN(_1044_ ) );
AOI21_X1 _1789_ ( .A(_1044_ ), .B1(\araddr [18] ), .B2(_1028_ ), .ZN(_1045_ ) );
INV_X1 _1790_ ( .A(_1038_ ), .ZN(_1046_ ) );
INV_X1 _1791_ ( .A(_1035_ ), .ZN(_1047_ ) );
NOR3_X2 _1792_ ( .A1(_1045_ ), .A2(_1046_ ), .A3(_1047_ ), .ZN(_1048_ ) );
AND2_X1 _1793_ ( .A1(_1037_ ), .A2(\araddr [19] ), .ZN(_1049_ ) );
AND2_X1 _1794_ ( .A1(_1049_ ), .A2(_1035_ ), .ZN(_1050_ ) );
AOI21_X1 _1795_ ( .A(_1050_ ), .B1(\araddr [20] ), .B2(_0898_ ), .ZN(_1051_ ) );
INV_X1 _1796_ ( .A(_1051_ ), .ZN(_1052_ ) );
OAI21_X1 _1797_ ( .A(_1026_ ), .B1(_1048_ ), .B2(_1052_ ), .ZN(_1053_ ) );
NAND2_X1 _1798_ ( .A1(_0898_ ), .A2(\araddr [24] ), .ZN(_1054_ ) );
AND3_X1 _1799_ ( .A1(_0897_ ), .A2(\araddr [21] ), .A3(pc_$_SDFFE_PP0P__Q_8_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_1055_ ) );
AOI21_X1 _1800_ ( .A(_1055_ ), .B1(\araddr [22] ), .B2(_0898_ ), .ZN(_1056_ ) );
OR3_X1 _1801_ ( .A1(_1056_ ), .A2(_1024_ ), .A3(_1025_ ), .ZN(_1057_ ) );
AND4_X2 _1802_ ( .A1(_1041_ ), .A2(_1053_ ), .A3(_1054_ ), .A4(_1057_ ), .ZN(_1058_ ) );
INV_X1 _1803_ ( .A(_1058_ ), .ZN(_1059_ ) );
OAI211_X1 _1804_ ( .A(_0902_ ), .B(_0908_ ), .C1(_1040_ ), .C2(_1059_ ), .ZN(_1060_ ) );
NOR4_X1 _1805_ ( .A1(_0896_ ), .A2(\araddr [28] ), .A3(_0900_ ), .A4(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_1061_ ) );
NAND2_X1 _1806_ ( .A1(_0898_ ), .A2(\araddr [25] ), .ZN(_1062_ ) );
OR3_X1 _1807_ ( .A1(_0896_ ), .A2(_0904_ ), .A3(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_1063_ ) );
NAND2_X1 _1808_ ( .A1(_1062_ ), .A2(_1063_ ), .ZN(_1064_ ) );
AOI221_X4 _1809_ ( .A(_1061_ ), .B1(\araddr [28] ), .B2(_0903_ ), .C1(_0902_ ), .C2(_1064_ ), .ZN(_1065_ ) );
AND2_X2 _1810_ ( .A1(_1060_ ), .A2(_1065_ ), .ZN(_1066_ ) );
XOR2_X1 _1811_ ( .A(_0903_ ), .B(\araddr [29] ), .Z(_1067_ ) );
INV_X1 _1812_ ( .A(_1067_ ), .ZN(_1068_ ) );
NOR2_X1 _1813_ ( .A1(_1066_ ), .A2(_1068_ ), .ZN(_1069_ ) );
AND2_X1 _1814_ ( .A1(_0903_ ), .A2(\araddr [29] ), .ZN(_1070_ ) );
XNOR2_X1 _1815_ ( .A(_0903_ ), .B(\araddr [30] ), .ZN(_1071_ ) );
OR3_X2 _1816_ ( .A1(_1069_ ), .A2(_1070_ ), .A3(_1071_ ), .ZN(_1072_ ) );
XNOR2_X1 _1817_ ( .A(\pc_jump [0] ), .B(\pc [0] ), .ZN(_1073_ ) );
XNOR2_X1 _1818_ ( .A(\pc_jump [3] ), .B(\araddr [3] ), .ZN(_1074_ ) );
XNOR2_X1 _1819_ ( .A(\pc_jump [2] ), .B(\pc [2] ), .ZN(_1075_ ) );
XNOR2_X1 _1820_ ( .A(\pc_jump [1] ), .B(\pc [1] ), .ZN(_1076_ ) );
AND4_X1 _1821_ ( .A1(_1073_ ), .A2(_1074_ ), .A3(_1075_ ), .A4(_1076_ ), .ZN(_1077_ ) );
XNOR2_X1 _1822_ ( .A(\pc_jump [6] ), .B(\araddr [6] ), .ZN(_1078_ ) );
XNOR2_X1 _1823_ ( .A(\pc_jump [5] ), .B(\araddr [5] ), .ZN(_1079_ ) );
XNOR2_X1 _1824_ ( .A(\pc_jump [7] ), .B(\araddr [7] ), .ZN(_1080_ ) );
XNOR2_X1 _1825_ ( .A(\pc_jump [4] ), .B(\araddr [4] ), .ZN(_1081_ ) );
AND4_X1 _1826_ ( .A1(_1078_ ), .A2(_1079_ ), .A3(_1080_ ), .A4(_1081_ ), .ZN(_1082_ ) );
XNOR2_X1 _1827_ ( .A(\pc_jump [15] ), .B(\araddr [15] ), .ZN(_1083_ ) );
XNOR2_X1 _1828_ ( .A(\pc_jump [12] ), .B(\araddr [12] ), .ZN(_1084_ ) );
XNOR2_X1 _1829_ ( .A(\pc_jump [14] ), .B(\araddr [14] ), .ZN(_1085_ ) );
XNOR2_X1 _1830_ ( .A(\pc_jump [13] ), .B(\araddr [13] ), .ZN(_1086_ ) );
AND4_X1 _1831_ ( .A1(_1083_ ), .A2(_1084_ ), .A3(_1085_ ), .A4(_1086_ ), .ZN(_1087_ ) );
XNOR2_X1 _1832_ ( .A(\pc_jump [8] ), .B(\araddr [8] ), .ZN(_1088_ ) );
XNOR2_X1 _1833_ ( .A(\pc_jump [9] ), .B(\araddr [9] ), .ZN(_1089_ ) );
XNOR2_X1 _1834_ ( .A(\pc_jump [10] ), .B(\araddr [10] ), .ZN(_1090_ ) );
XNOR2_X1 _1835_ ( .A(\pc_jump [11] ), .B(\araddr [11] ), .ZN(_1091_ ) );
AND4_X1 _1836_ ( .A1(_1088_ ), .A2(_1089_ ), .A3(_1090_ ), .A4(_1091_ ), .ZN(_1092_ ) );
AND4_X1 _1837_ ( .A1(_1077_ ), .A2(_1082_ ), .A3(_1087_ ), .A4(_1092_ ), .ZN(_1093_ ) );
XNOR2_X1 _1838_ ( .A(\pc_jump [30] ), .B(\araddr [30] ), .ZN(_1094_ ) );
XNOR2_X1 _1839_ ( .A(\pc_jump [31] ), .B(\araddr [31] ), .ZN(_1095_ ) );
XNOR2_X1 _1840_ ( .A(\pc_jump [28] ), .B(\araddr [28] ), .ZN(_1096_ ) );
XNOR2_X1 _1841_ ( .A(\pc_jump [29] ), .B(\araddr [29] ), .ZN(_1097_ ) );
AND4_X1 _1842_ ( .A1(_1094_ ), .A2(_1095_ ), .A3(_1096_ ), .A4(_1097_ ), .ZN(_1098_ ) );
XNOR2_X1 _1843_ ( .A(\pc_jump [24] ), .B(\araddr [24] ), .ZN(_1099_ ) );
XNOR2_X1 _1844_ ( .A(\pc_jump [26] ), .B(\araddr [26] ), .ZN(_1100_ ) );
XNOR2_X1 _1845_ ( .A(\pc_jump [27] ), .B(\araddr [27] ), .ZN(_1101_ ) );
XNOR2_X1 _1846_ ( .A(\pc_jump [25] ), .B(\araddr [25] ), .ZN(_1102_ ) );
AND4_X1 _1847_ ( .A1(_1099_ ), .A2(_1100_ ), .A3(_1101_ ), .A4(_1102_ ), .ZN(_1103_ ) );
XNOR2_X1 _1848_ ( .A(\pc_jump [18] ), .B(\araddr [18] ), .ZN(_1104_ ) );
XNOR2_X1 _1849_ ( .A(\pc_jump [16] ), .B(\araddr [16] ), .ZN(_1105_ ) );
XNOR2_X1 _1850_ ( .A(\pc_jump [19] ), .B(\araddr [19] ), .ZN(_1106_ ) );
XNOR2_X1 _1851_ ( .A(\pc_jump [17] ), .B(\araddr [17] ), .ZN(_1107_ ) );
NAND4_X1 _1852_ ( .A1(_1104_ ), .A2(_1105_ ), .A3(_1106_ ), .A4(_1107_ ), .ZN(_1108_ ) );
XNOR2_X1 _1853_ ( .A(\pc_jump [23] ), .B(\araddr [23] ), .ZN(_1109_ ) );
XNOR2_X1 _1854_ ( .A(\pc_jump [22] ), .B(\araddr [22] ), .ZN(_1110_ ) );
NAND2_X1 _1855_ ( .A1(_1109_ ), .A2(_1110_ ), .ZN(_1111_ ) );
XOR2_X1 _1856_ ( .A(\pc_jump [20] ), .B(\araddr [20] ), .Z(_1112_ ) );
XOR2_X1 _1857_ ( .A(\pc_jump [21] ), .B(\araddr [21] ), .Z(_1113_ ) );
NOR4_X1 _1858_ ( .A1(_1108_ ), .A2(_1111_ ), .A3(_1112_ ), .A4(_1113_ ), .ZN(_1114_ ) );
NAND4_X1 _1859_ ( .A1(_1093_ ), .A2(_1098_ ), .A3(_1103_ ), .A4(_1114_ ), .ZN(_1115_ ) );
AND2_X2 _1860_ ( .A1(_1115_ ), .A2(check_quest ), .ZN(_1116_ ) );
INV_X1 _1861_ ( .A(_1116_ ), .ZN(_1117_ ) );
BUF_X4 _1862_ ( .A(_1117_ ), .Z(_1118_ ) );
OAI21_X1 _1863_ ( .A(_1071_ ), .B1(_1069_ ), .B2(_1070_ ), .ZN(_1119_ ) );
NAND3_X1 _1864_ ( .A1(_1072_ ), .A2(_1118_ ), .A3(_1119_ ), .ZN(_1120_ ) );
INV_X2 _1865_ ( .A(fanout_net_11 ), .ZN(_1121_ ) );
BUF_X4 _1866_ ( .A(_1121_ ), .Z(_1122_ ) );
BUF_X4 _1867_ ( .A(_1118_ ), .Z(_1123_ ) );
OAI211_X1 _1868_ ( .A(_1120_ ), .B(_1122_ ), .C1(\pc_jump [30] ), .C2(_1123_ ), .ZN(_1124_ ) );
NAND2_X1 _1869_ ( .A1(fanout_net_11 ), .A2(\mtvec [30] ), .ZN(_1125_ ) );
AOI21_X1 _1870_ ( .A(fanout_net_1 ), .B1(_1124_ ), .B2(_1125_ ), .ZN(_0003_ ) );
NOR2_X1 _1871_ ( .A1(_1121_ ), .A2(\mtvec [29] ), .ZN(_1126_ ) );
BUF_X4 _1872_ ( .A(_1116_ ), .Z(_1127_ ) );
AND3_X1 _1873_ ( .A1(_1060_ ), .A2(_1065_ ), .A3(_1068_ ), .ZN(_1128_ ) );
OR3_X1 _1874_ ( .A1(_1069_ ), .A2(_1127_ ), .A3(_1128_ ), .ZN(_1129_ ) );
BUF_X4 _1875_ ( .A(_1127_ ), .Z(_1130_ ) );
AOI21_X1 _1876_ ( .A(fanout_net_11 ), .B1(_1130_ ), .B2(\pc_jump [29] ), .ZN(_1131_ ) );
AOI211_X1 _1877_ ( .A(fanout_net_1 ), .B(_1126_ ), .C1(_1129_ ), .C2(_1131_ ), .ZN(_0004_ ) );
NAND2_X1 _1878_ ( .A1(_1016_ ), .A2(_1033_ ), .ZN(_1132_ ) );
AOI21_X1 _1879_ ( .A(_1046_ ), .B1(_1132_ ), .B2(_1045_ ), .ZN(_1133_ ) );
OR3_X1 _1880_ ( .A1(_1133_ ), .A2(_1047_ ), .A3(_1049_ ), .ZN(_1134_ ) );
OAI21_X1 _1881_ ( .A(_1047_ ), .B1(_1133_ ), .B2(_1049_ ), .ZN(_1135_ ) );
AOI21_X1 _1882_ ( .A(_1127_ ), .B1(_1134_ ), .B2(_1135_ ), .ZN(_1136_ ) );
AOI211_X1 _1883_ ( .A(fanout_net_11 ), .B(_1136_ ), .C1(\pc_jump [20] ), .C2(_1130_ ), .ZN(_1137_ ) );
BUF_X4 _1884_ ( .A(_1121_ ), .Z(_1138_ ) );
NOR2_X1 _1885_ ( .A1(_1138_ ), .A2(\mtvec [20] ), .ZN(_1139_ ) );
NOR3_X1 _1886_ ( .A1(_1137_ ), .A2(fanout_net_1 ), .A3(_1139_ ), .ZN(_0005_ ) );
AND3_X1 _1887_ ( .A1(_1132_ ), .A2(_1046_ ), .A3(_1045_ ), .ZN(_1140_ ) );
NOR3_X1 _1888_ ( .A1(_1140_ ), .A2(_1133_ ), .A3(_1127_ ), .ZN(_1141_ ) );
AOI211_X1 _1889_ ( .A(fanout_net_11 ), .B(_1141_ ), .C1(\pc_jump [19] ), .C2(_1130_ ), .ZN(_1142_ ) );
NOR2_X1 _1890_ ( .A1(_1138_ ), .A2(\mtvec [19] ), .ZN(_1143_ ) );
NOR3_X1 _1891_ ( .A1(_1142_ ), .A2(fanout_net_1 ), .A3(_1143_ ), .ZN(_0006_ ) );
INV_X1 _1892_ ( .A(_1032_ ), .ZN(_1144_ ) );
AOI21_X1 _1893_ ( .A(_1144_ ), .B1(_0996_ ), .B2(_1014_ ), .ZN(_1145_ ) );
OR2_X1 _1894_ ( .A1(_1145_ ), .A2(_1043_ ), .ZN(_1146_ ) );
OAI21_X1 _1895_ ( .A(_1117_ ), .B1(_1146_ ), .B2(_1029_ ), .ZN(_1147_ ) );
AOI21_X1 _1896_ ( .A(_1147_ ), .B1(_1029_ ), .B2(_1146_ ), .ZN(_1148_ ) );
AOI211_X1 _1897_ ( .A(fanout_net_11 ), .B(_1148_ ), .C1(\pc_jump [18] ), .C2(_1130_ ), .ZN(_1149_ ) );
NOR2_X1 _1898_ ( .A1(_1138_ ), .A2(\mtvec [18] ), .ZN(_1150_ ) );
NOR3_X1 _1899_ ( .A1(_1149_ ), .A2(fanout_net_1 ), .A3(_1150_ ), .ZN(_0007_ ) );
AND3_X1 _1900_ ( .A1(_0996_ ), .A2(_1014_ ), .A3(_1144_ ), .ZN(_1151_ ) );
NOR3_X1 _1901_ ( .A1(_1151_ ), .A2(_1145_ ), .A3(_1127_ ), .ZN(_1152_ ) );
AOI211_X1 _1902_ ( .A(fanout_net_11 ), .B(_1152_ ), .C1(\pc_jump [17] ), .C2(_1130_ ), .ZN(_1153_ ) );
NOR2_X1 _1903_ ( .A1(_1138_ ), .A2(\mtvec [17] ), .ZN(_1154_ ) );
NOR3_X1 _1904_ ( .A1(_1153_ ), .A2(fanout_net_1 ), .A3(_1154_ ), .ZN(_0008_ ) );
OAI21_X1 _1905_ ( .A(_0943_ ), .B1(_0987_ ), .B2(_0995_ ), .ZN(_1155_ ) );
AOI21_X1 _1906_ ( .A(_0929_ ), .B1(_1155_ ), .B2(_1005_ ), .ZN(_1156_ ) );
OAI21_X1 _1907_ ( .A(_0919_ ), .B1(_1156_ ), .B2(_1010_ ), .ZN(_1157_ ) );
INV_X1 _1908_ ( .A(_1012_ ), .ZN(_1158_ ) );
AND3_X1 _1909_ ( .A1(_1157_ ), .A2(_0915_ ), .A3(_1158_ ), .ZN(_1159_ ) );
AOI21_X1 _1910_ ( .A(_0915_ ), .B1(_1157_ ), .B2(_1158_ ), .ZN(_1160_ ) );
OR3_X1 _1911_ ( .A1(_1159_ ), .A2(_1160_ ), .A3(_1116_ ), .ZN(_1161_ ) );
OAI211_X1 _1912_ ( .A(_1161_ ), .B(_1122_ ), .C1(\pc_jump [16] ), .C2(_1123_ ), .ZN(_1162_ ) );
NAND2_X1 _1913_ ( .A1(fanout_net_11 ), .A2(\mtvec [16] ), .ZN(_1163_ ) );
AOI21_X1 _1914_ ( .A(fanout_net_1 ), .B1(_1162_ ), .B2(_1163_ ), .ZN(_0009_ ) );
INV_X1 _1915_ ( .A(_1157_ ), .ZN(_1164_ ) );
NOR3_X1 _1916_ ( .A1(_1156_ ), .A2(_0919_ ), .A3(_1010_ ), .ZN(_1165_ ) );
OAI21_X1 _1917_ ( .A(_1118_ ), .B1(_1164_ ), .B2(_1165_ ), .ZN(_1166_ ) );
OAI211_X1 _1918_ ( .A(_1166_ ), .B(_1122_ ), .C1(\pc_jump [15] ), .C2(_1123_ ), .ZN(_1167_ ) );
NAND2_X1 _1919_ ( .A1(fanout_net_11 ), .A2(\mtvec [15] ), .ZN(_1168_ ) );
AOI21_X1 _1920_ ( .A(fanout_net_1 ), .B1(_1167_ ), .B2(_1168_ ), .ZN(_0010_ ) );
NAND2_X1 _1921_ ( .A1(_1155_ ), .A2(_1005_ ), .ZN(_1169_ ) );
NAND2_X1 _1922_ ( .A1(_1169_ ), .A2(_0924_ ), .ZN(_1170_ ) );
OR2_X1 _1923_ ( .A1(_0923_ ), .A2(_1008_ ), .ZN(_1171_ ) );
AND2_X1 _1924_ ( .A1(_0927_ ), .A2(_0928_ ), .ZN(_1172_ ) );
AND3_X1 _1925_ ( .A1(_1170_ ), .A2(_1171_ ), .A3(_1172_ ), .ZN(_1173_ ) );
AOI21_X1 _1926_ ( .A(_1172_ ), .B1(_1170_ ), .B2(_1171_ ), .ZN(_1174_ ) );
OR3_X1 _1927_ ( .A1(_1173_ ), .A2(_1174_ ), .A3(_1116_ ), .ZN(_1175_ ) );
OAI211_X1 _1928_ ( .A(_1175_ ), .B(_1122_ ), .C1(\pc_jump [14] ), .C2(_1123_ ), .ZN(_1176_ ) );
NAND2_X1 _1929_ ( .A1(fanout_net_11 ), .A2(\mtvec [14] ), .ZN(_1177_ ) );
AOI21_X1 _1930_ ( .A(fanout_net_1 ), .B1(_1176_ ), .B2(_1177_ ), .ZN(_0011_ ) );
XOR2_X1 _1931_ ( .A(_1169_ ), .B(_0924_ ), .Z(_1178_ ) );
MUX2_X1 _1932_ ( .A(\pc_jump [13] ), .B(_1178_ ), .S(_1117_ ), .Z(_1179_ ) );
MUX2_X1 _1933_ ( .A(\mtvec [13] ), .B(_1179_ ), .S(_1121_ ), .Z(_1180_ ) );
INV_X1 _1934_ ( .A(fanout_net_1 ), .ZN(_1181_ ) );
AND2_X1 _1935_ ( .A1(_1180_ ), .A2(_1181_ ), .ZN(_0012_ ) );
OAI21_X1 _1936_ ( .A(_0936_ ), .B1(_0987_ ), .B2(_0995_ ), .ZN(_1182_ ) );
AOI21_X1 _1937_ ( .A(_0999_ ), .B1(_0935_ ), .B2(_0997_ ), .ZN(_1183_ ) );
NAND2_X1 _1938_ ( .A1(_1182_ ), .A2(_1183_ ), .ZN(_1184_ ) );
NAND2_X1 _1939_ ( .A1(_1184_ ), .A2(_0942_ ), .ZN(_1185_ ) );
INV_X1 _1940_ ( .A(_1003_ ), .ZN(_1186_ ) );
AND3_X1 _1941_ ( .A1(_1185_ ), .A2(_0939_ ), .A3(_1186_ ), .ZN(_1187_ ) );
AOI21_X1 _1942_ ( .A(_0939_ ), .B1(_1185_ ), .B2(_1186_ ), .ZN(_1188_ ) );
OR3_X1 _1943_ ( .A1(_1187_ ), .A2(_1188_ ), .A3(_1116_ ), .ZN(_1189_ ) );
OAI211_X1 _1944_ ( .A(_1189_ ), .B(_1122_ ), .C1(\pc_jump [12] ), .C2(_1123_ ), .ZN(_1190_ ) );
NAND2_X1 _1945_ ( .A1(fanout_net_11 ), .A2(\mtvec [12] ), .ZN(_1191_ ) );
AOI21_X1 _1946_ ( .A(fanout_net_1 ), .B1(_1190_ ), .B2(_1191_ ), .ZN(_0013_ ) );
OR2_X1 _1947_ ( .A1(_1184_ ), .A2(_0942_ ), .ZN(_1192_ ) );
AND3_X1 _1948_ ( .A1(_1192_ ), .A2(_1118_ ), .A3(_1185_ ), .ZN(_1193_ ) );
AOI211_X1 _1949_ ( .A(fanout_net_11 ), .B(_1193_ ), .C1(\pc_jump [11] ), .C2(_1130_ ), .ZN(_1194_ ) );
NOR2_X1 _1950_ ( .A1(_1138_ ), .A2(\mtvec [11] ), .ZN(_1195_ ) );
NOR3_X1 _1951_ ( .A1(_1194_ ), .A2(fanout_net_1 ), .A3(_1195_ ), .ZN(_0014_ ) );
NOR2_X1 _1952_ ( .A1(_1040_ ), .A2(_1059_ ), .ZN(_1196_ ) );
INV_X1 _1953_ ( .A(_1196_ ), .ZN(_1197_ ) );
AND2_X4 _1954_ ( .A1(_1197_ ), .A2(_0908_ ), .ZN(_1198_ ) );
OAI21_X2 _1955_ ( .A(_0901_ ), .B1(_1198_ ), .B2(_1064_ ), .ZN(_1199_ ) );
NAND2_X1 _1956_ ( .A1(_0903_ ), .A2(\araddr [27] ), .ZN(_1200_ ) );
AND3_X2 _1957_ ( .A1(_1199_ ), .A2(_0899_ ), .A3(_1200_ ), .ZN(_1201_ ) );
AOI21_X1 _1958_ ( .A(_0899_ ), .B1(_1199_ ), .B2(_1200_ ), .ZN(_1202_ ) );
OR3_X2 _1959_ ( .A1(_1201_ ), .A2(_1202_ ), .A3(_1116_ ), .ZN(_1203_ ) );
OAI211_X1 _1960_ ( .A(_1203_ ), .B(_1122_ ), .C1(\pc_jump [28] ), .C2(_1123_ ), .ZN(_1204_ ) );
NAND2_X1 _1961_ ( .A1(fanout_net_11 ), .A2(\mtvec [28] ), .ZN(_1205_ ) );
AOI21_X1 _1962_ ( .A(fanout_net_1 ), .B1(_1204_ ), .B2(_1205_ ), .ZN(_0015_ ) );
NOR2_X1 _1963_ ( .A1(_0987_ ), .A2(_0995_ ), .ZN(_1206_ ) );
INV_X1 _1964_ ( .A(_0932_ ), .ZN(_1207_ ) );
NOR2_X1 _1965_ ( .A1(_1206_ ), .A2(_1207_ ), .ZN(_0040_ ) );
OR3_X1 _1966_ ( .A1(_0040_ ), .A2(_0997_ ), .A3(_0935_ ), .ZN(_0041_ ) );
OAI21_X1 _1967_ ( .A(_0935_ ), .B1(_0040_ ), .B2(_0997_ ), .ZN(_0042_ ) );
AND3_X1 _1968_ ( .A1(_0041_ ), .A2(_1117_ ), .A3(_0042_ ), .ZN(_0043_ ) );
AOI211_X1 _1969_ ( .A(fanout_net_11 ), .B(_0043_ ), .C1(\pc_jump [10] ), .C2(_1130_ ), .ZN(_0044_ ) );
NOR2_X1 _1970_ ( .A1(_1138_ ), .A2(\mtvec [10] ), .ZN(_0045_ ) );
NOR3_X1 _1971_ ( .A1(_0044_ ), .A2(fanout_net_1 ), .A3(_0045_ ), .ZN(_0016_ ) );
NOR3_X1 _1972_ ( .A1(_0987_ ), .A2(_0995_ ), .A3(_0932_ ), .ZN(_0046_ ) );
OAI21_X1 _1973_ ( .A(_1118_ ), .B1(_0040_ ), .B2(_0046_ ), .ZN(_0047_ ) );
BUF_X4 _1974_ ( .A(_1121_ ), .Z(_0048_ ) );
OAI211_X1 _1975_ ( .A(_0047_ ), .B(_0048_ ), .C1(\pc_jump [9] ), .C2(_1123_ ), .ZN(_0049_ ) );
NAND2_X1 _1976_ ( .A1(fanout_net_11 ), .A2(\mtvec [9] ), .ZN(_0050_ ) );
AOI21_X1 _1977_ ( .A(fanout_net_1 ), .B1(_0049_ ), .B2(_0050_ ), .ZN(_0017_ ) );
NOR2_X1 _1978_ ( .A1(_0972_ ), .A2(_0986_ ), .ZN(_0051_ ) );
NOR2_X1 _1979_ ( .A1(_0051_ ), .A2(_0990_ ), .ZN(_0052_ ) );
NOR2_X1 _1980_ ( .A1(_0052_ ), .A2(_0978_ ), .ZN(_0053_ ) );
OR3_X1 _1981_ ( .A1(_0053_ ), .A2(_0975_ ), .A3(_0993_ ), .ZN(_0054_ ) );
OAI21_X1 _1982_ ( .A(_0975_ ), .B1(_0053_ ), .B2(_0993_ ), .ZN(_0055_ ) );
AOI21_X1 _1983_ ( .A(_1127_ ), .B1(_0054_ ), .B2(_0055_ ), .ZN(_0056_ ) );
AOI211_X1 _1984_ ( .A(fanout_net_11 ), .B(_0056_ ), .C1(\pc_jump [8] ), .C2(_1130_ ), .ZN(_0057_ ) );
NOR2_X1 _1985_ ( .A1(_1138_ ), .A2(\mtvec [8] ), .ZN(_0058_ ) );
NOR3_X1 _1986_ ( .A1(_0057_ ), .A2(fanout_net_1 ), .A3(_0058_ ), .ZN(_0018_ ) );
NOR3_X1 _1987_ ( .A1(_0051_ ), .A2(_0977_ ), .A3(_0990_ ), .ZN(_0059_ ) );
OAI21_X1 _1988_ ( .A(_1118_ ), .B1(_0053_ ), .B2(_0059_ ), .ZN(_0060_ ) );
OAI211_X1 _1989_ ( .A(_0060_ ), .B(_0048_ ), .C1(\pc_jump [7] ), .C2(_1123_ ), .ZN(_0061_ ) );
NAND2_X1 _1990_ ( .A1(fanout_net_11 ), .A2(\mtvec [7] ), .ZN(_0062_ ) );
AOI21_X1 _1991_ ( .A(fanout_net_1 ), .B1(_0061_ ), .B2(_0062_ ), .ZN(_0019_ ) );
OR2_X1 _1992_ ( .A1(_0972_ ), .A2(_0980_ ), .ZN(_0063_ ) );
NOR2_X1 _1993_ ( .A1(_0984_ ), .A2(_0983_ ), .ZN(_0064_ ) );
AND3_X1 _1994_ ( .A1(_0063_ ), .A2(_0064_ ), .A3(_0988_ ), .ZN(_0065_ ) );
AOI21_X1 _1995_ ( .A(_0064_ ), .B1(_0063_ ), .B2(_0988_ ), .ZN(_0066_ ) );
OR3_X1 _1996_ ( .A1(_0065_ ), .A2(_0066_ ), .A3(_1116_ ), .ZN(_0067_ ) );
BUF_X4 _1997_ ( .A(_1118_ ), .Z(_0068_ ) );
OAI211_X1 _1998_ ( .A(_0067_ ), .B(_0048_ ), .C1(\pc_jump [6] ), .C2(_0068_ ), .ZN(_0069_ ) );
NAND2_X1 _1999_ ( .A1(fanout_net_11 ), .A2(\mtvec [6] ), .ZN(_0070_ ) );
AOI21_X1 _2000_ ( .A(fanout_net_1 ), .B1(_0069_ ), .B2(_0070_ ), .ZN(_0020_ ) );
XNOR2_X1 _2001_ ( .A(_0972_ ), .B(_0980_ ), .ZN(_0071_ ) );
NAND2_X1 _2002_ ( .A1(_0071_ ), .A2(_0068_ ), .ZN(_0072_ ) );
OAI211_X1 _2003_ ( .A(_0072_ ), .B(_0048_ ), .C1(\pc_jump [5] ), .C2(_0068_ ), .ZN(_0073_ ) );
NAND2_X1 _2004_ ( .A1(fanout_net_11 ), .A2(\mtvec [5] ), .ZN(_0074_ ) );
AOI21_X1 _2005_ ( .A(fanout_net_1 ), .B1(_0073_ ), .B2(_0074_ ), .ZN(_0021_ ) );
NOR2_X1 _2006_ ( .A1(_0967_ ), .A2(_0970_ ), .ZN(_0075_ ) );
OAI21_X1 _2007_ ( .A(_0968_ ), .B1(_0075_ ), .B2(_0951_ ), .ZN(_0076_ ) );
INV_X1 _2008_ ( .A(_0951_ ), .ZN(_0077_ ) );
OAI211_X1 _2009_ ( .A(_0947_ ), .B(_0077_ ), .C1(_0967_ ), .C2(_0970_ ), .ZN(_0078_ ) );
NAND3_X1 _2010_ ( .A1(_0076_ ), .A2(_1117_ ), .A3(_0078_ ), .ZN(_0079_ ) );
OAI211_X1 _2011_ ( .A(_0079_ ), .B(_1121_ ), .C1(\pc_jump [4] ), .C2(_1117_ ), .ZN(_0080_ ) );
NAND2_X1 _2012_ ( .A1(fanout_net_11 ), .A2(\mtvec [4] ), .ZN(_0081_ ) );
AOI21_X1 _2013_ ( .A(fanout_net_1 ), .B1(_0080_ ), .B2(_0081_ ), .ZN(_0022_ ) );
AND2_X1 _2014_ ( .A1(fanout_net_11 ), .A2(\mtvec [3] ), .ZN(_0082_ ) );
XOR2_X1 _2015_ ( .A(_0967_ ), .B(_0970_ ), .Z(_0083_ ) );
MUX2_X1 _2016_ ( .A(\pc_jump [3] ), .B(_0083_ ), .S(_1117_ ), .Z(_0084_ ) );
AOI21_X1 _2017_ ( .A(_0082_ ), .B1(_0084_ ), .B2(_1138_ ), .ZN(_0085_ ) );
NOR2_X1 _2018_ ( .A1(_0085_ ), .A2(fanout_net_1 ), .ZN(_0023_ ) );
AND2_X1 _2019_ ( .A1(\state [1] ), .A2(readyFromIDU ), .ZN(readyFromIDU_$_AND__B_Y ) );
AND3_X1 _2020_ ( .A1(_0080_ ), .A2(_0081_ ), .A3(readyFromIDU_$_AND__B_Y ), .ZN(_0086_ ) );
BUF_X2 _2021_ ( .A(_0946_ ), .Z(_0087_ ) );
BUF_X4 _2022_ ( .A(_0087_ ), .Z(_0088_ ) );
BUF_X2 _2023_ ( .A(_0088_ ), .Z(_0089_ ) );
INV_X1 _2024_ ( .A(readyFromIDU_$_AND__B_Y ), .ZN(_0090_ ) );
AOI211_X1 _2025_ ( .A(fanout_net_1 ), .B(_0086_ ), .C1(_0089_ ), .C2(_0090_ ), .ZN(_0024_ ) );
OAI21_X1 _2026_ ( .A(_1118_ ), .B1(_0964_ ), .B2(_0960_ ), .ZN(_0091_ ) );
NOR2_X1 _2027_ ( .A1(_0091_ ), .A2(_0965_ ), .ZN(_0092_ ) );
AOI211_X1 _2028_ ( .A(fanout_net_11 ), .B(_0092_ ), .C1(\pc_jump [2] ), .C2(_1130_ ), .ZN(_0093_ ) );
NOR2_X1 _2029_ ( .A1(_1138_ ), .A2(\mtvec [2] ), .ZN(_0094_ ) );
NOR3_X1 _2030_ ( .A1(_0093_ ), .A2(fanout_net_1 ), .A3(_0094_ ), .ZN(_0025_ ) );
AOI211_X1 _2031_ ( .A(_0082_ ), .B(_0090_ ), .C1(_0084_ ), .C2(_1121_ ), .ZN(_0095_ ) );
BUF_X4 _2032_ ( .A(_0969_ ), .Z(_0096_ ) );
BUF_X2 _2033_ ( .A(_0096_ ), .Z(_0097_ ) );
AOI211_X1 _2034_ ( .A(fanout_net_1 ), .B(_0095_ ), .C1(_0097_ ), .C2(_0090_ ), .ZN(_0026_ ) );
XNOR2_X1 _2035_ ( .A(_0963_ ), .B(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B ), .ZN(_0098_ ) );
NAND2_X1 _2036_ ( .A1(_0068_ ), .A2(_0098_ ), .ZN(_0099_ ) );
OAI211_X1 _2037_ ( .A(_0099_ ), .B(_0048_ ), .C1(\pc_jump [1] ), .C2(_0068_ ), .ZN(_0100_ ) );
NAND2_X1 _2038_ ( .A1(fanout_net_11 ), .A2(\mtvec [1] ), .ZN(_0101_ ) );
AOI21_X1 _2039_ ( .A(fanout_net_1 ), .B1(_0100_ ), .B2(_0101_ ), .ZN(_0027_ ) );
OR3_X4 _2040_ ( .A1(_1198_ ), .A2(_0901_ ), .A3(_1064_ ), .ZN(_0102_ ) );
AND3_X2 _2041_ ( .A1(_0102_ ), .A2(_1117_ ), .A3(_1199_ ), .ZN(_0103_ ) );
AOI211_X2 _2042_ ( .A(fanout_net_11 ), .B(_0103_ ), .C1(\pc_jump [27] ), .C2(_1130_ ), .ZN(_0104_ ) );
NOR2_X1 _2043_ ( .A1(_1122_ ), .A2(\mtvec [27] ), .ZN(_0105_ ) );
NOR3_X1 _2044_ ( .A1(_0104_ ), .A2(fanout_net_1 ), .A3(_0105_ ), .ZN(_0028_ ) );
NAND4_X1 _2045_ ( .A1(_1115_ ), .A2(_1122_ ), .A3(check_quest ), .A4(\pc_jump [0] ), .ZN(_0106_ ) );
NAND2_X1 _2046_ ( .A1(fanout_net_11 ), .A2(\mtvec [0] ), .ZN(_0107_ ) );
AOI21_X1 _2047_ ( .A(fanout_net_1 ), .B1(_0106_ ), .B2(_0107_ ), .ZN(_0029_ ) );
OAI21_X1 _2048_ ( .A(_0907_ ), .B1(_1040_ ), .B2(_1059_ ), .ZN(_0108_ ) );
AND3_X1 _2049_ ( .A1(_0108_ ), .A2(_0905_ ), .A3(_1062_ ), .ZN(_0109_ ) );
AOI21_X1 _2050_ ( .A(_0905_ ), .B1(_0108_ ), .B2(_1062_ ), .ZN(_0110_ ) );
OR3_X1 _2051_ ( .A1(_0109_ ), .A2(_0110_ ), .A3(_1116_ ), .ZN(_0111_ ) );
OAI211_X1 _2052_ ( .A(_0111_ ), .B(_0048_ ), .C1(\pc_jump [26] ), .C2(_0068_ ), .ZN(_0112_ ) );
NAND2_X1 _2053_ ( .A1(fanout_net_11 ), .A2(\mtvec [26] ), .ZN(_0113_ ) );
AOI21_X1 _2054_ ( .A(fanout_net_1 ), .B1(_0112_ ), .B2(_0113_ ), .ZN(_0030_ ) );
OR3_X1 _2055_ ( .A1(_1040_ ), .A2(_1059_ ), .A3(_0907_ ), .ZN(_0114_ ) );
AND3_X1 _2056_ ( .A1(_0114_ ), .A2(_1117_ ), .A3(_0108_ ), .ZN(_0115_ ) );
AOI211_X1 _2057_ ( .A(fanout_net_11 ), .B(_0115_ ), .C1(\pc_jump [25] ), .C2(_1127_ ), .ZN(_0116_ ) );
NOR2_X1 _2058_ ( .A1(_1122_ ), .A2(\mtvec [25] ), .ZN(_0117_ ) );
NOR3_X1 _2059_ ( .A1(_0116_ ), .A2(fanout_net_1 ), .A3(_0117_ ), .ZN(_0031_ ) );
NAND2_X1 _2060_ ( .A1(_1016_ ), .A2(_1039_ ), .ZN(_0118_ ) );
NOR2_X1 _2061_ ( .A1(_1048_ ), .A2(_1052_ ), .ZN(_0119_ ) );
AOI21_X1 _2062_ ( .A(_1021_ ), .B1(_0118_ ), .B2(_0119_ ), .ZN(_0120_ ) );
AND2_X1 _2063_ ( .A1(_0903_ ), .A2(\araddr [22] ), .ZN(_0121_ ) );
OR3_X1 _2064_ ( .A1(_0120_ ), .A2(_0121_ ), .A3(_1055_ ), .ZN(_0122_ ) );
NAND2_X1 _2065_ ( .A1(_0122_ ), .A2(_1023_ ), .ZN(_0123_ ) );
AND3_X1 _2066_ ( .A1(_0123_ ), .A2(_1041_ ), .A3(_1025_ ), .ZN(_0124_ ) );
AOI21_X1 _2067_ ( .A(_1025_ ), .B1(_0123_ ), .B2(_1041_ ), .ZN(_0125_ ) );
OAI21_X1 _2068_ ( .A(_1118_ ), .B1(_0124_ ), .B2(_0125_ ), .ZN(_0126_ ) );
OAI211_X1 _2069_ ( .A(_0126_ ), .B(_0048_ ), .C1(\pc_jump [24] ), .C2(_0068_ ), .ZN(_0127_ ) );
NAND2_X1 _2070_ ( .A1(fanout_net_11 ), .A2(\mtvec [24] ), .ZN(_0128_ ) );
AOI21_X1 _2071_ ( .A(fanout_net_1 ), .B1(_0127_ ), .B2(_0128_ ), .ZN(_0032_ ) );
XNOR2_X1 _2072_ ( .A(_0122_ ), .B(_1023_ ), .ZN(_0129_ ) );
NOR2_X1 _2073_ ( .A1(_0129_ ), .A2(_1127_ ), .ZN(_0130_ ) );
AOI211_X1 _2074_ ( .A(fanout_net_11 ), .B(_0130_ ), .C1(\pc_jump [23] ), .C2(_1127_ ), .ZN(_0131_ ) );
NOR2_X1 _2075_ ( .A1(_1122_ ), .A2(\mtvec [23] ), .ZN(_0132_ ) );
NOR3_X1 _2076_ ( .A1(_0131_ ), .A2(reset ), .A3(_0132_ ), .ZN(_0033_ ) );
INV_X1 _2077_ ( .A(_1018_ ), .ZN(_0133_ ) );
AOI21_X1 _2078_ ( .A(_0133_ ), .B1(_0118_ ), .B2(_0119_ ), .ZN(_0134_ ) );
AND2_X1 _2079_ ( .A1(_0903_ ), .A2(\araddr [21] ), .ZN(_0135_ ) );
OR2_X1 _2080_ ( .A1(_0134_ ), .A2(_0135_ ), .ZN(_0136_ ) );
XNOR2_X1 _2081_ ( .A(_0136_ ), .B(_1019_ ), .ZN(_0137_ ) );
NAND2_X1 _2082_ ( .A1(_0137_ ), .A2(_0068_ ), .ZN(_0138_ ) );
OAI211_X1 _2083_ ( .A(_0138_ ), .B(_0048_ ), .C1(\pc_jump [22] ), .C2(_0068_ ), .ZN(_0139_ ) );
NAND2_X1 _2084_ ( .A1(fanout_net_11 ), .A2(\mtvec [22] ), .ZN(_0140_ ) );
AOI21_X1 _2085_ ( .A(reset ), .B1(_0139_ ), .B2(_0140_ ), .ZN(_0034_ ) );
AND3_X1 _2086_ ( .A1(_0118_ ), .A2(_0133_ ), .A3(_0119_ ), .ZN(_0141_ ) );
OAI21_X1 _2087_ ( .A(_1118_ ), .B1(_0141_ ), .B2(_0134_ ), .ZN(_0142_ ) );
OAI211_X1 _2088_ ( .A(_0142_ ), .B(_0048_ ), .C1(\pc_jump [21] ), .C2(_0068_ ), .ZN(_0143_ ) );
NAND2_X1 _2089_ ( .A1(to_reset ), .A2(\mtvec [21] ), .ZN(_0144_ ) );
AOI21_X1 _2090_ ( .A(reset ), .B1(_0143_ ), .B2(_0144_ ), .ZN(_0035_ ) );
NAND2_X1 _2091_ ( .A1(to_reset ), .A2(\mtvec [31] ), .ZN(_0145_ ) );
OR3_X4 _2092_ ( .A1(_1066_ ), .A2(_1068_ ), .A3(_1071_ ), .ZN(_0146_ ) );
OAI21_X1 _2093_ ( .A(_0903_ ), .B1(\araddr [30] ), .B2(\araddr [29] ), .ZN(_0147_ ) );
XOR2_X1 _2094_ ( .A(_0903_ ), .B(\araddr [31] ), .Z(_0148_ ) );
AND3_X4 _2095_ ( .A1(_0146_ ), .A2(_0147_ ), .A3(_0148_ ), .ZN(_0149_ ) );
AOI21_X1 _2096_ ( .A(_0148_ ), .B1(_0146_ ), .B2(_0147_ ), .ZN(_0150_ ) );
NOR3_X1 _2097_ ( .A1(_0149_ ), .A2(_0150_ ), .A3(_1127_ ), .ZN(_0151_ ) );
OAI21_X1 _2098_ ( .A(_0048_ ), .B1(_1123_ ), .B2(\pc_jump [31] ), .ZN(_0152_ ) );
OAI211_X1 _2099_ ( .A(_1181_ ), .B(_0145_ ), .C1(_0151_ ), .C2(_0152_ ), .ZN(_0036_ ) );
INV_X1 _2100_ ( .A(\rid [1] ), .ZN(_0153_ ) );
NAND2_X1 _2101_ ( .A1(_0153_ ), .A2(\rid [0] ), .ZN(_0154_ ) );
NOR3_X1 _2102_ ( .A1(_0154_ ), .A2(\rid [3] ), .A3(\rid [2] ), .ZN(_0155_ ) );
NOR2_X1 _2103_ ( .A1(\rresp [1] ), .A2(\rresp [0] ), .ZN(_0156_ ) );
AND2_X1 _2104_ ( .A1(_0156_ ), .A2(rvalid ), .ZN(_0157_ ) );
AND2_X1 _2105_ ( .A1(_0155_ ), .A2(_0157_ ), .ZN(_0158_ ) );
NAND2_X1 _2106_ ( .A1(_0158_ ), .A2(rlast ), .ZN(_0159_ ) );
INV_X1 _2107_ ( .A(\tmp_offset [2] ), .ZN(_0160_ ) );
NAND3_X1 _2108_ ( .A1(_0159_ ), .A2(_1181_ ), .A3(_0160_ ), .ZN(_0161_ ) );
INV_X1 _2109_ ( .A(_0161_ ), .ZN(_0037_ ) );
NOR3_X1 _2110_ ( .A1(reset ), .A2(\state [2] ), .A3(\state [1] ), .ZN(_0038_ ) );
NOR2_X1 _2111_ ( .A1(to_reset ), .A2(stall_quest_exception_IFU ), .ZN(_0162_ ) );
AOI211_X1 _2112_ ( .A(reset ), .B(_0162_ ), .C1(to_reset ), .C2(readyFromIDU_$_AND__B_Y ), .ZN(_0039_ ) );
NOR2_X1 _2113_ ( .A1(reset ), .A2(stall_quest_fencei ), .ZN(_0163_ ) );
AND2_X1 _2114_ ( .A1(_0163_ ), .A2(\myicache.wen ), .ZN(wen_$_ANDNOT__A_Y ) );
NOR2_X1 _2115_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .ZN(_0164_ ) );
BUF_X4 _2116_ ( .A(_0164_ ), .Z(_0165_ ) );
BUF_X2 _2117_ ( .A(_0165_ ), .Z(_0166_ ) );
AND3_X1 _2118_ ( .A1(_0163_ ), .A2(_0166_ ), .A3(\myicache.wen ), .ZN(_0000_ ) );
INV_X1 _2119_ ( .A(_0163_ ), .ZN(_0167_ ) );
NAND2_X1 _2120_ ( .A1(_0089_ ), .A2(\araddr [3] ), .ZN(_0168_ ) );
INV_X1 _2121_ ( .A(\myicache.wen ), .ZN(_0169_ ) );
BUF_X4 _2122_ ( .A(_0169_ ), .Z(_0170_ ) );
NOR3_X1 _2123_ ( .A1(_0167_ ), .A2(_0168_ ), .A3(_0170_ ), .ZN(_0001_ ) );
NAND2_X1 _2124_ ( .A1(_0097_ ), .A2(\araddr [4] ), .ZN(_0171_ ) );
NOR3_X1 _2125_ ( .A1(_0167_ ), .A2(_0171_ ), .A3(_0170_ ), .ZN(_0002_ ) );
INV_X1 _2126_ ( .A(\state [0] ), .ZN(_0172_ ) );
NOR3_X1 _2127_ ( .A1(_0172_ ), .A2(reset ), .A3(stall_quest_fencei ), .ZN(arvalid ) );
INV_X1 _2128_ ( .A(\state [1] ), .ZN(_0173_ ) );
NOR2_X1 _2129_ ( .A1(_0173_ ), .A2(readyFromIDU ), .ZN(_0174_ ) );
NOR2_X1 _2130_ ( .A1(_0173_ ), .A2(to_reset ), .ZN(_0175_ ) );
INV_X1 _2131_ ( .A(_0175_ ), .ZN(_0176_ ) );
INV_X1 _2132_ ( .A(check_assert_$_DFFE_PP__Q_E_$_ANDNOT__Y_B_$_MUX__Y_A ), .ZN(_0177_ ) );
NAND2_X1 _2133_ ( .A1(_0173_ ), .A2(_0177_ ), .ZN(_0178_ ) );
AOI211_X1 _2134_ ( .A(reset ), .B(_0174_ ), .C1(_0176_ ), .C2(_0178_ ), .ZN(check_assert_$_DFFE_PP__Q_E ) );
OR2_X1 _2135_ ( .A1(_0000_ ), .A2(_0167_ ), .ZN(\myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
OAI21_X1 _2136_ ( .A(_0163_ ), .B1(_0168_ ), .B2(_0170_ ), .ZN(\myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
OAI21_X1 _2137_ ( .A(_0163_ ), .B1(_0171_ ), .B2(_0170_ ), .ZN(\myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _2138_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .ZN(_0179_ ) );
OAI21_X1 _2139_ ( .A(_0163_ ), .B1(_0179_ ), .B2(_0170_ ), .ZN(\myicache.valid[3]_$_DFFE_PP__Q_E ) );
INV_X1 _2140_ ( .A(\pc [1] ), .ZN(_0180_ ) );
OAI211_X1 _2141_ ( .A(_0180_ ), .B(tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ), .C1(_0959_ ), .C2(\tmp_offset [2] ), .ZN(_0181_ ) );
NOR2_X1 _2142_ ( .A1(_0160_ ), .A2(\pc [2] ), .ZN(_0182_ ) );
NOR2_X1 _2143_ ( .A1(_0181_ ), .A2(_0182_ ), .ZN(_0183_ ) );
AND2_X1 _2144_ ( .A1(_0158_ ), .A2(_0183_ ), .ZN(_0184_ ) );
INV_X1 _2145_ ( .A(_0184_ ), .ZN(_0185_ ) );
CLKBUF_X2 _2146_ ( .A(_0185_ ), .Z(_0186_ ) );
OR2_X1 _2147_ ( .A1(_0186_ ), .A2(\rdata [8] ), .ZN(_0187_ ) );
INV_X1 _2148_ ( .A(\state [2] ), .ZN(_0188_ ) );
BUF_X4 _2149_ ( .A(_0188_ ), .Z(_0189_ ) );
BUF_X4 _2150_ ( .A(_0185_ ), .Z(_0190_ ) );
BUF_X4 _2151_ ( .A(_0190_ ), .Z(_0191_ ) );
AOI21_X1 _2152_ ( .A(_0189_ ), .B1(_0191_ ), .B2(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_0192_ ) );
NAND2_X1 _2153_ ( .A1(_0187_ ), .A2(_0192_ ), .ZN(_0193_ ) );
AND3_X1 _2154_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .A3(\myicache.data[6][8] ), .ZN(_0194_ ) );
AND3_X1 _2155_ ( .A1(_0088_ ), .A2(\araddr [3] ), .A3(\myicache.data[2][8] ), .ZN(_0195_ ) );
AOI211_X1 _2156_ ( .A(_0194_ ), .B(_0195_ ), .C1(\myicache.data[0][8] ), .C2(_0166_ ), .ZN(_0196_ ) );
NAND2_X1 _2157_ ( .A1(_0169_ ), .A2(\pc [2] ), .ZN(_0197_ ) );
BUF_X4 _2158_ ( .A(_0197_ ), .Z(_0198_ ) );
BUF_X2 _2159_ ( .A(_0198_ ), .Z(_0199_ ) );
NAND2_X1 _2160_ ( .A1(\tmp_offset [2] ), .A2(\myicache.wen ), .ZN(_0200_ ) );
BUF_X4 _2161_ ( .A(_0200_ ), .Z(_0201_ ) );
BUF_X4 _2162_ ( .A(_0201_ ), .Z(_0202_ ) );
NAND3_X1 _2163_ ( .A1(_0097_ ), .A2(\araddr [4] ), .A3(\myicache.data[4][8] ), .ZN(_0203_ ) );
NAND4_X1 _2164_ ( .A1(_0196_ ), .A2(_0199_ ), .A3(_0202_ ), .A4(_0203_ ), .ZN(_0204_ ) );
NOR2_X2 _2165_ ( .A1(\state [2] ), .A2(\state [1] ), .ZN(_0205_ ) );
BUF_X4 _2166_ ( .A(_0205_ ), .Z(_0206_ ) );
BUF_X4 _2167_ ( .A(_0087_ ), .Z(_0207_ ) );
BUF_X4 _2168_ ( .A(_0207_ ), .Z(_0208_ ) );
NAND3_X1 _2169_ ( .A1(_0208_ ), .A2(\araddr [3] ), .A3(\myicache.data[3][8] ), .ZN(_0209_ ) );
NAND3_X1 _2170_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .A3(\myicache.data[7][8] ), .ZN(_0210_ ) );
AND2_X1 _2171_ ( .A1(_0209_ ), .A2(_0210_ ), .ZN(_0211_ ) );
NAND2_X1 _2172_ ( .A1(_0197_ ), .A2(_0200_ ), .ZN(_0212_ ) );
BUF_X2 _2173_ ( .A(_0212_ ), .Z(_0213_ ) );
BUF_X4 _2174_ ( .A(_0969_ ), .Z(_0214_ ) );
BUF_X4 _2175_ ( .A(_0214_ ), .Z(_0215_ ) );
NAND3_X1 _2176_ ( .A1(_0215_ ), .A2(\araddr [4] ), .A3(\myicache.data[5][8] ), .ZN(_0216_ ) );
BUF_X4 _2177_ ( .A(_0096_ ), .Z(_0217_ ) );
NAND3_X1 _2178_ ( .A1(_0217_ ), .A2(_0089_ ), .A3(\myicache.data[1][8] ), .ZN(_0218_ ) );
NAND4_X1 _2179_ ( .A1(_0211_ ), .A2(_0213_ ), .A3(_0216_ ), .A4(_0218_ ), .ZN(_0219_ ) );
NAND3_X1 _2180_ ( .A1(_0204_ ), .A2(_0206_ ), .A3(_0219_ ), .ZN(_0220_ ) );
NAND2_X1 _2181_ ( .A1(_0193_ ), .A2(_0220_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ) );
OR2_X1 _2182_ ( .A1(_0186_ ), .A2(\rdata [31] ), .ZN(_0221_ ) );
AOI21_X1 _2183_ ( .A(_0189_ ), .B1(_0191_ ), .B2(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_0222_ ) );
NAND2_X1 _2184_ ( .A1(_0221_ ), .A2(_0222_ ), .ZN(_0223_ ) );
AND3_X1 _2185_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .A3(\myicache.data[6][31] ), .ZN(_0224_ ) );
AND3_X1 _2186_ ( .A1(_0088_ ), .A2(\araddr [3] ), .A3(\myicache.data[2][31] ), .ZN(_0225_ ) );
AOI211_X1 _2187_ ( .A(_0224_ ), .B(_0225_ ), .C1(\myicache.data[0][31] ), .C2(_0166_ ), .ZN(_0226_ ) );
NAND3_X1 _2188_ ( .A1(_0097_ ), .A2(\araddr [4] ), .A3(\myicache.data[4][31] ), .ZN(_0227_ ) );
NAND4_X1 _2189_ ( .A1(_0226_ ), .A2(_0199_ ), .A3(_0202_ ), .A4(_0227_ ), .ZN(_0228_ ) );
BUF_X4 _2190_ ( .A(_0207_ ), .Z(_0229_ ) );
NAND3_X1 _2191_ ( .A1(_0229_ ), .A2(\araddr [3] ), .A3(\myicache.data[3][31] ), .ZN(_0230_ ) );
NAND3_X1 _2192_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .A3(\myicache.data[7][31] ), .ZN(_0231_ ) );
AND2_X1 _2193_ ( .A1(_0230_ ), .A2(_0231_ ), .ZN(_0232_ ) );
NAND3_X1 _2194_ ( .A1(_0215_ ), .A2(\araddr [4] ), .A3(\myicache.data[5][31] ), .ZN(_0233_ ) );
BUF_X4 _2195_ ( .A(_0096_ ), .Z(_0234_ ) );
NAND3_X1 _2196_ ( .A1(_0234_ ), .A2(_0089_ ), .A3(\myicache.data[1][31] ), .ZN(_0235_ ) );
NAND4_X1 _2197_ ( .A1(_0232_ ), .A2(_0213_ ), .A3(_0233_ ), .A4(_0235_ ), .ZN(_0236_ ) );
NAND3_X1 _2198_ ( .A1(_0228_ ), .A2(_0206_ ), .A3(_0236_ ), .ZN(_0237_ ) );
NAND2_X1 _2199_ ( .A1(_0223_ ), .A2(_0237_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ) );
AND3_X1 _2200_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .A3(\myicache.data[6][30] ), .ZN(_0238_ ) );
AND3_X1 _2201_ ( .A1(_0207_ ), .A2(\araddr [3] ), .A3(\myicache.data[2][30] ), .ZN(_0239_ ) );
BUF_X4 _2202_ ( .A(_0165_ ), .Z(_0240_ ) );
AOI211_X1 _2203_ ( .A(_0238_ ), .B(_0239_ ), .C1(\myicache.data[0][30] ), .C2(_0240_ ), .ZN(_0241_ ) );
BUF_X4 _2204_ ( .A(_0096_ ), .Z(_0242_ ) );
NAND3_X1 _2205_ ( .A1(_0242_ ), .A2(\araddr [4] ), .A3(\myicache.data[4][30] ), .ZN(_0243_ ) );
NAND4_X1 _2206_ ( .A1(_0241_ ), .A2(_0198_ ), .A3(_0201_ ), .A4(_0243_ ), .ZN(_0244_ ) );
NAND3_X1 _2207_ ( .A1(_0088_ ), .A2(\araddr [3] ), .A3(\myicache.data[3][30] ), .ZN(_0245_ ) );
NAND3_X1 _2208_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .A3(\myicache.data[7][30] ), .ZN(_0246_ ) );
AND2_X1 _2209_ ( .A1(_0245_ ), .A2(_0246_ ), .ZN(_0247_ ) );
BUF_X2 _2210_ ( .A(_0212_ ), .Z(_0248_ ) );
NAND3_X1 _2211_ ( .A1(_0242_ ), .A2(\araddr [4] ), .A3(\myicache.data[5][30] ), .ZN(_0249_ ) );
NAND3_X1 _2212_ ( .A1(_0242_ ), .A2(_0208_ ), .A3(\myicache.data[1][30] ), .ZN(_0250_ ) );
NAND4_X1 _2213_ ( .A1(_0247_ ), .A2(_0248_ ), .A3(_0249_ ), .A4(_0250_ ), .ZN(_0251_ ) );
NAND3_X1 _2214_ ( .A1(_0244_ ), .A2(_0205_ ), .A3(_0251_ ), .ZN(_0252_ ) );
NOR2_X1 _2215_ ( .A1(_0191_ ), .A2(\rdata [30] ), .ZN(_0253_ ) );
OAI21_X1 _2216_ ( .A(\state [2] ), .B1(_0184_ ), .B2(_0933_ ), .ZN(_0254_ ) );
OAI21_X1 _2217_ ( .A(_0252_ ), .B1(_0253_ ), .B2(_0254_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ) );
OR2_X1 _2218_ ( .A1(_0186_ ), .A2(\rdata [21] ), .ZN(_0255_ ) );
AOI21_X1 _2219_ ( .A(_0189_ ), .B1(_0191_ ), .B2(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0256_ ) );
NAND2_X1 _2220_ ( .A1(_0255_ ), .A2(_0256_ ), .ZN(_0257_ ) );
AND3_X1 _2221_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .A3(\myicache.data[6][21] ), .ZN(_0258_ ) );
AND3_X1 _2222_ ( .A1(_0088_ ), .A2(\araddr [3] ), .A3(\myicache.data[2][21] ), .ZN(_0259_ ) );
AOI211_X1 _2223_ ( .A(_0258_ ), .B(_0259_ ), .C1(\myicache.data[0][21] ), .C2(_0166_ ), .ZN(_0260_ ) );
NAND3_X1 _2224_ ( .A1(_0097_ ), .A2(\araddr [4] ), .A3(\myicache.data[4][21] ), .ZN(_0261_ ) );
NAND4_X1 _2225_ ( .A1(_0260_ ), .A2(_0199_ ), .A3(_0202_ ), .A4(_0261_ ), .ZN(_0262_ ) );
NAND3_X1 _2226_ ( .A1(_0229_ ), .A2(\araddr [3] ), .A3(\myicache.data[3][21] ), .ZN(_0263_ ) );
NAND3_X1 _2227_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .A3(\myicache.data[7][21] ), .ZN(_0264_ ) );
AND2_X1 _2228_ ( .A1(_0263_ ), .A2(_0264_ ), .ZN(_0265_ ) );
NAND3_X1 _2229_ ( .A1(_0215_ ), .A2(\araddr [4] ), .A3(\myicache.data[5][21] ), .ZN(_0266_ ) );
NAND3_X1 _2230_ ( .A1(_0234_ ), .A2(_0089_ ), .A3(\myicache.data[1][21] ), .ZN(_0267_ ) );
NAND4_X1 _2231_ ( .A1(_0265_ ), .A2(_0213_ ), .A3(_0266_ ), .A4(_0267_ ), .ZN(_0268_ ) );
NAND3_X1 _2232_ ( .A1(_0262_ ), .A2(_0206_ ), .A3(_0268_ ), .ZN(_0269_ ) );
NAND2_X1 _2233_ ( .A1(_0257_ ), .A2(_0269_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ) );
OR2_X1 _2234_ ( .A1(_0186_ ), .A2(\rdata [20] ), .ZN(_0270_ ) );
AOI21_X1 _2235_ ( .A(_0189_ ), .B1(_0191_ ), .B2(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0271_ ) );
NAND2_X1 _2236_ ( .A1(_0270_ ), .A2(_0271_ ), .ZN(_0272_ ) );
AND3_X1 _2237_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .A3(\myicache.data[6][20] ), .ZN(_0273_ ) );
CLKBUF_X2 _2238_ ( .A(_0087_ ), .Z(_0274_ ) );
AND3_X1 _2239_ ( .A1(_0274_ ), .A2(\araddr [3] ), .A3(\myicache.data[2][20] ), .ZN(_0275_ ) );
AOI211_X1 _2240_ ( .A(_0273_ ), .B(_0275_ ), .C1(\myicache.data[0][20] ), .C2(_0166_ ), .ZN(_0276_ ) );
NAND3_X1 _2241_ ( .A1(_0097_ ), .A2(\araddr [4] ), .A3(\myicache.data[4][20] ), .ZN(_0277_ ) );
NAND4_X1 _2242_ ( .A1(_0276_ ), .A2(_0199_ ), .A3(_0202_ ), .A4(_0277_ ), .ZN(_0278_ ) );
NAND3_X1 _2243_ ( .A1(_0229_ ), .A2(\araddr [3] ), .A3(\myicache.data[3][20] ), .ZN(_0279_ ) );
NAND3_X1 _2244_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .A3(\myicache.data[7][20] ), .ZN(_0280_ ) );
AND2_X1 _2245_ ( .A1(_0279_ ), .A2(_0280_ ), .ZN(_0281_ ) );
BUF_X4 _2246_ ( .A(_0248_ ), .Z(_0282_ ) );
NAND3_X1 _2247_ ( .A1(_0215_ ), .A2(\araddr [4] ), .A3(\myicache.data[5][20] ), .ZN(_0283_ ) );
NAND3_X1 _2248_ ( .A1(_0234_ ), .A2(_0089_ ), .A3(\myicache.data[1][20] ), .ZN(_0284_ ) );
NAND4_X1 _2249_ ( .A1(_0281_ ), .A2(_0282_ ), .A3(_0283_ ), .A4(_0284_ ), .ZN(_0285_ ) );
NAND3_X1 _2250_ ( .A1(_0278_ ), .A2(_0206_ ), .A3(_0285_ ), .ZN(_0286_ ) );
NAND2_X1 _2251_ ( .A1(_0272_ ), .A2(_0286_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ) );
BUF_X4 _2252_ ( .A(_0188_ ), .Z(_0287_ ) );
NOR2_X1 _2253_ ( .A1(_0190_ ), .A2(\rdata [19] ), .ZN(_0288_ ) );
BUF_X4 _2254_ ( .A(_0185_ ), .Z(_0289_ ) );
AOI211_X1 _2255_ ( .A(_0287_ ), .B(_0288_ ), .C1(pc_$_SDFFE_PP0P__Q_10_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ), .C2(_0289_ ), .ZN(_0290_ ) );
INV_X1 _2256_ ( .A(_0205_ ), .ZN(_0291_ ) );
AND3_X1 _2257_ ( .A1(\araddr [3] ), .A2(\araddr [4] ), .A3(\myicache.data[6][19] ), .ZN(_0292_ ) );
AND3_X1 _2258_ ( .A1(_0087_ ), .A2(\araddr [3] ), .A3(\myicache.data[2][19] ), .ZN(_0293_ ) );
AOI211_X1 _2259_ ( .A(_0292_ ), .B(_0293_ ), .C1(\myicache.data[0][19] ), .C2(_0165_ ), .ZN(_0294_ ) );
NAND3_X1 _2260_ ( .A1(_0096_ ), .A2(\araddr [4] ), .A3(\myicache.data[4][19] ), .ZN(_0295_ ) );
AND4_X1 _2261_ ( .A1(_0198_ ), .A2(_0294_ ), .A3(_0201_ ), .A4(_0295_ ), .ZN(_0296_ ) );
NAND3_X1 _2262_ ( .A1(_0214_ ), .A2(\araddr [4] ), .A3(\myicache.data[5][19] ), .ZN(_0297_ ) );
AND2_X1 _2263_ ( .A1(_0248_ ), .A2(_0297_ ), .ZN(_0298_ ) );
AND3_X1 _2264_ ( .A1(\araddr [3] ), .A2(fanout_net_7 ), .A3(\myicache.data[7][19] ), .ZN(_0299_ ) );
AND3_X1 _2265_ ( .A1(_0207_ ), .A2(\araddr [3] ), .A3(\myicache.data[3][19] ), .ZN(_0300_ ) );
AOI211_X1 _2266_ ( .A(_0299_ ), .B(_0300_ ), .C1(\myicache.data[1][19] ), .C2(_0165_ ), .ZN(_0301_ ) );
AOI211_X1 _2267_ ( .A(_0291_ ), .B(_0296_ ), .C1(_0298_ ), .C2(_0301_ ), .ZN(_0302_ ) );
OR2_X1 _2268_ ( .A1(_0290_ ), .A2(_0302_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ) );
OR2_X1 _2269_ ( .A1(_0186_ ), .A2(\rdata [18] ), .ZN(_0303_ ) );
AOI21_X1 _2270_ ( .A(_0189_ ), .B1(_0191_ ), .B2(pc_$_SDFFE_PP0P__Q_12_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0304_ ) );
NAND2_X1 _2271_ ( .A1(_0303_ ), .A2(_0304_ ), .ZN(_0305_ ) );
AND3_X1 _2272_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[6][18] ), .ZN(_0306_ ) );
AND3_X1 _2273_ ( .A1(_0274_ ), .A2(fanout_net_3 ), .A3(\myicache.data[2][18] ), .ZN(_0307_ ) );
AOI211_X1 _2274_ ( .A(_0306_ ), .B(_0307_ ), .C1(\myicache.data[0][18] ), .C2(_0166_ ), .ZN(_0308_ ) );
NAND3_X1 _2275_ ( .A1(_0097_ ), .A2(fanout_net_7 ), .A3(\myicache.data[4][18] ), .ZN(_0309_ ) );
NAND4_X1 _2276_ ( .A1(_0308_ ), .A2(_0199_ ), .A3(_0202_ ), .A4(_0309_ ), .ZN(_0310_ ) );
NAND3_X1 _2277_ ( .A1(_0229_ ), .A2(fanout_net_3 ), .A3(\myicache.data[3][18] ), .ZN(_0311_ ) );
NAND3_X1 _2278_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[7][18] ), .ZN(_0312_ ) );
AND2_X1 _2279_ ( .A1(_0311_ ), .A2(_0312_ ), .ZN(_0313_ ) );
BUF_X4 _2280_ ( .A(_0214_ ), .Z(_0314_ ) );
NAND3_X1 _2281_ ( .A1(_0314_ ), .A2(fanout_net_7 ), .A3(\myicache.data[5][18] ), .ZN(_0315_ ) );
NAND3_X1 _2282_ ( .A1(_0234_ ), .A2(_0089_ ), .A3(\myicache.data[1][18] ), .ZN(_0316_ ) );
NAND4_X1 _2283_ ( .A1(_0313_ ), .A2(_0282_ ), .A3(_0315_ ), .A4(_0316_ ), .ZN(_0317_ ) );
NAND3_X1 _2284_ ( .A1(_0310_ ), .A2(_0206_ ), .A3(_0317_ ), .ZN(_0318_ ) );
NAND2_X1 _2285_ ( .A1(_0305_ ), .A2(_0318_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ) );
NOR2_X1 _2286_ ( .A1(_0190_ ), .A2(\rdata [17] ), .ZN(_0319_ ) );
AOI211_X1 _2287_ ( .A(_0287_ ), .B(_0319_ ), .C1(pc_$_SDFFE_PP0P__Q_12_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ORNOT__Y_B_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ), .C2(_0289_ ), .ZN(_0320_ ) );
AND3_X1 _2288_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[6][17] ), .ZN(_0321_ ) );
AND3_X1 _2289_ ( .A1(_0087_ ), .A2(fanout_net_3 ), .A3(\myicache.data[2][17] ), .ZN(_0322_ ) );
AOI211_X1 _2290_ ( .A(_0321_ ), .B(_0322_ ), .C1(\myicache.data[0][17] ), .C2(_0164_ ), .ZN(_0323_ ) );
NAND3_X1 _2291_ ( .A1(_0096_ ), .A2(fanout_net_7 ), .A3(\myicache.data[4][17] ), .ZN(_0324_ ) );
AND4_X1 _2292_ ( .A1(_0197_ ), .A2(_0323_ ), .A3(_0200_ ), .A4(_0324_ ), .ZN(_0325_ ) );
NAND3_X1 _2293_ ( .A1(_0214_ ), .A2(fanout_net_7 ), .A3(\myicache.data[5][17] ), .ZN(_0326_ ) );
AND2_X1 _2294_ ( .A1(_0248_ ), .A2(_0326_ ), .ZN(_0327_ ) );
AND3_X1 _2295_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[7][17] ), .ZN(_0328_ ) );
AND3_X1 _2296_ ( .A1(_0207_ ), .A2(fanout_net_3 ), .A3(\myicache.data[3][17] ), .ZN(_0329_ ) );
AOI211_X1 _2297_ ( .A(_0328_ ), .B(_0329_ ), .C1(\myicache.data[1][17] ), .C2(_0165_ ), .ZN(_0330_ ) );
AOI211_X1 _2298_ ( .A(_0291_ ), .B(_0325_ ), .C1(_0327_ ), .C2(_0330_ ), .ZN(_0331_ ) );
OR2_X1 _2299_ ( .A1(_0320_ ), .A2(_0331_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ) );
NOR2_X1 _2300_ ( .A1(_0190_ ), .A2(\rdata [16] ), .ZN(_0332_ ) );
AOI211_X1 _2301_ ( .A(_0287_ ), .B(_0332_ ), .C1(pc_$_SDFFE_PP0P__Q_14_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .C2(_0289_ ), .ZN(_0333_ ) );
AND3_X1 _2302_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[6][16] ), .ZN(_0334_ ) );
AND3_X1 _2303_ ( .A1(_0087_ ), .A2(fanout_net_3 ), .A3(\myicache.data[2][16] ), .ZN(_0335_ ) );
AOI211_X1 _2304_ ( .A(_0334_ ), .B(_0335_ ), .C1(\myicache.data[0][16] ), .C2(_0164_ ), .ZN(_0336_ ) );
NAND3_X1 _2305_ ( .A1(_0096_ ), .A2(fanout_net_7 ), .A3(\myicache.data[4][16] ), .ZN(_0337_ ) );
AND4_X1 _2306_ ( .A1(_0197_ ), .A2(_0336_ ), .A3(_0200_ ), .A4(_0337_ ), .ZN(_0338_ ) );
NAND3_X1 _2307_ ( .A1(_0214_ ), .A2(fanout_net_7 ), .A3(\myicache.data[5][16] ), .ZN(_0339_ ) );
AND2_X1 _2308_ ( .A1(_0248_ ), .A2(_0339_ ), .ZN(_0340_ ) );
AND3_X1 _2309_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[7][16] ), .ZN(_0341_ ) );
AND3_X1 _2310_ ( .A1(_0207_ ), .A2(fanout_net_3 ), .A3(\myicache.data[3][16] ), .ZN(_0342_ ) );
AOI211_X1 _2311_ ( .A(_0341_ ), .B(_0342_ ), .C1(\myicache.data[1][16] ), .C2(_0165_ ), .ZN(_0343_ ) );
AOI211_X1 _2312_ ( .A(_0291_ ), .B(_0338_ ), .C1(_0340_ ), .C2(_0343_ ), .ZN(_0344_ ) );
OR2_X1 _2313_ ( .A1(_0333_ ), .A2(_0344_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ) );
OR2_X1 _2314_ ( .A1(_0186_ ), .A2(\rdata [15] ), .ZN(_0345_ ) );
AOI21_X1 _2315_ ( .A(_0189_ ), .B1(_0191_ ), .B2(pc_$_SDFFE_PP0P__Q_14_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0346_ ) );
NAND2_X1 _2316_ ( .A1(_0345_ ), .A2(_0346_ ), .ZN(_0347_ ) );
AND3_X1 _2317_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[6][15] ), .ZN(_0348_ ) );
AND3_X1 _2318_ ( .A1(_0274_ ), .A2(fanout_net_3 ), .A3(\myicache.data[2][15] ), .ZN(_0349_ ) );
AOI211_X1 _2319_ ( .A(_0348_ ), .B(_0349_ ), .C1(\myicache.data[0][15] ), .C2(_0166_ ), .ZN(_0350_ ) );
NAND3_X1 _2320_ ( .A1(_0097_ ), .A2(fanout_net_7 ), .A3(\myicache.data[4][15] ), .ZN(_0351_ ) );
NAND4_X1 _2321_ ( .A1(_0350_ ), .A2(_0199_ ), .A3(_0202_ ), .A4(_0351_ ), .ZN(_0352_ ) );
NAND3_X1 _2322_ ( .A1(_0229_ ), .A2(fanout_net_3 ), .A3(\myicache.data[3][15] ), .ZN(_0353_ ) );
NAND3_X1 _2323_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[7][15] ), .ZN(_0354_ ) );
AND2_X1 _2324_ ( .A1(_0353_ ), .A2(_0354_ ), .ZN(_0355_ ) );
NAND3_X1 _2325_ ( .A1(_0314_ ), .A2(fanout_net_7 ), .A3(\myicache.data[5][15] ), .ZN(_0356_ ) );
NAND3_X1 _2326_ ( .A1(_0234_ ), .A2(_0089_ ), .A3(\myicache.data[1][15] ), .ZN(_0357_ ) );
NAND4_X1 _2327_ ( .A1(_0355_ ), .A2(_0282_ ), .A3(_0356_ ), .A4(_0357_ ), .ZN(_0358_ ) );
NAND3_X1 _2328_ ( .A1(_0352_ ), .A2(_0206_ ), .A3(_0358_ ), .ZN(_0359_ ) );
NAND2_X1 _2329_ ( .A1(_0347_ ), .A2(_0359_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ) );
NOR2_X1 _2330_ ( .A1(_0185_ ), .A2(\rdata [14] ), .ZN(_0360_ ) );
AOI211_X1 _2331_ ( .A(_0287_ ), .B(_0360_ ), .C1(pc_$_SDFFE_PP0P__Q_16_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .C2(_0289_ ), .ZN(_0361_ ) );
AND3_X1 _2332_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[6][14] ), .ZN(_0362_ ) );
AND3_X1 _2333_ ( .A1(_0087_ ), .A2(fanout_net_3 ), .A3(\myicache.data[2][14] ), .ZN(_0363_ ) );
AOI211_X1 _2334_ ( .A(_0362_ ), .B(_0363_ ), .C1(\myicache.data[0][14] ), .C2(_0164_ ), .ZN(_0364_ ) );
NAND3_X1 _2335_ ( .A1(_0096_ ), .A2(fanout_net_7 ), .A3(\myicache.data[4][14] ), .ZN(_0365_ ) );
AND4_X1 _2336_ ( .A1(_0197_ ), .A2(_0364_ ), .A3(_0200_ ), .A4(_0365_ ), .ZN(_0366_ ) );
NAND3_X1 _2337_ ( .A1(_0214_ ), .A2(fanout_net_7 ), .A3(\myicache.data[5][14] ), .ZN(_0367_ ) );
AND2_X1 _2338_ ( .A1(_0248_ ), .A2(_0367_ ), .ZN(_0368_ ) );
AND3_X1 _2339_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[7][14] ), .ZN(_0369_ ) );
AND3_X1 _2340_ ( .A1(_0207_ ), .A2(fanout_net_3 ), .A3(\myicache.data[3][14] ), .ZN(_0370_ ) );
AOI211_X1 _2341_ ( .A(_0369_ ), .B(_0370_ ), .C1(\myicache.data[1][14] ), .C2(_0165_ ), .ZN(_0371_ ) );
AOI211_X1 _2342_ ( .A(_0291_ ), .B(_0366_ ), .C1(_0368_ ), .C2(_0371_ ), .ZN(_0372_ ) );
OR2_X1 _2343_ ( .A1(_0361_ ), .A2(_0372_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ) );
NOR2_X1 _2344_ ( .A1(_0185_ ), .A2(\rdata [13] ), .ZN(_0373_ ) );
AOI211_X1 _2345_ ( .A(_0188_ ), .B(_0373_ ), .C1(pc_$_SDFFE_PP0P__Q_16_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ), .C2(_0186_ ), .ZN(_0374_ ) );
AND3_X1 _2346_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[6][13] ), .ZN(_0375_ ) );
AND3_X1 _2347_ ( .A1(_0946_ ), .A2(fanout_net_3 ), .A3(\myicache.data[2][13] ), .ZN(_0376_ ) );
AOI211_X1 _2348_ ( .A(_0375_ ), .B(_0376_ ), .C1(\myicache.data[0][13] ), .C2(_0164_ ), .ZN(_0377_ ) );
NAND3_X1 _2349_ ( .A1(_0096_ ), .A2(fanout_net_7 ), .A3(\myicache.data[4][13] ), .ZN(_0378_ ) );
AND4_X1 _2350_ ( .A1(_0197_ ), .A2(_0377_ ), .A3(_0200_ ), .A4(_0378_ ), .ZN(_0379_ ) );
NAND3_X1 _2351_ ( .A1(_0214_ ), .A2(fanout_net_7 ), .A3(\myicache.data[5][13] ), .ZN(_0380_ ) );
AND2_X1 _2352_ ( .A1(_0248_ ), .A2(_0380_ ), .ZN(_0381_ ) );
AND3_X1 _2353_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[7][13] ), .ZN(_0382_ ) );
AND3_X1 _2354_ ( .A1(_0087_ ), .A2(fanout_net_3 ), .A3(\myicache.data[3][13] ), .ZN(_0383_ ) );
AOI211_X1 _2355_ ( .A(_0382_ ), .B(_0383_ ), .C1(\myicache.data[1][13] ), .C2(_0165_ ), .ZN(_0384_ ) );
AOI211_X1 _2356_ ( .A(_0291_ ), .B(_0379_ ), .C1(_0381_ ), .C2(_0384_ ), .ZN(_0385_ ) );
OR2_X1 _2357_ ( .A1(_0374_ ), .A2(_0385_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ) );
OR2_X1 _2358_ ( .A1(_0186_ ), .A2(\rdata [12] ), .ZN(_0386_ ) );
AOI21_X1 _2359_ ( .A(_0189_ ), .B1(_0191_ ), .B2(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0387_ ) );
NAND2_X1 _2360_ ( .A1(_0386_ ), .A2(_0387_ ), .ZN(_0388_ ) );
AND3_X1 _2361_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[6][12] ), .ZN(_0389_ ) );
AND3_X1 _2362_ ( .A1(_0274_ ), .A2(fanout_net_3 ), .A3(\myicache.data[2][12] ), .ZN(_0390_ ) );
BUF_X4 _2363_ ( .A(_0165_ ), .Z(_0391_ ) );
AOI211_X1 _2364_ ( .A(_0389_ ), .B(_0390_ ), .C1(\myicache.data[0][12] ), .C2(_0391_ ), .ZN(_0392_ ) );
NAND3_X1 _2365_ ( .A1(_0097_ ), .A2(fanout_net_7 ), .A3(\myicache.data[4][12] ), .ZN(_0393_ ) );
NAND4_X1 _2366_ ( .A1(_0392_ ), .A2(_0199_ ), .A3(_0202_ ), .A4(_0393_ ), .ZN(_0394_ ) );
NAND3_X1 _2367_ ( .A1(_0229_ ), .A2(fanout_net_3 ), .A3(\myicache.data[3][12] ), .ZN(_0395_ ) );
NAND3_X1 _2368_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[7][12] ), .ZN(_0396_ ) );
AND2_X1 _2369_ ( .A1(_0395_ ), .A2(_0396_ ), .ZN(_0397_ ) );
NAND3_X1 _2370_ ( .A1(_0314_ ), .A2(fanout_net_7 ), .A3(\myicache.data[5][12] ), .ZN(_0398_ ) );
NAND3_X1 _2371_ ( .A1(_0234_ ), .A2(_0089_ ), .A3(\myicache.data[1][12] ), .ZN(_0399_ ) );
NAND4_X1 _2372_ ( .A1(_0397_ ), .A2(_0282_ ), .A3(_0398_ ), .A4(_0399_ ), .ZN(_0400_ ) );
NAND3_X1 _2373_ ( .A1(_0394_ ), .A2(_0206_ ), .A3(_0400_ ), .ZN(_0401_ ) );
NAND2_X1 _2374_ ( .A1(_0388_ ), .A2(_0401_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ) );
NOR2_X1 _2375_ ( .A1(_0185_ ), .A2(\rdata [29] ), .ZN(_0402_ ) );
AOI211_X1 _2376_ ( .A(_0188_ ), .B(_0402_ ), .C1(pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_0186_ ), .ZN(_0403_ ) );
AND3_X1 _2377_ ( .A1(fanout_net_3 ), .A2(fanout_net_7 ), .A3(\myicache.data[6][29] ), .ZN(_0404_ ) );
AND3_X1 _2378_ ( .A1(_0946_ ), .A2(fanout_net_3 ), .A3(\myicache.data[2][29] ), .ZN(_0405_ ) );
AOI211_X1 _2379_ ( .A(_0404_ ), .B(_0405_ ), .C1(\myicache.data[0][29] ), .C2(_0164_ ), .ZN(_0406_ ) );
NAND3_X1 _2380_ ( .A1(_0969_ ), .A2(fanout_net_8 ), .A3(\myicache.data[4][29] ), .ZN(_0407_ ) );
AND4_X1 _2381_ ( .A1(_0197_ ), .A2(_0406_ ), .A3(_0200_ ), .A4(_0407_ ), .ZN(_0408_ ) );
NAND3_X1 _2382_ ( .A1(_0214_ ), .A2(fanout_net_8 ), .A3(\myicache.data[5][29] ), .ZN(_0409_ ) );
AND2_X1 _2383_ ( .A1(_0248_ ), .A2(_0409_ ), .ZN(_0410_ ) );
AND3_X1 _2384_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[7][29] ), .ZN(_0411_ ) );
AND3_X1 _2385_ ( .A1(_0087_ ), .A2(fanout_net_4 ), .A3(\myicache.data[3][29] ), .ZN(_0412_ ) );
AOI211_X1 _2386_ ( .A(_0411_ ), .B(_0412_ ), .C1(\myicache.data[1][29] ), .C2(_0165_ ), .ZN(_0413_ ) );
AOI211_X1 _2387_ ( .A(_0291_ ), .B(_0408_ ), .C1(_0410_ ), .C2(_0413_ ), .ZN(_0414_ ) );
OR2_X1 _2388_ ( .A1(_0403_ ), .A2(_0414_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ) );
OR2_X1 _2389_ ( .A1(_0186_ ), .A2(\rdata [11] ), .ZN(_0415_ ) );
BUF_X4 _2390_ ( .A(_0190_ ), .Z(_0416_ ) );
AOI21_X1 _2391_ ( .A(_0189_ ), .B1(_0416_ ), .B2(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_0417_ ) );
NAND2_X1 _2392_ ( .A1(_0415_ ), .A2(_0417_ ), .ZN(_0418_ ) );
AND3_X1 _2393_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[6][11] ), .ZN(_0419_ ) );
AND3_X1 _2394_ ( .A1(_0274_ ), .A2(fanout_net_4 ), .A3(\myicache.data[2][11] ), .ZN(_0420_ ) );
AOI211_X1 _2395_ ( .A(_0419_ ), .B(_0420_ ), .C1(\myicache.data[0][11] ), .C2(_0391_ ), .ZN(_0421_ ) );
BUF_X4 _2396_ ( .A(_0214_ ), .Z(_0422_ ) );
NAND3_X1 _2397_ ( .A1(_0422_ ), .A2(fanout_net_8 ), .A3(\myicache.data[4][11] ), .ZN(_0423_ ) );
NAND4_X1 _2398_ ( .A1(_0421_ ), .A2(_0199_ ), .A3(_0202_ ), .A4(_0423_ ), .ZN(_0424_ ) );
NAND3_X1 _2399_ ( .A1(_0229_ ), .A2(fanout_net_4 ), .A3(\myicache.data[3][11] ), .ZN(_0425_ ) );
NAND3_X1 _2400_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[7][11] ), .ZN(_0426_ ) );
AND2_X1 _2401_ ( .A1(_0425_ ), .A2(_0426_ ), .ZN(_0427_ ) );
NAND3_X1 _2402_ ( .A1(_0314_ ), .A2(fanout_net_8 ), .A3(\myicache.data[5][11] ), .ZN(_0428_ ) );
BUF_X4 _2403_ ( .A(_0088_ ), .Z(_0429_ ) );
NAND3_X1 _2404_ ( .A1(_0234_ ), .A2(_0429_ ), .A3(\myicache.data[1][11] ), .ZN(_0430_ ) );
NAND4_X1 _2405_ ( .A1(_0427_ ), .A2(_0282_ ), .A3(_0428_ ), .A4(_0430_ ), .ZN(_0431_ ) );
NAND3_X1 _2406_ ( .A1(_0424_ ), .A2(_0206_ ), .A3(_0431_ ), .ZN(_0432_ ) );
NAND2_X1 _2407_ ( .A1(_0418_ ), .A2(_0432_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ) );
CLKBUF_X2 _2408_ ( .A(_0185_ ), .Z(_0433_ ) );
OR2_X1 _2409_ ( .A1(_0433_ ), .A2(\rdata [10] ), .ZN(_0434_ ) );
BUF_X4 _2410_ ( .A(_0188_ ), .Z(_0435_ ) );
AOI21_X1 _2411_ ( .A(_0435_ ), .B1(_0416_ ), .B2(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_0436_ ) );
NAND2_X1 _2412_ ( .A1(_0434_ ), .A2(_0436_ ), .ZN(_0437_ ) );
AND3_X1 _2413_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[6][10] ), .ZN(_0438_ ) );
AND3_X1 _2414_ ( .A1(_0274_ ), .A2(fanout_net_4 ), .A3(\myicache.data[2][10] ), .ZN(_0439_ ) );
AOI211_X1 _2415_ ( .A(_0438_ ), .B(_0439_ ), .C1(\myicache.data[0][10] ), .C2(_0391_ ), .ZN(_0440_ ) );
NAND3_X1 _2416_ ( .A1(_0422_ ), .A2(fanout_net_8 ), .A3(\myicache.data[4][10] ), .ZN(_0441_ ) );
NAND4_X1 _2417_ ( .A1(_0440_ ), .A2(_0199_ ), .A3(_0202_ ), .A4(_0441_ ), .ZN(_0442_ ) );
NAND3_X1 _2418_ ( .A1(_0229_ ), .A2(fanout_net_4 ), .A3(\myicache.data[3][10] ), .ZN(_0443_ ) );
NAND3_X1 _2419_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[7][10] ), .ZN(_0444_ ) );
AND2_X1 _2420_ ( .A1(_0443_ ), .A2(_0444_ ), .ZN(_0445_ ) );
NAND3_X1 _2421_ ( .A1(_0314_ ), .A2(fanout_net_8 ), .A3(\myicache.data[5][10] ), .ZN(_0446_ ) );
NAND3_X1 _2422_ ( .A1(_0234_ ), .A2(_0429_ ), .A3(\myicache.data[1][10] ), .ZN(_0447_ ) );
NAND4_X1 _2423_ ( .A1(_0445_ ), .A2(_0282_ ), .A3(_0446_ ), .A4(_0447_ ), .ZN(_0448_ ) );
NAND3_X1 _2424_ ( .A1(_0442_ ), .A2(_0206_ ), .A3(_0448_ ), .ZN(_0449_ ) );
NAND2_X1 _2425_ ( .A1(_0437_ ), .A2(_0449_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ) );
AND3_X1 _2426_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[6][9] ), .ZN(_0450_ ) );
AND3_X1 _2427_ ( .A1(_0207_ ), .A2(fanout_net_4 ), .A3(\myicache.data[2][9] ), .ZN(_0451_ ) );
AOI211_X1 _2428_ ( .A(_0450_ ), .B(_0451_ ), .C1(\myicache.data[0][9] ), .C2(_0240_ ), .ZN(_0452_ ) );
NAND3_X1 _2429_ ( .A1(_0242_ ), .A2(fanout_net_8 ), .A3(\myicache.data[4][9] ), .ZN(_0453_ ) );
NAND4_X1 _2430_ ( .A1(_0452_ ), .A2(_0198_ ), .A3(_0201_ ), .A4(_0453_ ), .ZN(_0454_ ) );
NAND3_X1 _2431_ ( .A1(_0088_ ), .A2(fanout_net_4 ), .A3(\myicache.data[3][9] ), .ZN(_0455_ ) );
NAND3_X1 _2432_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[7][9] ), .ZN(_0456_ ) );
AND2_X1 _2433_ ( .A1(_0455_ ), .A2(_0456_ ), .ZN(_0457_ ) );
NAND3_X1 _2434_ ( .A1(_0242_ ), .A2(fanout_net_8 ), .A3(\myicache.data[5][9] ), .ZN(_0458_ ) );
NAND3_X1 _2435_ ( .A1(_0242_ ), .A2(_0208_ ), .A3(\myicache.data[1][9] ), .ZN(_0459_ ) );
NAND4_X1 _2436_ ( .A1(_0457_ ), .A2(_0248_ ), .A3(_0458_ ), .A4(_0459_ ), .ZN(_0460_ ) );
NAND3_X1 _2437_ ( .A1(_0454_ ), .A2(_0205_ ), .A3(_0460_ ), .ZN(_0461_ ) );
NOR2_X1 _2438_ ( .A1(_0191_ ), .A2(\rdata [9] ), .ZN(_0462_ ) );
OAI21_X1 _2439_ ( .A(\state [2] ), .B1(_0184_ ), .B2(_0955_ ), .ZN(_0463_ ) );
OAI21_X1 _2440_ ( .A(_0461_ ), .B1(_0462_ ), .B2(_0463_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ) );
OR2_X1 _2441_ ( .A1(_0433_ ), .A2(\rdata [7] ), .ZN(_0464_ ) );
AOI21_X1 _2442_ ( .A(_0435_ ), .B1(_0416_ ), .B2(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_0465_ ) );
NAND2_X1 _2443_ ( .A1(_0464_ ), .A2(_0465_ ), .ZN(_0466_ ) );
AND3_X1 _2444_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[6][7] ), .ZN(_0467_ ) );
AND3_X1 _2445_ ( .A1(_0274_ ), .A2(fanout_net_4 ), .A3(\myicache.data[2][7] ), .ZN(_0468_ ) );
AOI211_X1 _2446_ ( .A(_0467_ ), .B(_0468_ ), .C1(\myicache.data[0][7] ), .C2(_0391_ ), .ZN(_0469_ ) );
BUF_X4 _2447_ ( .A(_0198_ ), .Z(_0470_ ) );
BUF_X4 _2448_ ( .A(_0201_ ), .Z(_0471_ ) );
NAND3_X1 _2449_ ( .A1(_0422_ ), .A2(fanout_net_8 ), .A3(\myicache.data[4][7] ), .ZN(_0472_ ) );
NAND4_X1 _2450_ ( .A1(_0469_ ), .A2(_0470_ ), .A3(_0471_ ), .A4(_0472_ ), .ZN(_0473_ ) );
NAND3_X1 _2451_ ( .A1(_0229_ ), .A2(fanout_net_4 ), .A3(\myicache.data[3][7] ), .ZN(_0474_ ) );
NAND3_X1 _2452_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[7][7] ), .ZN(_0475_ ) );
AND2_X1 _2453_ ( .A1(_0474_ ), .A2(_0475_ ), .ZN(_0476_ ) );
NAND3_X1 _2454_ ( .A1(_0314_ ), .A2(fanout_net_8 ), .A3(\myicache.data[5][7] ), .ZN(_0477_ ) );
NAND3_X1 _2455_ ( .A1(_0234_ ), .A2(_0429_ ), .A3(\myicache.data[1][7] ), .ZN(_0478_ ) );
NAND4_X1 _2456_ ( .A1(_0476_ ), .A2(_0282_ ), .A3(_0477_ ), .A4(_0478_ ), .ZN(_0479_ ) );
NAND3_X1 _2457_ ( .A1(_0473_ ), .A2(_0206_ ), .A3(_0479_ ), .ZN(_0480_ ) );
NAND2_X1 _2458_ ( .A1(_0466_ ), .A2(_0480_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ) );
OR2_X1 _2459_ ( .A1(_0433_ ), .A2(\rdata [6] ), .ZN(_0481_ ) );
AOI21_X1 _2460_ ( .A(_0435_ ), .B1(_0416_ ), .B2(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_0482_ ) );
NAND2_X1 _2461_ ( .A1(_0481_ ), .A2(_0482_ ), .ZN(_0483_ ) );
AND3_X1 _2462_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[6][6] ), .ZN(_0484_ ) );
AND3_X1 _2463_ ( .A1(_0274_ ), .A2(fanout_net_4 ), .A3(\myicache.data[2][6] ), .ZN(_0485_ ) );
AOI211_X1 _2464_ ( .A(_0484_ ), .B(_0485_ ), .C1(\myicache.data[0][6] ), .C2(_0391_ ), .ZN(_0486_ ) );
NAND3_X1 _2465_ ( .A1(_0422_ ), .A2(fanout_net_8 ), .A3(\myicache.data[4][6] ), .ZN(_0487_ ) );
NAND4_X1 _2466_ ( .A1(_0486_ ), .A2(_0470_ ), .A3(_0471_ ), .A4(_0487_ ), .ZN(_0488_ ) );
BUF_X4 _2467_ ( .A(_0205_ ), .Z(_0489_ ) );
NAND3_X1 _2468_ ( .A1(_0229_ ), .A2(fanout_net_4 ), .A3(\myicache.data[3][6] ), .ZN(_0490_ ) );
NAND3_X1 _2469_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[7][6] ), .ZN(_0491_ ) );
AND2_X1 _2470_ ( .A1(_0490_ ), .A2(_0491_ ), .ZN(_0492_ ) );
NAND3_X1 _2471_ ( .A1(_0314_ ), .A2(fanout_net_8 ), .A3(\myicache.data[5][6] ), .ZN(_0493_ ) );
NAND3_X1 _2472_ ( .A1(_0234_ ), .A2(_0429_ ), .A3(\myicache.data[1][6] ), .ZN(_0494_ ) );
NAND4_X1 _2473_ ( .A1(_0492_ ), .A2(_0282_ ), .A3(_0493_ ), .A4(_0494_ ), .ZN(_0495_ ) );
NAND3_X1 _2474_ ( .A1(_0488_ ), .A2(_0489_ ), .A3(_0495_ ), .ZN(_0496_ ) );
NAND2_X1 _2475_ ( .A1(_0483_ ), .A2(_0496_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ) );
OR2_X1 _2476_ ( .A1(_0433_ ), .A2(\rdata [5] ), .ZN(_0497_ ) );
AOI21_X1 _2477_ ( .A(_0435_ ), .B1(_0416_ ), .B2(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_0498_ ) );
NAND2_X1 _2478_ ( .A1(_0497_ ), .A2(_0498_ ), .ZN(_0499_ ) );
AND3_X1 _2479_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[6][5] ), .ZN(_0500_ ) );
AND3_X1 _2480_ ( .A1(_0274_ ), .A2(fanout_net_4 ), .A3(\myicache.data[2][5] ), .ZN(_0501_ ) );
AOI211_X1 _2481_ ( .A(_0500_ ), .B(_0501_ ), .C1(\myicache.data[0][5] ), .C2(_0391_ ), .ZN(_0502_ ) );
NAND3_X1 _2482_ ( .A1(_0422_ ), .A2(fanout_net_8 ), .A3(\myicache.data[4][5] ), .ZN(_0503_ ) );
NAND4_X1 _2483_ ( .A1(_0502_ ), .A2(_0470_ ), .A3(_0471_ ), .A4(_0503_ ), .ZN(_0504_ ) );
BUF_X4 _2484_ ( .A(_0207_ ), .Z(_0505_ ) );
NAND3_X1 _2485_ ( .A1(_0505_ ), .A2(fanout_net_4 ), .A3(\myicache.data[3][5] ), .ZN(_0506_ ) );
NAND3_X1 _2486_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[7][5] ), .ZN(_0507_ ) );
AND2_X1 _2487_ ( .A1(_0506_ ), .A2(_0507_ ), .ZN(_0508_ ) );
NAND3_X1 _2488_ ( .A1(_0314_ ), .A2(fanout_net_8 ), .A3(\myicache.data[5][5] ), .ZN(_0509_ ) );
BUF_X4 _2489_ ( .A(_0096_ ), .Z(_0510_ ) );
NAND3_X1 _2490_ ( .A1(_0510_ ), .A2(_0429_ ), .A3(\myicache.data[1][5] ), .ZN(_0511_ ) );
NAND4_X1 _2491_ ( .A1(_0508_ ), .A2(_0282_ ), .A3(_0509_ ), .A4(_0511_ ), .ZN(_0512_ ) );
NAND3_X1 _2492_ ( .A1(_0504_ ), .A2(_0489_ ), .A3(_0512_ ), .ZN(_0513_ ) );
NAND2_X1 _2493_ ( .A1(_0499_ ), .A2(_0513_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ) );
OR2_X1 _2494_ ( .A1(_0433_ ), .A2(\rdata [4] ), .ZN(_0514_ ) );
AOI21_X1 _2495_ ( .A(_0435_ ), .B1(_0416_ ), .B2(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_0515_ ) );
NAND2_X1 _2496_ ( .A1(_0514_ ), .A2(_0515_ ), .ZN(_0516_ ) );
AND3_X1 _2497_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[6][4] ), .ZN(_0517_ ) );
AND3_X1 _2498_ ( .A1(_0274_ ), .A2(fanout_net_4 ), .A3(\myicache.data[2][4] ), .ZN(_0518_ ) );
AOI211_X1 _2499_ ( .A(_0517_ ), .B(_0518_ ), .C1(\myicache.data[0][4] ), .C2(_0391_ ), .ZN(_0519_ ) );
NAND3_X1 _2500_ ( .A1(_0422_ ), .A2(fanout_net_8 ), .A3(\myicache.data[4][4] ), .ZN(_0520_ ) );
NAND4_X1 _2501_ ( .A1(_0519_ ), .A2(_0470_ ), .A3(_0471_ ), .A4(_0520_ ), .ZN(_0521_ ) );
NAND3_X1 _2502_ ( .A1(_0505_ ), .A2(fanout_net_4 ), .A3(\myicache.data[3][4] ), .ZN(_0522_ ) );
NAND3_X1 _2503_ ( .A1(fanout_net_4 ), .A2(fanout_net_8 ), .A3(\myicache.data[7][4] ), .ZN(_0523_ ) );
AND2_X1 _2504_ ( .A1(_0522_ ), .A2(_0523_ ), .ZN(_0524_ ) );
NAND3_X1 _2505_ ( .A1(_0314_ ), .A2(fanout_net_9 ), .A3(\myicache.data[5][4] ), .ZN(_0525_ ) );
NAND3_X1 _2506_ ( .A1(_0510_ ), .A2(_0429_ ), .A3(\myicache.data[1][4] ), .ZN(_0526_ ) );
NAND4_X1 _2507_ ( .A1(_0524_ ), .A2(_0282_ ), .A3(_0525_ ), .A4(_0526_ ), .ZN(_0527_ ) );
NAND3_X1 _2508_ ( .A1(_0521_ ), .A2(_0489_ ), .A3(_0527_ ), .ZN(_0528_ ) );
NAND2_X1 _2509_ ( .A1(_0516_ ), .A2(_0528_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ) );
OR2_X1 _2510_ ( .A1(_0433_ ), .A2(\rdata [3] ), .ZN(_0529_ ) );
AOI21_X1 _2511_ ( .A(_0435_ ), .B1(_0416_ ), .B2(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_0530_ ) );
NAND2_X1 _2512_ ( .A1(_0529_ ), .A2(_0530_ ), .ZN(_0531_ ) );
AND3_X1 _2513_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[6][3] ), .ZN(_0532_ ) );
CLKBUF_X2 _2514_ ( .A(_0087_ ), .Z(_0533_ ) );
AND3_X1 _2515_ ( .A1(_0533_ ), .A2(fanout_net_5 ), .A3(\myicache.data[2][3] ), .ZN(_0534_ ) );
AOI211_X1 _2516_ ( .A(_0532_ ), .B(_0534_ ), .C1(\myicache.data[0][3] ), .C2(_0391_ ), .ZN(_0535_ ) );
NAND3_X1 _2517_ ( .A1(_0422_ ), .A2(fanout_net_9 ), .A3(\myicache.data[4][3] ), .ZN(_0536_ ) );
NAND4_X1 _2518_ ( .A1(_0535_ ), .A2(_0470_ ), .A3(_0471_ ), .A4(_0536_ ), .ZN(_0537_ ) );
NAND3_X1 _2519_ ( .A1(_0505_ ), .A2(fanout_net_5 ), .A3(\myicache.data[3][3] ), .ZN(_0538_ ) );
NAND3_X1 _2520_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[7][3] ), .ZN(_0539_ ) );
AND2_X1 _2521_ ( .A1(_0538_ ), .A2(_0539_ ), .ZN(_0540_ ) );
BUF_X4 _2522_ ( .A(_0212_ ), .Z(_0541_ ) );
NAND3_X1 _2523_ ( .A1(_0314_ ), .A2(fanout_net_9 ), .A3(\myicache.data[5][3] ), .ZN(_0542_ ) );
NAND3_X1 _2524_ ( .A1(_0510_ ), .A2(_0429_ ), .A3(\myicache.data[1][3] ), .ZN(_0543_ ) );
NAND4_X1 _2525_ ( .A1(_0540_ ), .A2(_0541_ ), .A3(_0542_ ), .A4(_0543_ ), .ZN(_0544_ ) );
NAND3_X1 _2526_ ( .A1(_0537_ ), .A2(_0489_ ), .A3(_0544_ ), .ZN(_0545_ ) );
NAND2_X1 _2527_ ( .A1(_0531_ ), .A2(_0545_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ) );
OR2_X1 _2528_ ( .A1(_0433_ ), .A2(\rdata [2] ), .ZN(_0546_ ) );
AOI21_X1 _2529_ ( .A(_0435_ ), .B1(_0416_ ), .B2(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_0547_ ) );
NAND2_X1 _2530_ ( .A1(_0546_ ), .A2(_0547_ ), .ZN(_0548_ ) );
AND3_X1 _2531_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[6][2] ), .ZN(_0549_ ) );
AND3_X1 _2532_ ( .A1(_0533_ ), .A2(fanout_net_5 ), .A3(\myicache.data[2][2] ), .ZN(_0550_ ) );
AOI211_X1 _2533_ ( .A(_0549_ ), .B(_0550_ ), .C1(\myicache.data[0][2] ), .C2(_0391_ ), .ZN(_0551_ ) );
NAND3_X1 _2534_ ( .A1(_0422_ ), .A2(fanout_net_9 ), .A3(\myicache.data[4][2] ), .ZN(_0552_ ) );
NAND4_X1 _2535_ ( .A1(_0551_ ), .A2(_0470_ ), .A3(_0471_ ), .A4(_0552_ ), .ZN(_0553_ ) );
NAND3_X1 _2536_ ( .A1(_0505_ ), .A2(fanout_net_5 ), .A3(\myicache.data[3][2] ), .ZN(_0554_ ) );
NAND3_X1 _2537_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[7][2] ), .ZN(_0555_ ) );
AND2_X1 _2538_ ( .A1(_0554_ ), .A2(_0555_ ), .ZN(_0556_ ) );
NAND3_X1 _2539_ ( .A1(_0217_ ), .A2(fanout_net_9 ), .A3(\myicache.data[5][2] ), .ZN(_0557_ ) );
NAND3_X1 _2540_ ( .A1(_0510_ ), .A2(_0429_ ), .A3(\myicache.data[1][2] ), .ZN(_0558_ ) );
NAND4_X1 _2541_ ( .A1(_0556_ ), .A2(_0541_ ), .A3(_0557_ ), .A4(_0558_ ), .ZN(_0559_ ) );
NAND3_X1 _2542_ ( .A1(_0553_ ), .A2(_0489_ ), .A3(_0559_ ), .ZN(_0560_ ) );
NAND2_X1 _2543_ ( .A1(_0548_ ), .A2(_0560_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ) );
OR2_X1 _2544_ ( .A1(_0433_ ), .A2(\rdata [1] ), .ZN(_0561_ ) );
AOI21_X1 _2545_ ( .A(_0435_ ), .B1(_0416_ ), .B2(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_0562_ ) );
NAND2_X1 _2546_ ( .A1(_0561_ ), .A2(_0562_ ), .ZN(_0563_ ) );
AND3_X1 _2547_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[6][1] ), .ZN(_0564_ ) );
AND3_X1 _2548_ ( .A1(_0533_ ), .A2(fanout_net_5 ), .A3(\myicache.data[2][1] ), .ZN(_0565_ ) );
AOI211_X1 _2549_ ( .A(_0564_ ), .B(_0565_ ), .C1(\myicache.data[0][1] ), .C2(_0391_ ), .ZN(_0566_ ) );
NAND3_X1 _2550_ ( .A1(_0422_ ), .A2(fanout_net_9 ), .A3(\myicache.data[4][1] ), .ZN(_0567_ ) );
NAND4_X1 _2551_ ( .A1(_0566_ ), .A2(_0470_ ), .A3(_0471_ ), .A4(_0567_ ), .ZN(_0568_ ) );
NAND3_X1 _2552_ ( .A1(_0505_ ), .A2(fanout_net_5 ), .A3(\myicache.data[3][1] ), .ZN(_0569_ ) );
NAND3_X1 _2553_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[7][1] ), .ZN(_0570_ ) );
AND2_X1 _2554_ ( .A1(_0569_ ), .A2(_0570_ ), .ZN(_0571_ ) );
NAND3_X1 _2555_ ( .A1(_0217_ ), .A2(fanout_net_9 ), .A3(\myicache.data[5][1] ), .ZN(_0572_ ) );
NAND3_X1 _2556_ ( .A1(_0510_ ), .A2(_0429_ ), .A3(\myicache.data[1][1] ), .ZN(_0573_ ) );
NAND4_X1 _2557_ ( .A1(_0571_ ), .A2(_0541_ ), .A3(_0572_ ), .A4(_0573_ ), .ZN(_0574_ ) );
NAND3_X1 _2558_ ( .A1(_0568_ ), .A2(_0489_ ), .A3(_0574_ ), .ZN(_0575_ ) );
NAND2_X1 _2559_ ( .A1(_0563_ ), .A2(_0575_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ) );
OR2_X1 _2560_ ( .A1(_0433_ ), .A2(\rdata [28] ), .ZN(_0576_ ) );
AOI21_X1 _2561_ ( .A(_0435_ ), .B1(_0416_ ), .B2(pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_0577_ ) );
NAND2_X1 _2562_ ( .A1(_0576_ ), .A2(_0577_ ), .ZN(_0578_ ) );
AND3_X1 _2563_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[6][28] ), .ZN(_0579_ ) );
AND3_X1 _2564_ ( .A1(_0533_ ), .A2(fanout_net_5 ), .A3(\myicache.data[2][28] ), .ZN(_0580_ ) );
AOI211_X1 _2565_ ( .A(_0579_ ), .B(_0580_ ), .C1(\myicache.data[0][28] ), .C2(_0240_ ), .ZN(_0581_ ) );
NAND3_X1 _2566_ ( .A1(_0422_ ), .A2(fanout_net_9 ), .A3(\myicache.data[4][28] ), .ZN(_0582_ ) );
NAND4_X1 _2567_ ( .A1(_0581_ ), .A2(_0470_ ), .A3(_0471_ ), .A4(_0582_ ), .ZN(_0583_ ) );
NAND3_X1 _2568_ ( .A1(_0505_ ), .A2(fanout_net_5 ), .A3(\myicache.data[3][28] ), .ZN(_0584_ ) );
NAND3_X1 _2569_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[7][28] ), .ZN(_0585_ ) );
AND2_X1 _2570_ ( .A1(_0584_ ), .A2(_0585_ ), .ZN(_0586_ ) );
NAND3_X1 _2571_ ( .A1(_0217_ ), .A2(fanout_net_9 ), .A3(\myicache.data[5][28] ), .ZN(_0587_ ) );
NAND3_X1 _2572_ ( .A1(_0510_ ), .A2(_0429_ ), .A3(\myicache.data[1][28] ), .ZN(_0588_ ) );
NAND4_X1 _2573_ ( .A1(_0586_ ), .A2(_0541_ ), .A3(_0587_ ), .A4(_0588_ ), .ZN(_0589_ ) );
NAND3_X1 _2574_ ( .A1(_0583_ ), .A2(_0489_ ), .A3(_0589_ ), .ZN(_0590_ ) );
NAND2_X1 _2575_ ( .A1(_0578_ ), .A2(_0590_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ) );
OR2_X1 _2576_ ( .A1(_0433_ ), .A2(\rdata [0] ), .ZN(_0591_ ) );
AOI21_X1 _2577_ ( .A(_0435_ ), .B1(_0289_ ), .B2(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_0592_ ) );
NAND2_X1 _2578_ ( .A1(_0591_ ), .A2(_0592_ ), .ZN(_0593_ ) );
AND3_X1 _2579_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[6][0] ), .ZN(_0594_ ) );
AND3_X1 _2580_ ( .A1(_0533_ ), .A2(fanout_net_5 ), .A3(\myicache.data[2][0] ), .ZN(_0595_ ) );
AOI211_X1 _2581_ ( .A(_0594_ ), .B(_0595_ ), .C1(\myicache.data[0][0] ), .C2(_0240_ ), .ZN(_0596_ ) );
NAND3_X1 _2582_ ( .A1(_0215_ ), .A2(fanout_net_9 ), .A3(\myicache.data[4][0] ), .ZN(_0597_ ) );
NAND4_X1 _2583_ ( .A1(_0596_ ), .A2(_0470_ ), .A3(_0471_ ), .A4(_0597_ ), .ZN(_0598_ ) );
NAND3_X1 _2584_ ( .A1(_0505_ ), .A2(fanout_net_5 ), .A3(\myicache.data[3][0] ), .ZN(_0599_ ) );
NAND3_X1 _2585_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[7][0] ), .ZN(_0600_ ) );
AND2_X1 _2586_ ( .A1(_0599_ ), .A2(_0600_ ), .ZN(_0601_ ) );
NAND3_X1 _2587_ ( .A1(_0217_ ), .A2(fanout_net_9 ), .A3(\myicache.data[5][0] ), .ZN(_0602_ ) );
NAND3_X1 _2588_ ( .A1(_0510_ ), .A2(_0208_ ), .A3(\myicache.data[1][0] ), .ZN(_0603_ ) );
NAND4_X1 _2589_ ( .A1(_0601_ ), .A2(_0541_ ), .A3(_0602_ ), .A4(_0603_ ), .ZN(_0604_ ) );
NAND3_X1 _2590_ ( .A1(_0598_ ), .A2(_0489_ ), .A3(_0604_ ), .ZN(_0605_ ) );
NAND2_X1 _2591_ ( .A1(_0593_ ), .A2(_0605_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ) );
OR2_X1 _2592_ ( .A1(_0190_ ), .A2(\rdata [27] ), .ZN(_0606_ ) );
AOI21_X1 _2593_ ( .A(_0287_ ), .B1(_0289_ ), .B2(pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_0607_ ) );
NAND2_X1 _2594_ ( .A1(_0606_ ), .A2(_0607_ ), .ZN(_0608_ ) );
AND3_X1 _2595_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[6][27] ), .ZN(_0609_ ) );
AND3_X1 _2596_ ( .A1(_0533_ ), .A2(fanout_net_5 ), .A3(\myicache.data[2][27] ), .ZN(_0610_ ) );
AOI211_X1 _2597_ ( .A(_0609_ ), .B(_0610_ ), .C1(\myicache.data[0][27] ), .C2(_0240_ ), .ZN(_0611_ ) );
NAND3_X1 _2598_ ( .A1(_0215_ ), .A2(fanout_net_9 ), .A3(\myicache.data[4][27] ), .ZN(_0612_ ) );
NAND4_X1 _2599_ ( .A1(_0611_ ), .A2(_0470_ ), .A3(_0471_ ), .A4(_0612_ ), .ZN(_0613_ ) );
NAND3_X1 _2600_ ( .A1(_0505_ ), .A2(fanout_net_5 ), .A3(\myicache.data[3][27] ), .ZN(_0614_ ) );
NAND3_X1 _2601_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[7][27] ), .ZN(_0615_ ) );
AND2_X1 _2602_ ( .A1(_0614_ ), .A2(_0615_ ), .ZN(_0616_ ) );
NAND3_X1 _2603_ ( .A1(_0217_ ), .A2(fanout_net_9 ), .A3(\myicache.data[5][27] ), .ZN(_0617_ ) );
NAND3_X1 _2604_ ( .A1(_0510_ ), .A2(_0208_ ), .A3(\myicache.data[1][27] ), .ZN(_0618_ ) );
NAND4_X1 _2605_ ( .A1(_0616_ ), .A2(_0541_ ), .A3(_0617_ ), .A4(_0618_ ), .ZN(_0619_ ) );
NAND3_X1 _2606_ ( .A1(_0613_ ), .A2(_0489_ ), .A3(_0619_ ), .ZN(_0620_ ) );
NAND2_X1 _2607_ ( .A1(_0608_ ), .A2(_0620_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ) );
AND3_X1 _2608_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[6][26] ), .ZN(_0621_ ) );
AND3_X1 _2609_ ( .A1(_0207_ ), .A2(fanout_net_5 ), .A3(\myicache.data[2][26] ), .ZN(_0622_ ) );
AOI211_X1 _2610_ ( .A(_0621_ ), .B(_0622_ ), .C1(\myicache.data[0][26] ), .C2(_0240_ ), .ZN(_0623_ ) );
NAND3_X1 _2611_ ( .A1(_0242_ ), .A2(fanout_net_9 ), .A3(\myicache.data[4][26] ), .ZN(_0624_ ) );
NAND4_X1 _2612_ ( .A1(_0623_ ), .A2(_0198_ ), .A3(_0201_ ), .A4(_0624_ ), .ZN(_0625_ ) );
NAND3_X1 _2613_ ( .A1(_0088_ ), .A2(fanout_net_5 ), .A3(\myicache.data[3][26] ), .ZN(_0626_ ) );
NAND3_X1 _2614_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[7][26] ), .ZN(_0627_ ) );
AND2_X1 _2615_ ( .A1(_0626_ ), .A2(_0627_ ), .ZN(_0628_ ) );
NAND3_X1 _2616_ ( .A1(_0242_ ), .A2(fanout_net_9 ), .A3(\myicache.data[5][26] ), .ZN(_0629_ ) );
NAND3_X1 _2617_ ( .A1(_0214_ ), .A2(_0208_ ), .A3(\myicache.data[1][26] ), .ZN(_0630_ ) );
NAND4_X1 _2618_ ( .A1(_0628_ ), .A2(_0248_ ), .A3(_0629_ ), .A4(_0630_ ), .ZN(_0631_ ) );
NAND3_X1 _2619_ ( .A1(_0625_ ), .A2(_0205_ ), .A3(_0631_ ), .ZN(_0632_ ) );
NOR2_X1 _2620_ ( .A1(_0191_ ), .A2(\rdata [26] ), .ZN(_0633_ ) );
OAI21_X1 _2621_ ( .A(\state [2] ), .B1(_0184_ ), .B2(_0982_ ), .ZN(_0634_ ) );
OAI21_X1 _2622_ ( .A(_0632_ ), .B1(_0633_ ), .B2(_0634_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ) );
OR2_X1 _2623_ ( .A1(_0190_ ), .A2(\rdata [25] ), .ZN(_0635_ ) );
AOI21_X1 _2624_ ( .A(_0287_ ), .B1(_0289_ ), .B2(pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_0636_ ) );
NAND2_X1 _2625_ ( .A1(_0635_ ), .A2(_0636_ ), .ZN(_0637_ ) );
AND3_X1 _2626_ ( .A1(fanout_net_5 ), .A2(fanout_net_9 ), .A3(\myicache.data[6][25] ), .ZN(_0638_ ) );
AND3_X1 _2627_ ( .A1(_0533_ ), .A2(fanout_net_5 ), .A3(\myicache.data[2][25] ), .ZN(_0639_ ) );
AOI211_X1 _2628_ ( .A(_0638_ ), .B(_0639_ ), .C1(\myicache.data[0][25] ), .C2(_0240_ ), .ZN(_0640_ ) );
NAND3_X1 _2629_ ( .A1(_0215_ ), .A2(fanout_net_6 ), .A3(\myicache.data[4][25] ), .ZN(_0641_ ) );
NAND4_X1 _2630_ ( .A1(_0640_ ), .A2(_0198_ ), .A3(_0201_ ), .A4(_0641_ ), .ZN(_0642_ ) );
NAND3_X1 _2631_ ( .A1(_0505_ ), .A2(fanout_net_2 ), .A3(\myicache.data[3][25] ), .ZN(_0643_ ) );
NAND3_X1 _2632_ ( .A1(fanout_net_2 ), .A2(fanout_net_6 ), .A3(\myicache.data[7][25] ), .ZN(_0644_ ) );
AND2_X1 _2633_ ( .A1(_0643_ ), .A2(_0644_ ), .ZN(_0645_ ) );
NAND3_X1 _2634_ ( .A1(_0217_ ), .A2(fanout_net_6 ), .A3(\myicache.data[5][25] ), .ZN(_0646_ ) );
NAND3_X1 _2635_ ( .A1(_0510_ ), .A2(_0208_ ), .A3(\myicache.data[1][25] ), .ZN(_0647_ ) );
NAND4_X1 _2636_ ( .A1(_0645_ ), .A2(_0541_ ), .A3(_0646_ ), .A4(_0647_ ), .ZN(_0648_ ) );
NAND3_X1 _2637_ ( .A1(_0642_ ), .A2(_0489_ ), .A3(_0648_ ), .ZN(_0649_ ) );
NAND2_X1 _2638_ ( .A1(_0637_ ), .A2(_0649_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ) );
OR2_X1 _2639_ ( .A1(_0190_ ), .A2(\rdata [24] ), .ZN(_0650_ ) );
AOI21_X1 _2640_ ( .A(_0287_ ), .B1(_0289_ ), .B2(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0651_ ) );
NAND2_X1 _2641_ ( .A1(_0650_ ), .A2(_0651_ ), .ZN(_0652_ ) );
AND3_X1 _2642_ ( .A1(fanout_net_2 ), .A2(fanout_net_6 ), .A3(\myicache.data[6][24] ), .ZN(_0653_ ) );
AND3_X1 _2643_ ( .A1(_0533_ ), .A2(fanout_net_2 ), .A3(\myicache.data[2][24] ), .ZN(_0654_ ) );
AOI211_X1 _2644_ ( .A(_0653_ ), .B(_0654_ ), .C1(\myicache.data[0][24] ), .C2(_0240_ ), .ZN(_0655_ ) );
NAND3_X1 _2645_ ( .A1(_0215_ ), .A2(fanout_net_6 ), .A3(\myicache.data[4][24] ), .ZN(_0656_ ) );
NAND4_X1 _2646_ ( .A1(_0655_ ), .A2(_0198_ ), .A3(_0201_ ), .A4(_0656_ ), .ZN(_0657_ ) );
NAND3_X1 _2647_ ( .A1(_0505_ ), .A2(fanout_net_2 ), .A3(\myicache.data[3][24] ), .ZN(_0658_ ) );
NAND3_X1 _2648_ ( .A1(fanout_net_2 ), .A2(fanout_net_6 ), .A3(\myicache.data[7][24] ), .ZN(_0659_ ) );
AND2_X1 _2649_ ( .A1(_0658_ ), .A2(_0659_ ), .ZN(_0660_ ) );
NAND3_X1 _2650_ ( .A1(_0217_ ), .A2(fanout_net_6 ), .A3(\myicache.data[5][24] ), .ZN(_0661_ ) );
NAND3_X1 _2651_ ( .A1(_0510_ ), .A2(_0208_ ), .A3(\myicache.data[1][24] ), .ZN(_0662_ ) );
NAND4_X1 _2652_ ( .A1(_0660_ ), .A2(_0541_ ), .A3(_0661_ ), .A4(_0662_ ), .ZN(_0663_ ) );
NAND3_X1 _2653_ ( .A1(_0657_ ), .A2(_0205_ ), .A3(_0663_ ), .ZN(_0664_ ) );
NAND2_X1 _2654_ ( .A1(_0652_ ), .A2(_0664_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ) );
OR2_X1 _2655_ ( .A1(_0190_ ), .A2(\rdata [23] ), .ZN(_0665_ ) );
AOI21_X1 _2656_ ( .A(_0287_ ), .B1(_0289_ ), .B2(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_A_$_OR__Y_B ), .ZN(_0666_ ) );
NAND2_X1 _2657_ ( .A1(_0665_ ), .A2(_0666_ ), .ZN(_0667_ ) );
AND3_X1 _2658_ ( .A1(fanout_net_2 ), .A2(fanout_net_6 ), .A3(\myicache.data[6][23] ), .ZN(_0668_ ) );
AND3_X1 _2659_ ( .A1(_0533_ ), .A2(fanout_net_2 ), .A3(\myicache.data[2][23] ), .ZN(_0669_ ) );
AOI211_X1 _2660_ ( .A(_0668_ ), .B(_0669_ ), .C1(\myicache.data[0][23] ), .C2(_0240_ ), .ZN(_0670_ ) );
NAND3_X1 _2661_ ( .A1(_0215_ ), .A2(fanout_net_6 ), .A3(\myicache.data[4][23] ), .ZN(_0671_ ) );
NAND4_X1 _2662_ ( .A1(_0670_ ), .A2(_0198_ ), .A3(_0201_ ), .A4(_0671_ ), .ZN(_0672_ ) );
NAND3_X1 _2663_ ( .A1(_0088_ ), .A2(fanout_net_2 ), .A3(\myicache.data[3][23] ), .ZN(_0673_ ) );
NAND3_X1 _2664_ ( .A1(fanout_net_2 ), .A2(fanout_net_6 ), .A3(\myicache.data[7][23] ), .ZN(_0674_ ) );
AND2_X1 _2665_ ( .A1(_0673_ ), .A2(_0674_ ), .ZN(_0675_ ) );
NAND3_X1 _2666_ ( .A1(_0217_ ), .A2(fanout_net_6 ), .A3(\myicache.data[5][23] ), .ZN(_0676_ ) );
NAND3_X1 _2667_ ( .A1(_0242_ ), .A2(_0208_ ), .A3(\myicache.data[1][23] ), .ZN(_0677_ ) );
NAND4_X1 _2668_ ( .A1(_0675_ ), .A2(_0541_ ), .A3(_0676_ ), .A4(_0677_ ), .ZN(_0678_ ) );
NAND3_X1 _2669_ ( .A1(_0672_ ), .A2(_0205_ ), .A3(_0678_ ), .ZN(_0679_ ) );
NAND2_X1 _2670_ ( .A1(_0667_ ), .A2(_0679_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ) );
OR2_X1 _2671_ ( .A1(_0190_ ), .A2(\rdata [22] ), .ZN(_0680_ ) );
AOI21_X1 _2672_ ( .A(_0287_ ), .B1(_0289_ ), .B2(pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .ZN(_0681_ ) );
NAND2_X1 _2673_ ( .A1(_0680_ ), .A2(_0681_ ), .ZN(_0682_ ) );
AND3_X1 _2674_ ( .A1(fanout_net_2 ), .A2(fanout_net_6 ), .A3(\myicache.data[6][22] ), .ZN(_0683_ ) );
AND3_X1 _2675_ ( .A1(_0533_ ), .A2(fanout_net_2 ), .A3(\myicache.data[2][22] ), .ZN(_0684_ ) );
AOI211_X1 _2676_ ( .A(_0683_ ), .B(_0684_ ), .C1(\myicache.data[0][22] ), .C2(_0240_ ), .ZN(_0685_ ) );
NAND3_X1 _2677_ ( .A1(_0215_ ), .A2(fanout_net_6 ), .A3(\myicache.data[4][22] ), .ZN(_0686_ ) );
NAND4_X1 _2678_ ( .A1(_0685_ ), .A2(_0198_ ), .A3(_0201_ ), .A4(_0686_ ), .ZN(_0687_ ) );
NAND3_X1 _2679_ ( .A1(_0088_ ), .A2(fanout_net_2 ), .A3(\myicache.data[3][22] ), .ZN(_0688_ ) );
NAND3_X1 _2680_ ( .A1(fanout_net_2 ), .A2(fanout_net_6 ), .A3(\myicache.data[7][22] ), .ZN(_0689_ ) );
AND2_X1 _2681_ ( .A1(_0688_ ), .A2(_0689_ ), .ZN(_0690_ ) );
NAND3_X1 _2682_ ( .A1(_0217_ ), .A2(fanout_net_6 ), .A3(\myicache.data[5][22] ), .ZN(_0691_ ) );
NAND3_X1 _2683_ ( .A1(_0242_ ), .A2(_0208_ ), .A3(\myicache.data[1][22] ), .ZN(_0692_ ) );
NAND4_X1 _2684_ ( .A1(_0690_ ), .A2(_0541_ ), .A3(_0691_ ), .A4(_0692_ ), .ZN(_0693_ ) );
NAND3_X1 _2685_ ( .A1(_0687_ ), .A2(_0205_ ), .A3(_0693_ ), .ZN(_0694_ ) );
NAND2_X1 _2686_ ( .A1(_0682_ ), .A2(_0694_ ), .ZN(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ) );
AOI21_X1 _2687_ ( .A(_0090_ ), .B1(_1123_ ), .B2(_1138_ ), .ZN(pc_$_SDFFE_PP0P__Q_30_E ) );
INV_X1 _2688_ ( .A(fanout_net_10 ), .ZN(_0695_ ) );
OR2_X1 _2689_ ( .A1(_0695_ ), .A2(\myicache.tag[1][12] ), .ZN(_0696_ ) );
INV_X1 _2690_ ( .A(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_0697_ ) );
OAI211_X1 _2691_ ( .A(_0696_ ), .B(_0697_ ), .C1(fanout_net_10 ), .C2(\myicache.tag[0][12] ), .ZN(_0698_ ) );
OR2_X1 _2692_ ( .A1(_0695_ ), .A2(\myicache.tag[3][12] ), .ZN(_0699_ ) );
OAI211_X1 _2693_ ( .A(_0699_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_10 ), .C2(\myicache.tag[2][12] ), .ZN(_0700_ ) );
AND3_X1 _2694_ ( .A1(_0698_ ), .A2(_0700_ ), .A3(\araddr [17] ), .ZN(_0701_ ) );
MUX2_X1 _2695_ ( .A(\myicache.tag[2][10] ), .B(\myicache.tag[3][10] ), .S(fanout_net_10 ), .Z(_0702_ ) );
OR2_X1 _2696_ ( .A1(_0702_ ), .A2(_0697_ ), .ZN(_0703_ ) );
MUX2_X1 _2697_ ( .A(\myicache.tag[0][10] ), .B(\myicache.tag[1][10] ), .S(fanout_net_10 ), .Z(_0704_ ) );
OR2_X1 _2698_ ( .A1(_0704_ ), .A2(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_0705_ ) );
AND3_X1 _2699_ ( .A1(_0703_ ), .A2(_0705_ ), .A3(_0918_ ), .ZN(_0706_ ) );
OR2_X1 _2700_ ( .A1(_0695_ ), .A2(\myicache.tag[1][18] ), .ZN(_0707_ ) );
OAI211_X1 _2701_ ( .A(_0707_ ), .B(_0697_ ), .C1(fanout_net_10 ), .C2(\myicache.tag[0][18] ), .ZN(_0708_ ) );
OR2_X1 _2702_ ( .A1(_0695_ ), .A2(\myicache.tag[3][18] ), .ZN(_0709_ ) );
OAI211_X1 _2703_ ( .A(_0709_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_10 ), .C2(\myicache.tag[2][18] ), .ZN(_0710_ ) );
AND3_X1 _2704_ ( .A1(_0708_ ), .A2(_0710_ ), .A3(\araddr [23] ), .ZN(_0711_ ) );
AOI21_X1 _2705_ ( .A(\araddr [17] ), .B1(_0698_ ), .B2(_0700_ ), .ZN(_0712_ ) );
OR4_X1 _2706_ ( .A1(_0701_ ), .A2(_0706_ ), .A3(_0711_ ), .A4(_0712_ ), .ZN(_0713_ ) );
NAND2_X1 _2707_ ( .A1(_0708_ ), .A2(_0710_ ), .ZN(_0714_ ) );
NAND2_X1 _2708_ ( .A1(_0714_ ), .A2(_1022_ ), .ZN(_0715_ ) );
MUX2_X1 _2709_ ( .A(\myicache.tag[2][22] ), .B(\myicache.tag[3][22] ), .S(fanout_net_10 ), .Z(_0716_ ) );
AND2_X1 _2710_ ( .A1(_0716_ ), .A2(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_0717_ ) );
BUF_X2 _2711_ ( .A(_0697_ ), .Z(_0718_ ) );
BUF_X2 _2712_ ( .A(_0718_ ), .Z(_0719_ ) );
MUX2_X1 _2713_ ( .A(\myicache.tag[0][22] ), .B(\myicache.tag[1][22] ), .S(fanout_net_10 ), .Z(_0720_ ) );
AOI21_X1 _2714_ ( .A(_0717_ ), .B1(_0719_ ), .B2(_0720_ ), .ZN(_0721_ ) );
OAI21_X1 _2715_ ( .A(_0715_ ), .B1(_0721_ ), .B2(\araddr [27] ), .ZN(_0722_ ) );
MUX2_X1 _2716_ ( .A(\myicache.tag[2][5] ), .B(\myicache.tag[3][5] ), .S(fanout_net_10 ), .Z(_0723_ ) );
OR2_X1 _2717_ ( .A1(_0723_ ), .A2(_0718_ ), .ZN(_0724_ ) );
MUX2_X1 _2718_ ( .A(\myicache.tag[0][5] ), .B(\myicache.tag[1][5] ), .S(fanout_net_10 ), .Z(_0725_ ) );
OAI21_X1 _2719_ ( .A(_0724_ ), .B1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_0725_ ), .ZN(_0726_ ) );
MUX2_X1 _2720_ ( .A(\myicache.tag[0][20] ), .B(\myicache.tag[1][20] ), .S(fanout_net_10 ), .Z(_0727_ ) );
MUX2_X1 _2721_ ( .A(\myicache.tag[2][20] ), .B(\myicache.tag[3][20] ), .S(fanout_net_10 ), .Z(_0728_ ) );
MUX2_X1 _2722_ ( .A(_0727_ ), .B(_0728_ ), .S(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_0729_ ) );
OAI22_X1 _2723_ ( .A1(_0726_ ), .A2(\araddr [10] ), .B1(_0906_ ), .B2(_0729_ ), .ZN(_0730_ ) );
OR3_X1 _2724_ ( .A1(_0713_ ), .A2(_0722_ ), .A3(_0730_ ), .ZN(_0731_ ) );
CLKBUF_X2 _2725_ ( .A(_0695_ ), .Z(_0732_ ) );
OR2_X1 _2726_ ( .A1(_0732_ ), .A2(\myicache.tag[1][9] ), .ZN(_0733_ ) );
OAI211_X1 _2727_ ( .A(_0733_ ), .B(_0718_ ), .C1(fanout_net_10 ), .C2(\myicache.tag[0][9] ), .ZN(_0734_ ) );
OR2_X1 _2728_ ( .A1(_0732_ ), .A2(\myicache.tag[3][9] ), .ZN(_0735_ ) );
OAI211_X1 _2729_ ( .A(_0735_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_10 ), .C2(\myicache.tag[2][9] ), .ZN(_0736_ ) );
NAND3_X1 _2730_ ( .A1(_0734_ ), .A2(_0736_ ), .A3(\araddr [14] ), .ZN(_0737_ ) );
MUX2_X1 _2731_ ( .A(\myicache.tag[2][13] ), .B(\myicache.tag[3][13] ), .S(fanout_net_10 ), .Z(_0738_ ) );
OR2_X1 _2732_ ( .A1(_0738_ ), .A2(_0719_ ), .ZN(_0739_ ) );
MUX2_X1 _2733_ ( .A(\myicache.tag[0][13] ), .B(\myicache.tag[1][13] ), .S(fanout_net_10 ), .Z(_0740_ ) );
OAI21_X1 _2734_ ( .A(_0739_ ), .B1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_0740_ ), .ZN(_0741_ ) );
MUX2_X1 _2735_ ( .A(\myicache.tag[2][16] ), .B(\myicache.tag[3][16] ), .S(fanout_net_10 ), .Z(_0742_ ) );
OR2_X1 _2736_ ( .A1(_0742_ ), .A2(_0719_ ), .ZN(_0743_ ) );
MUX2_X1 _2737_ ( .A(\myicache.tag[0][16] ), .B(\myicache.tag[1][16] ), .S(fanout_net_10 ), .Z(_0744_ ) );
OAI21_X1 _2738_ ( .A(_0743_ ), .B1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_0744_ ), .ZN(_0745_ ) );
OAI221_X1 _2739_ ( .A(_0737_ ), .B1(_0741_ ), .B2(\araddr [18] ), .C1(_0745_ ), .C2(\araddr [21] ), .ZN(_0746_ ) );
MUX2_X1 _2740_ ( .A(\myicache.tag[0][7] ), .B(\myicache.tag[1][7] ), .S(fanout_net_10 ), .Z(_0747_ ) );
MUX2_X1 _2741_ ( .A(\myicache.tag[2][7] ), .B(\myicache.tag[3][7] ), .S(fanout_net_10 ), .Z(_0748_ ) );
MUX2_X1 _2742_ ( .A(_0747_ ), .B(_0748_ ), .S(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_0749_ ) );
NOR2_X1 _2743_ ( .A1(_0749_ ), .A2(_1001_ ), .ZN(_0750_ ) );
MUX2_X1 _2744_ ( .A(\myicache.tag[2][11] ), .B(\myicache.tag[3][11] ), .S(fanout_net_10 ), .Z(_0751_ ) );
AND2_X1 _2745_ ( .A1(_0751_ ), .A2(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_0752_ ) );
MUX2_X1 _2746_ ( .A(\myicache.tag[0][11] ), .B(\myicache.tag[1][11] ), .S(fanout_net_10 ), .Z(_0753_ ) );
AOI21_X1 _2747_ ( .A(_0752_ ), .B1(_0718_ ), .B2(_0753_ ), .ZN(_0754_ ) );
AND2_X1 _2748_ ( .A1(_0754_ ), .A2(\araddr [16] ), .ZN(_0755_ ) );
MUX2_X1 _2749_ ( .A(\myicache.tag[2][0] ), .B(\myicache.tag[3][0] ), .S(fanout_net_10 ), .Z(_0756_ ) );
OR2_X1 _2750_ ( .A1(_0756_ ), .A2(_0718_ ), .ZN(_0757_ ) );
MUX2_X1 _2751_ ( .A(\myicache.tag[0][0] ), .B(\myicache.tag[1][0] ), .S(fanout_net_10 ), .Z(_0758_ ) );
OR2_X1 _2752_ ( .A1(_0758_ ), .A2(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_0759_ ) );
AND3_X1 _2753_ ( .A1(_0757_ ), .A2(_0759_ ), .A3(pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_0760_ ) );
AOI21_X1 _2754_ ( .A(\araddr [14] ), .B1(_0734_ ), .B2(_0736_ ), .ZN(_0761_ ) );
OR4_X1 _2755_ ( .A1(_0750_ ), .A2(_0755_ ), .A3(_0760_ ), .A4(_0761_ ), .ZN(_0762_ ) );
NOR3_X1 _2756_ ( .A1(_0731_ ), .A2(_0746_ ), .A3(_0762_ ), .ZN(_0763_ ) );
NOR2_X1 _2757_ ( .A1(_0754_ ), .A2(\araddr [16] ), .ZN(_0764_ ) );
AOI21_X1 _2758_ ( .A(_0764_ ), .B1(\araddr [18] ), .B2(_0741_ ), .ZN(_0765_ ) );
MUX2_X1 _2759_ ( .A(\myicache.tag[0][3] ), .B(\myicache.tag[1][3] ), .S(fanout_net_10 ), .Z(_0766_ ) );
MUX2_X1 _2760_ ( .A(\myicache.tag[2][3] ), .B(\myicache.tag[3][3] ), .S(fanout_net_10 ), .Z(_0767_ ) );
MUX2_X1 _2761_ ( .A(_0766_ ), .B(_0767_ ), .S(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_0768_ ) );
XNOR2_X1 _2762_ ( .A(_0768_ ), .B(\araddr [8] ), .ZN(_0769_ ) );
AOI22_X1 _2763_ ( .A1(_0745_ ), .A2(\araddr [21] ), .B1(_0749_ ), .B2(_1001_ ), .ZN(_0770_ ) );
MUX2_X1 _2764_ ( .A(\myicache.tag[2][15] ), .B(\myicache.tag[3][15] ), .S(fanout_net_10 ), .Z(_0771_ ) );
OR2_X1 _2765_ ( .A1(_0771_ ), .A2(_0718_ ), .ZN(_0772_ ) );
MUX2_X1 _2766_ ( .A(\myicache.tag[0][15] ), .B(\myicache.tag[1][15] ), .S(fanout_net_10 ), .Z(_0773_ ) );
OAI21_X1 _2767_ ( .A(_0772_ ), .B1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_0773_ ), .ZN(_0774_ ) );
AOI22_X1 _2768_ ( .A1(\araddr [27] ), .A2(_0721_ ), .B1(_0774_ ), .B2(\araddr [20] ), .ZN(_0775_ ) );
NAND4_X1 _2769_ ( .A1(_0765_ ), .A2(_0769_ ), .A3(_0770_ ), .A4(_0775_ ), .ZN(_0776_ ) );
CLKBUF_X2 _2770_ ( .A(_0695_ ), .Z(_0777_ ) );
OR2_X1 _2771_ ( .A1(_0777_ ), .A2(\myicache.tag[1][1] ), .ZN(_0778_ ) );
OAI211_X1 _2772_ ( .A(_0778_ ), .B(_0719_ ), .C1(fanout_net_10 ), .C2(\myicache.tag[0][1] ), .ZN(_0779_ ) );
OR2_X1 _2773_ ( .A1(_0777_ ), .A2(\myicache.tag[3][1] ), .ZN(_0780_ ) );
OAI211_X1 _2774_ ( .A(_0780_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[2][1] ), .ZN(_0781_ ) );
AOI21_X1 _2775_ ( .A(\araddr [6] ), .B1(_0779_ ), .B2(_0781_ ), .ZN(_0782_ ) );
AOI21_X1 _2776_ ( .A(_0918_ ), .B1(_0703_ ), .B2(_0705_ ), .ZN(_0783_ ) );
OR2_X1 _2777_ ( .A1(_0732_ ), .A2(\myicache.tag[1][6] ), .ZN(_0784_ ) );
OAI211_X1 _2778_ ( .A(_0784_ ), .B(_0718_ ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[0][6] ), .ZN(_0785_ ) );
OR2_X1 _2779_ ( .A1(_0695_ ), .A2(\myicache.tag[3][6] ), .ZN(_0786_ ) );
OAI211_X1 _2780_ ( .A(_0786_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[2][6] ), .ZN(_0787_ ) );
AND3_X1 _2781_ ( .A1(_0785_ ), .A2(_0787_ ), .A3(\araddr [11] ), .ZN(_0788_ ) );
AOI21_X1 _2782_ ( .A(\araddr [11] ), .B1(_0785_ ), .B2(_0787_ ), .ZN(_0789_ ) );
OR4_X1 _2783_ ( .A1(_0782_ ), .A2(_0783_ ), .A3(_0788_ ), .A4(_0789_ ), .ZN(_0790_ ) );
OR2_X1 _2784_ ( .A1(_0774_ ), .A2(\araddr [20] ), .ZN(_0791_ ) );
NAND2_X1 _2785_ ( .A1(_0729_ ), .A2(_0906_ ), .ZN(_0792_ ) );
NAND3_X1 _2786_ ( .A1(_0779_ ), .A2(_0781_ ), .A3(\araddr [6] ), .ZN(_0793_ ) );
NAND2_X1 _2787_ ( .A1(_0726_ ), .A2(\araddr [10] ), .ZN(_0794_ ) );
NAND4_X1 _2788_ ( .A1(_0791_ ), .A2(_0792_ ), .A3(_0793_ ), .A4(_0794_ ), .ZN(_0795_ ) );
NOR3_X1 _2789_ ( .A1(_0776_ ), .A2(_0790_ ), .A3(_0795_ ), .ZN(_0796_ ) );
AND2_X1 _2790_ ( .A1(_0763_ ), .A2(_0796_ ), .ZN(_0797_ ) );
OR2_X1 _2791_ ( .A1(_0777_ ), .A2(\myicache.tag[1][21] ), .ZN(_0798_ ) );
OAI211_X1 _2792_ ( .A(_0798_ ), .B(_0719_ ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[0][21] ), .ZN(_0799_ ) );
OR2_X1 _2793_ ( .A1(_0777_ ), .A2(\myicache.tag[3][21] ), .ZN(_0800_ ) );
OAI211_X1 _2794_ ( .A(_0800_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[2][21] ), .ZN(_0801_ ) );
NAND2_X1 _2795_ ( .A1(_0799_ ), .A2(_0801_ ), .ZN(_0802_ ) );
XNOR2_X1 _2796_ ( .A(_0802_ ), .B(\araddr [26] ), .ZN(_0803_ ) );
OR2_X1 _2797_ ( .A1(_0777_ ), .A2(\myicache.tag[1][14] ), .ZN(_0804_ ) );
OAI211_X1 _2798_ ( .A(_0804_ ), .B(_0719_ ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[0][14] ), .ZN(_0805_ ) );
OR2_X1 _2799_ ( .A1(_0732_ ), .A2(\myicache.tag[3][14] ), .ZN(_0806_ ) );
OAI211_X1 _2800_ ( .A(_0806_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[2][14] ), .ZN(_0807_ ) );
NAND2_X1 _2801_ ( .A1(_0805_ ), .A2(_0807_ ), .ZN(_0808_ ) );
XNOR2_X1 _2802_ ( .A(_0808_ ), .B(\araddr [19] ), .ZN(_0809_ ) );
OR2_X1 _2803_ ( .A1(_0732_ ), .A2(\myicache.tag[1][26] ), .ZN(_0810_ ) );
OAI211_X1 _2804_ ( .A(_0810_ ), .B(_0719_ ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[0][26] ), .ZN(_0811_ ) );
OR2_X1 _2805_ ( .A1(_0732_ ), .A2(\myicache.tag[3][26] ), .ZN(_0812_ ) );
OAI211_X1 _2806_ ( .A(_0812_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[2][26] ), .ZN(_0813_ ) );
NAND2_X1 _2807_ ( .A1(_0811_ ), .A2(_0813_ ), .ZN(_0814_ ) );
XNOR2_X1 _2808_ ( .A(_0814_ ), .B(\araddr [31] ), .ZN(_0815_ ) );
OR2_X1 _2809_ ( .A1(_0732_ ), .A2(\myicache.tag[1][23] ), .ZN(_0816_ ) );
OAI211_X1 _2810_ ( .A(_0816_ ), .B(_0718_ ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[0][23] ), .ZN(_0817_ ) );
OR2_X1 _2811_ ( .A1(_0732_ ), .A2(\myicache.tag[3][23] ), .ZN(_0818_ ) );
OAI211_X1 _2812_ ( .A(_0818_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[2][23] ), .ZN(_0819_ ) );
NAND2_X1 _2813_ ( .A1(_0817_ ), .A2(_0819_ ), .ZN(_0820_ ) );
XNOR2_X1 _2814_ ( .A(_0820_ ), .B(\araddr [28] ), .ZN(_0821_ ) );
AND4_X1 _2815_ ( .A1(_0803_ ), .A2(_0809_ ), .A3(_0815_ ), .A4(_0821_ ), .ZN(_0822_ ) );
OR2_X1 _2816_ ( .A1(_0732_ ), .A2(\myicache.tag[1][2] ), .ZN(_0823_ ) );
OAI211_X1 _2817_ ( .A(_0823_ ), .B(_0719_ ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[0][2] ), .ZN(_0824_ ) );
OR2_X1 _2818_ ( .A1(_0732_ ), .A2(\myicache.tag[3][2] ), .ZN(_0825_ ) );
OAI211_X1 _2819_ ( .A(_0825_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[2][2] ), .ZN(_0826_ ) );
NAND2_X1 _2820_ ( .A1(_0824_ ), .A2(_0826_ ), .ZN(_0827_ ) );
XNOR2_X1 _2821_ ( .A(_0827_ ), .B(\araddr [7] ), .ZN(_0828_ ) );
OR2_X1 _2822_ ( .A1(_0695_ ), .A2(\myicache.tag[1][25] ), .ZN(_0829_ ) );
OAI211_X1 _2823_ ( .A(_0829_ ), .B(_0718_ ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[0][25] ), .ZN(_0830_ ) );
OR2_X1 _2824_ ( .A1(_0695_ ), .A2(\myicache.tag[3][25] ), .ZN(_0831_ ) );
OAI211_X1 _2825_ ( .A(_0831_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[2][25] ), .ZN(_0832_ ) );
NAND2_X1 _2826_ ( .A1(_0830_ ), .A2(_0832_ ), .ZN(_0833_ ) );
XNOR2_X1 _2827_ ( .A(_0833_ ), .B(\araddr [30] ), .ZN(_0834_ ) );
OR2_X1 _2828_ ( .A1(_0695_ ), .A2(\myicache.tag[3][4] ), .ZN(_0835_ ) );
OAI211_X1 _2829_ ( .A(_0835_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[2][4] ), .ZN(_0836_ ) );
OR2_X1 _2830_ ( .A1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myicache.tag[0][4] ), .ZN(_0837_ ) );
OAI211_X1 _2831_ ( .A(_0837_ ), .B(_0718_ ), .C1(_0777_ ), .C2(\myicache.tag[1][4] ), .ZN(_0838_ ) );
NAND2_X1 _2832_ ( .A1(_0836_ ), .A2(_0838_ ), .ZN(_0839_ ) );
XNOR2_X1 _2833_ ( .A(_0839_ ), .B(\araddr [9] ), .ZN(_0840_ ) );
AND2_X1 _2834_ ( .A1(_0834_ ), .A2(_0840_ ), .ZN(_0841_ ) );
MUX2_X1 _2835_ ( .A(\myicache.valid [0] ), .B(\myicache.valid [1] ), .S(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_0842_ ) );
MUX2_X1 _2836_ ( .A(\myicache.valid [2] ), .B(\myicache.valid [3] ), .S(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_0843_ ) );
MUX2_X1 _2837_ ( .A(_0842_ ), .B(_0843_ ), .S(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_0844_ ) );
OR2_X1 _2838_ ( .A1(_0777_ ), .A2(\myicache.tag[1][17] ), .ZN(_0845_ ) );
OAI211_X1 _2839_ ( .A(_0845_ ), .B(_0719_ ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[0][17] ), .ZN(_0846_ ) );
OR2_X1 _2840_ ( .A1(_0777_ ), .A2(\myicache.tag[3][17] ), .ZN(_0847_ ) );
OAI211_X1 _2841_ ( .A(_0847_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[2][17] ), .ZN(_0848_ ) );
NAND3_X1 _2842_ ( .A1(_0846_ ), .A2(_0848_ ), .A3(\araddr [22] ), .ZN(_0849_ ) );
AND4_X1 _2843_ ( .A1(_0828_ ), .A2(_0841_ ), .A3(_0844_ ), .A4(_0849_ ), .ZN(_0850_ ) );
MUX2_X1 _2844_ ( .A(\myicache.tag[0][24] ), .B(\myicache.tag[1][24] ), .S(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_0851_ ) );
MUX2_X1 _2845_ ( .A(\myicache.tag[2][24] ), .B(\myicache.tag[3][24] ), .S(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_0852_ ) );
MUX2_X1 _2846_ ( .A(_0851_ ), .B(_0852_ ), .S(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_0853_ ) );
XNOR2_X1 _2847_ ( .A(_0853_ ), .B(\araddr [29] ), .ZN(_0854_ ) );
MUX2_X1 _2848_ ( .A(\myicache.tag[0][8] ), .B(\myicache.tag[1][8] ), .S(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_0855_ ) );
MUX2_X1 _2849_ ( .A(\myicache.tag[2][8] ), .B(\myicache.tag[3][8] ), .S(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_0856_ ) );
MUX2_X1 _2850_ ( .A(_0855_ ), .B(_0856_ ), .S(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_0857_ ) );
XNOR2_X1 _2851_ ( .A(_0857_ ), .B(\araddr [13] ), .ZN(_0858_ ) );
AND2_X1 _2852_ ( .A1(_0854_ ), .A2(_0858_ ), .ZN(_0859_ ) );
AOI21_X1 _2853_ ( .A(pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_0757_ ), .B2(_0759_ ), .ZN(_0860_ ) );
OR2_X1 _2854_ ( .A1(_0777_ ), .A2(\myicache.tag[1][19] ), .ZN(_0861_ ) );
OAI211_X1 _2855_ ( .A(_0861_ ), .B(_0719_ ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[0][19] ), .ZN(_0862_ ) );
OR2_X1 _2856_ ( .A1(_0777_ ), .A2(\myicache.tag[3][19] ), .ZN(_0863_ ) );
OAI211_X1 _2857_ ( .A(_0863_ ), .B(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myicache.tag[2][19] ), .ZN(_0864_ ) );
AND3_X1 _2858_ ( .A1(_0862_ ), .A2(_0864_ ), .A3(\araddr [24] ), .ZN(_0865_ ) );
AOI21_X1 _2859_ ( .A(\araddr [22] ), .B1(_0846_ ), .B2(_0848_ ), .ZN(_0866_ ) );
AOI21_X1 _2860_ ( .A(\araddr [24] ), .B1(_0862_ ), .B2(_0864_ ), .ZN(_0867_ ) );
NOR4_X1 _2861_ ( .A1(_0860_ ), .A2(_0865_ ), .A3(_0866_ ), .A4(_0867_ ), .ZN(_0868_ ) );
AND4_X1 _2862_ ( .A1(_0822_ ), .A2(_0850_ ), .A3(_0859_ ), .A4(_0868_ ), .ZN(_0869_ ) );
AND2_X1 _2863_ ( .A1(_0797_ ), .A2(_0869_ ), .ZN(_0870_ ) );
OAI21_X1 _2864_ ( .A(_0189_ ), .B1(_0870_ ), .B2(_0172_ ), .ZN(rmem_quest ) );
AOI21_X1 _2865_ ( .A(_0173_ ), .B1(readyFromIDU ), .B2(to_reset ), .ZN(_0871_ ) );
AND2_X1 _2866_ ( .A1(\state [0] ), .A2(stall_quest_fencei ), .ZN(_0872_ ) );
NOR2_X1 _2867_ ( .A1(_0871_ ), .A2(_0872_ ), .ZN(_0873_ ) );
OAI211_X1 _2868_ ( .A(_0873_ ), .B(_1181_ ), .C1(\state [0] ), .C2(_0291_ ), .ZN(_0874_ ) );
INV_X1 _2869_ ( .A(_0870_ ), .ZN(_0875_ ) );
AOI21_X1 _2870_ ( .A(_0874_ ), .B1(_0875_ ), .B2(\state [0] ), .ZN(rmem_quest_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y ) );
INV_X1 _2871_ ( .A(_0797_ ), .ZN(_0876_ ) );
INV_X1 _2872_ ( .A(_0869_ ), .ZN(_0877_ ) );
OAI21_X1 _2873_ ( .A(arvalid ), .B1(_0876_ ), .B2(_0877_ ), .ZN(_0878_ ) );
NAND2_X1 _2874_ ( .A1(_0878_ ), .A2(_0189_ ), .ZN(rready ) );
NAND4_X1 _2875_ ( .A1(_0763_ ), .A2(_0869_ ), .A3(arvalid ), .A4(_0796_ ), .ZN(_0879_ ) );
AND4_X1 _2876_ ( .A1(\state [2] ), .A2(_0155_ ), .A3(rlast ), .A4(_0157_ ), .ZN(_0880_ ) );
OAI21_X1 _2877_ ( .A(_1181_ ), .B1(_0880_ ), .B2(_0174_ ), .ZN(_0881_ ) );
NAND2_X1 _2878_ ( .A1(_0879_ ), .A2(_0881_ ), .ZN(state_$_DFF_P__Q_1_D ) );
NOR2_X1 _2879_ ( .A1(_0878_ ), .A2(arready ), .ZN(_0882_ ) );
OR4_X1 _2880_ ( .A1(reset ), .A2(_0882_ ), .A3(readyFromIDU_$_AND__B_Y ), .A4(_0872_ ), .ZN(state_$_DFF_P__Q_2_D ) );
NAND3_X1 _2881_ ( .A1(_0159_ ), .A2(_1181_ ), .A3(\state [2] ), .ZN(_0883_ ) );
INV_X1 _2882_ ( .A(arready ), .ZN(_0884_ ) );
OAI21_X1 _2883_ ( .A(_0883_ ), .B1(_0878_ ), .B2(_0884_ ), .ZN(state_$_DFF_P__Q_D ) );
AND3_X1 _2884_ ( .A1(_0155_ ), .A2(\state [2] ), .A3(_0157_ ), .ZN(tmp_offset_$_SDFFE_PP0P__Q_E ) );
AOI21_X1 _2885_ ( .A(_0176_ ), .B1(_1115_ ), .B2(check_quest ), .ZN(validToIDU ) );
AND3_X1 _2886_ ( .A1(wen_$_ANDNOT__A_Y ), .A2(_0166_ ), .A3(_0213_ ), .ZN(wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
AND4_X1 _2887_ ( .A1(wen_$_ANDNOT__A_Y ), .A2(_0166_ ), .A3(_0199_ ), .A4(_0202_ ), .ZN(wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ) );
NOR4_X1 _2888_ ( .A1(_0213_ ), .A2(_0167_ ), .A3(_0170_ ), .A4(_0179_ ), .ZN(wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _2889_ ( .A1(fanout_net_2 ), .A2(wen_$_ANDNOT__A_Y ), .A3(fanout_net_6 ), .A4(_0213_ ), .ZN(wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ) );
AND4_X1 _2890_ ( .A1(fanout_net_2 ), .A2(wen_$_ANDNOT__A_Y ), .A3(_0089_ ), .A4(_0213_ ), .ZN(wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ) );
NOR4_X1 _2891_ ( .A1(_0213_ ), .A2(_0167_ ), .A3(_0170_ ), .A4(_0171_ ), .ZN(wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ) );
AND4_X1 _2892_ ( .A1(_0097_ ), .A2(wen_$_ANDNOT__A_Y ), .A3(fanout_net_6 ), .A4(_0213_ ), .ZN(wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ) );
NOR4_X1 _2893_ ( .A1(_0213_ ), .A2(_0167_ ), .A3(_0169_ ), .A4(_0168_ ), .ZN(wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ) );
AND3_X1 _2894_ ( .A1(_0163_ ), .A2(_0166_ ), .A3(\myicache.wen ), .ZN(wen_$_ANDNOT__A_Y_$_AND__B_Y ) );
NOR3_X1 _2895_ ( .A1(_0167_ ), .A2(_0168_ ), .A3(_0170_ ), .ZN(wen_$_ANDNOT__A_Y_$_AND__B_1_Y ) );
NOR3_X1 _2896_ ( .A1(_0167_ ), .A2(_0171_ ), .A3(_0170_ ), .ZN(wen_$_ANDNOT__A_Y_$_AND__B_2_Y ) );
NOR3_X1 _2897_ ( .A1(_0167_ ), .A2(_0170_ ), .A3(_0179_ ), .ZN(wen_$_ANDNOT__A_Y_$_AND__B_3_Y ) );
AND2_X1 _2898_ ( .A1(_0158_ ), .A2(rlast ), .ZN(_0885_ ) );
OAI221_X1 _2899_ ( .A(_0873_ ), .B1(\state [0] ), .B2(_0291_ ), .C1(_0885_ ), .C2(_0287_ ), .ZN(_0886_ ) );
AND4_X1 _2900_ ( .A1(_0177_ ), .A2(_0763_ ), .A3(_0869_ ), .A4(_0796_ ), .ZN(_0887_ ) );
AOI211_X1 _2901_ ( .A(_0886_ ), .B(_0887_ ), .C1(\state [0] ), .C2(_0884_ ), .ZN(wen_$_SDFFE_PP0P__Q_E ) );
CLKGATE_X1 _2902_ ( .CK(clock ), .E(wen_$_SDFFE_PP0P__Q_E ), .GCK(_1208_ ) );
CLKGATE_X1 _2903_ ( .CK(clock ), .E(tmp_offset_$_SDFFE_PP0P__Q_E ), .GCK(_1209_ ) );
CLKGATE_X1 _2904_ ( .CK(clock ), .E(pc_$_SDFFE_PP0P__Q_30_E ), .GCK(_1210_ ) );
CLKGATE_X1 _2905_ ( .CK(clock ), .E(readyFromIDU_$_AND__B_Y ), .GCK(_1211_ ) );
CLKGATE_X1 _2906_ ( .CK(clock ), .E(\myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_1212_ ) );
CLKGATE_X1 _2907_ ( .CK(clock ), .E(\myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_1213_ ) );
CLKGATE_X1 _2908_ ( .CK(clock ), .E(\myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_1214_ ) );
CLKGATE_X1 _2909_ ( .CK(clock ), .E(\myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_1215_ ) );
CLKGATE_X1 _2910_ ( .CK(clock ), .E(wen_$_ANDNOT__A_Y_$_AND__B_3_Y ), .GCK(_1216_ ) );
CLKGATE_X1 _2911_ ( .CK(clock ), .E(wen_$_ANDNOT__A_Y_$_AND__B_2_Y ), .GCK(_1217_ ) );
CLKGATE_X1 _2912_ ( .CK(clock ), .E(wen_$_ANDNOT__A_Y_$_AND__B_1_Y ), .GCK(_1218_ ) );
CLKGATE_X1 _2913_ ( .CK(clock ), .E(wen_$_ANDNOT__A_Y_$_AND__B_Y ), .GCK(_1219_ ) );
CLKGATE_X1 _2914_ ( .CK(clock ), .E(wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ), .GCK(_1220_ ) );
CLKGATE_X1 _2915_ ( .CK(clock ), .E(wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ), .GCK(_1221_ ) );
CLKGATE_X1 _2916_ ( .CK(clock ), .E(wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ), .GCK(_1222_ ) );
CLKGATE_X1 _2917_ ( .CK(clock ), .E(wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ), .GCK(_1223_ ) );
CLKGATE_X1 _2918_ ( .CK(clock ), .E(wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ), .GCK(_1224_ ) );
CLKGATE_X1 _2919_ ( .CK(clock ), .E(wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ), .GCK(_1225_ ) );
CLKGATE_X1 _2920_ ( .CK(clock ), .E(wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_1226_ ) );
CLKGATE_X1 _2921_ ( .CK(clock ), .E(wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ), .GCK(_1227_ ) );
CLKGATE_X1 _2922_ ( .CK(clock ), .E(rmem_quest_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y ), .GCK(_1228_ ) );
CLKGATE_X1 _2923_ ( .CK(clock ), .E(check_assert_$_DFFE_PP__Q_E ), .GCK(_1229_ ) );
LOGIC1_X1 _2924_ ( .Z(\arburst [0] ) );
LOGIC0_X1 _2925_ ( .Z(\araddr [0] ) );
DFF_X1 check_assert_$_DFFE_PP__Q ( .D(\state [1] ), .CK(_1229_ ), .Q(check_assert ), .QN(_1264_ ) );
DFF_X1 inst_$_DFFE_PP__Q ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ), .CK(_1228_ ), .Q(\inst [31] ), .QN(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_1 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ), .CK(_1228_ ), .Q(\inst [30] ), .QN(pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_10 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ), .CK(_1228_ ), .Q(\inst [21] ), .QN(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_11 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ), .CK(_1228_ ), .Q(\inst [20] ), .QN(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_12 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ), .CK(_1228_ ), .Q(\inst [19] ), .QN(pc_$_SDFFE_PP0P__Q_10_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_13 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ), .CK(_1228_ ), .Q(\inst [18] ), .QN(pc_$_SDFFE_PP0P__Q_12_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_14 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ), .CK(_1228_ ), .Q(\inst [17] ), .QN(pc_$_SDFFE_PP0P__Q_12_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ORNOT__Y_B_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_15 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ), .CK(_1228_ ), .Q(\inst [16] ), .QN(pc_$_SDFFE_PP0P__Q_14_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_16 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ), .CK(_1228_ ), .Q(\inst [15] ), .QN(pc_$_SDFFE_PP0P__Q_14_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_17 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ), .CK(_1228_ ), .Q(\inst [14] ), .QN(pc_$_SDFFE_PP0P__Q_16_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_18 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ), .CK(_1228_ ), .Q(\inst [13] ), .QN(pc_$_SDFFE_PP0P__Q_16_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_19 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ), .CK(_1228_ ), .Q(\inst [12] ), .QN(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_2 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ), .CK(_1228_ ), .Q(\inst [29] ), .QN(pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_20 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ), .CK(_1228_ ), .Q(\inst [11] ), .QN(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_21 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ), .CK(_1228_ ), .Q(\inst [10] ), .QN(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_22 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ), .CK(_1228_ ), .Q(\inst [9] ), .QN(pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_23 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ), .CK(_1228_ ), .Q(\inst [8] ), .QN(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_24 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ), .CK(_1228_ ), .Q(\inst [7] ), .QN(pc_$_SDFFE_PP0P__Q_18_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_25 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ), .CK(_1228_ ), .Q(\inst [6] ), .QN(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 inst_$_DFFE_PP__Q_26 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ), .CK(_1228_ ), .Q(\inst [5] ), .QN(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 inst_$_DFFE_PP__Q_27 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ), .CK(_1228_ ), .Q(\inst [4] ), .QN(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 inst_$_DFFE_PP__Q_28 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ), .CK(_1228_ ), .Q(\inst [3] ), .QN(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 inst_$_DFFE_PP__Q_29 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ), .CK(_1228_ ), .Q(\inst [2] ), .QN(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 inst_$_DFFE_PP__Q_3 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ), .CK(_1228_ ), .Q(\inst [28] ), .QN(pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_30 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ), .CK(_1228_ ), .Q(\inst [1] ), .QN(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 inst_$_DFFE_PP__Q_31 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ), .CK(_1228_ ), .Q(\inst [0] ), .QN(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 inst_$_DFFE_PP__Q_4 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ), .CK(_1228_ ), .Q(\inst [27] ), .QN(pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_5 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ), .CK(_1228_ ), .Q(\inst [26] ), .QN(pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_6 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ), .CK(_1228_ ), .Q(\inst [25] ), .QN(pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_7 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ), .CK(_1228_ ), .Q(\inst [24] ), .QN(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_8 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ), .CK(_1228_ ), .Q(\inst [23] ), .QN(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_A_$_OR__Y_B ) );
DFF_X1 inst_$_DFFE_PP__Q_9 ( .D(\pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__A_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ), .CK(_1228_ ), .Q(\inst [22] ), .QN(pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q ( .D(\rdata [19] ), .CK(_1227_ ), .Q(\myicache.data[0][19] ), .QN(_1265_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\rdata [18] ), .CK(_1227_ ), .Q(\myicache.data[0][18] ), .QN(_1266_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\rdata [9] ), .CK(_1227_ ), .Q(\myicache.data[0][9] ), .QN(_1267_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\rdata [8] ), .CK(_1227_ ), .Q(\myicache.data[0][8] ), .QN(_1268_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\rdata [7] ), .CK(_1227_ ), .Q(\myicache.data[0][7] ), .QN(_1269_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\rdata [6] ), .CK(_1227_ ), .Q(\myicache.data[0][6] ), .QN(_1270_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\rdata [5] ), .CK(_1227_ ), .Q(\myicache.data[0][5] ), .QN(_1271_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\rdata [4] ), .CK(_1227_ ), .Q(\myicache.data[0][4] ), .QN(_1272_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\rdata [3] ), .CK(_1227_ ), .Q(\myicache.data[0][3] ), .QN(_1273_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\rdata [2] ), .CK(_1227_ ), .Q(\myicache.data[0][2] ), .QN(_1274_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\rdata [1] ), .CK(_1227_ ), .Q(\myicache.data[0][1] ), .QN(_1275_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\rdata [0] ), .CK(_1227_ ), .Q(\myicache.data[0][0] ), .QN(_1276_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\rdata [17] ), .CK(_1227_ ), .Q(\myicache.data[0][17] ), .QN(_1277_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\rdata [31] ), .CK(_1227_ ), .Q(\myicache.data[0][31] ), .QN(_1278_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\rdata [30] ), .CK(_1227_ ), .Q(\myicache.data[0][30] ), .QN(_1279_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\rdata [29] ), .CK(_1227_ ), .Q(\myicache.data[0][29] ), .QN(_1280_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\rdata [28] ), .CK(_1227_ ), .Q(\myicache.data[0][28] ), .QN(_1281_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\rdata [27] ), .CK(_1227_ ), .Q(\myicache.data[0][27] ), .QN(_1282_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\rdata [26] ), .CK(_1227_ ), .Q(\myicache.data[0][26] ), .QN(_1283_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\rdata [25] ), .CK(_1227_ ), .Q(\myicache.data[0][25] ), .QN(_1284_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\rdata [24] ), .CK(_1227_ ), .Q(\myicache.data[0][24] ), .QN(_1285_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\rdata [23] ), .CK(_1227_ ), .Q(\myicache.data[0][23] ), .QN(_1286_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\rdata [22] ), .CK(_1227_ ), .Q(\myicache.data[0][22] ), .QN(_1287_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\rdata [16] ), .CK(_1227_ ), .Q(\myicache.data[0][16] ), .QN(_1288_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\rdata [21] ), .CK(_1227_ ), .Q(\myicache.data[0][21] ), .QN(_1289_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\rdata [20] ), .CK(_1227_ ), .Q(\myicache.data[0][20] ), .QN(_1290_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\rdata [15] ), .CK(_1227_ ), .Q(\myicache.data[0][15] ), .QN(_1291_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\rdata [14] ), .CK(_1227_ ), .Q(\myicache.data[0][14] ), .QN(_1292_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\rdata [13] ), .CK(_1227_ ), .Q(\myicache.data[0][13] ), .QN(_1293_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\rdata [12] ), .CK(_1227_ ), .Q(\myicache.data[0][12] ), .QN(_1294_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\rdata [11] ), .CK(_1227_ ), .Q(\myicache.data[0][11] ), .QN(_1295_ ) );
DFF_X1 \myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\rdata [10] ), .CK(_1227_ ), .Q(\myicache.data[0][10] ), .QN(_1296_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q ( .D(\rdata [31] ), .CK(_1226_ ), .Q(\myicache.data[1][31] ), .QN(_1297_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\rdata [30] ), .CK(_1226_ ), .Q(\myicache.data[1][30] ), .QN(_1298_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\rdata [21] ), .CK(_1226_ ), .Q(\myicache.data[1][21] ), .QN(_1299_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\rdata [20] ), .CK(_1226_ ), .Q(\myicache.data[1][20] ), .QN(_1300_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\rdata [19] ), .CK(_1226_ ), .Q(\myicache.data[1][19] ), .QN(_1301_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\rdata [18] ), .CK(_1226_ ), .Q(\myicache.data[1][18] ), .QN(_1302_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\rdata [17] ), .CK(_1226_ ), .Q(\myicache.data[1][17] ), .QN(_1303_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\rdata [16] ), .CK(_1226_ ), .Q(\myicache.data[1][16] ), .QN(_1304_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\rdata [15] ), .CK(_1226_ ), .Q(\myicache.data[1][15] ), .QN(_1305_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\rdata [14] ), .CK(_1226_ ), .Q(\myicache.data[1][14] ), .QN(_1306_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\rdata [13] ), .CK(_1226_ ), .Q(\myicache.data[1][13] ), .QN(_1307_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\rdata [12] ), .CK(_1226_ ), .Q(\myicache.data[1][12] ), .QN(_1308_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\rdata [29] ), .CK(_1226_ ), .Q(\myicache.data[1][29] ), .QN(_1309_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\rdata [11] ), .CK(_1226_ ), .Q(\myicache.data[1][11] ), .QN(_1310_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\rdata [10] ), .CK(_1226_ ), .Q(\myicache.data[1][10] ), .QN(_1311_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\rdata [9] ), .CK(_1226_ ), .Q(\myicache.data[1][9] ), .QN(_1312_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\rdata [8] ), .CK(_1226_ ), .Q(\myicache.data[1][8] ), .QN(_1313_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\rdata [7] ), .CK(_1226_ ), .Q(\myicache.data[1][7] ), .QN(_1314_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\rdata [6] ), .CK(_1226_ ), .Q(\myicache.data[1][6] ), .QN(_1315_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\rdata [5] ), .CK(_1226_ ), .Q(\myicache.data[1][5] ), .QN(_1316_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\rdata [4] ), .CK(_1226_ ), .Q(\myicache.data[1][4] ), .QN(_1317_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\rdata [3] ), .CK(_1226_ ), .Q(\myicache.data[1][3] ), .QN(_1318_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\rdata [2] ), .CK(_1226_ ), .Q(\myicache.data[1][2] ), .QN(_1319_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\rdata [28] ), .CK(_1226_ ), .Q(\myicache.data[1][28] ), .QN(_1320_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\rdata [1] ), .CK(_1226_ ), .Q(\myicache.data[1][1] ), .QN(_1321_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\rdata [0] ), .CK(_1226_ ), .Q(\myicache.data[1][0] ), .QN(_1322_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\rdata [27] ), .CK(_1226_ ), .Q(\myicache.data[1][27] ), .QN(_1323_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\rdata [26] ), .CK(_1226_ ), .Q(\myicache.data[1][26] ), .QN(_1324_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\rdata [25] ), .CK(_1226_ ), .Q(\myicache.data[1][25] ), .QN(_1325_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\rdata [24] ), .CK(_1226_ ), .Q(\myicache.data[1][24] ), .QN(_1326_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\rdata [23] ), .CK(_1226_ ), .Q(\myicache.data[1][23] ), .QN(_1327_ ) );
DFF_X1 \myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\rdata [22] ), .CK(_1226_ ), .Q(\myicache.data[1][22] ), .QN(_1328_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q ( .D(\rdata [31] ), .CK(_1225_ ), .Q(\myicache.data[2][31] ), .QN(_1329_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\rdata [30] ), .CK(_1225_ ), .Q(\myicache.data[2][30] ), .QN(_1330_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\rdata [21] ), .CK(_1225_ ), .Q(\myicache.data[2][21] ), .QN(_1331_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\rdata [20] ), .CK(_1225_ ), .Q(\myicache.data[2][20] ), .QN(_1332_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\rdata [19] ), .CK(_1225_ ), .Q(\myicache.data[2][19] ), .QN(_1333_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\rdata [18] ), .CK(_1225_ ), .Q(\myicache.data[2][18] ), .QN(_1334_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\rdata [17] ), .CK(_1225_ ), .Q(\myicache.data[2][17] ), .QN(_1335_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\rdata [16] ), .CK(_1225_ ), .Q(\myicache.data[2][16] ), .QN(_1336_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\rdata [15] ), .CK(_1225_ ), .Q(\myicache.data[2][15] ), .QN(_1337_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\rdata [14] ), .CK(_1225_ ), .Q(\myicache.data[2][14] ), .QN(_1338_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\rdata [13] ), .CK(_1225_ ), .Q(\myicache.data[2][13] ), .QN(_1339_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\rdata [12] ), .CK(_1225_ ), .Q(\myicache.data[2][12] ), .QN(_1340_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\rdata [29] ), .CK(_1225_ ), .Q(\myicache.data[2][29] ), .QN(_1341_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\rdata [11] ), .CK(_1225_ ), .Q(\myicache.data[2][11] ), .QN(_1342_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\rdata [10] ), .CK(_1225_ ), .Q(\myicache.data[2][10] ), .QN(_1343_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\rdata [9] ), .CK(_1225_ ), .Q(\myicache.data[2][9] ), .QN(_1344_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\rdata [8] ), .CK(_1225_ ), .Q(\myicache.data[2][8] ), .QN(_1345_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\rdata [7] ), .CK(_1225_ ), .Q(\myicache.data[2][7] ), .QN(_1346_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\rdata [6] ), .CK(_1225_ ), .Q(\myicache.data[2][6] ), .QN(_1347_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\rdata [5] ), .CK(_1225_ ), .Q(\myicache.data[2][5] ), .QN(_1348_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\rdata [4] ), .CK(_1225_ ), .Q(\myicache.data[2][4] ), .QN(_1349_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\rdata [3] ), .CK(_1225_ ), .Q(\myicache.data[2][3] ), .QN(_1350_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\rdata [2] ), .CK(_1225_ ), .Q(\myicache.data[2][2] ), .QN(_1351_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\rdata [28] ), .CK(_1225_ ), .Q(\myicache.data[2][28] ), .QN(_1352_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\rdata [1] ), .CK(_1225_ ), .Q(\myicache.data[2][1] ), .QN(_1353_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\rdata [0] ), .CK(_1225_ ), .Q(\myicache.data[2][0] ), .QN(_1354_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\rdata [27] ), .CK(_1225_ ), .Q(\myicache.data[2][27] ), .QN(_1355_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\rdata [26] ), .CK(_1225_ ), .Q(\myicache.data[2][26] ), .QN(_1356_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\rdata [25] ), .CK(_1225_ ), .Q(\myicache.data[2][25] ), .QN(_1357_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\rdata [24] ), .CK(_1225_ ), .Q(\myicache.data[2][24] ), .QN(_1358_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\rdata [23] ), .CK(_1225_ ), .Q(\myicache.data[2][23] ), .QN(_1359_ ) );
DFF_X1 \myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\rdata [22] ), .CK(_1225_ ), .Q(\myicache.data[2][22] ), .QN(_1360_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q ( .D(\rdata [31] ), .CK(_1224_ ), .Q(\myicache.data[3][31] ), .QN(_1361_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\rdata [30] ), .CK(_1224_ ), .Q(\myicache.data[3][30] ), .QN(_1362_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\rdata [21] ), .CK(_1224_ ), .Q(\myicache.data[3][21] ), .QN(_1363_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\rdata [20] ), .CK(_1224_ ), .Q(\myicache.data[3][20] ), .QN(_1364_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\rdata [19] ), .CK(_1224_ ), .Q(\myicache.data[3][19] ), .QN(_1365_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\rdata [18] ), .CK(_1224_ ), .Q(\myicache.data[3][18] ), .QN(_1366_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\rdata [17] ), .CK(_1224_ ), .Q(\myicache.data[3][17] ), .QN(_1367_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\rdata [16] ), .CK(_1224_ ), .Q(\myicache.data[3][16] ), .QN(_1368_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\rdata [15] ), .CK(_1224_ ), .Q(\myicache.data[3][15] ), .QN(_1369_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\rdata [14] ), .CK(_1224_ ), .Q(\myicache.data[3][14] ), .QN(_1370_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\rdata [13] ), .CK(_1224_ ), .Q(\myicache.data[3][13] ), .QN(_1371_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\rdata [12] ), .CK(_1224_ ), .Q(\myicache.data[3][12] ), .QN(_1372_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\rdata [29] ), .CK(_1224_ ), .Q(\myicache.data[3][29] ), .QN(_1373_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\rdata [11] ), .CK(_1224_ ), .Q(\myicache.data[3][11] ), .QN(_1374_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\rdata [10] ), .CK(_1224_ ), .Q(\myicache.data[3][10] ), .QN(_1375_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\rdata [9] ), .CK(_1224_ ), .Q(\myicache.data[3][9] ), .QN(_1376_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\rdata [8] ), .CK(_1224_ ), .Q(\myicache.data[3][8] ), .QN(_1377_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\rdata [7] ), .CK(_1224_ ), .Q(\myicache.data[3][7] ), .QN(_1378_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\rdata [6] ), .CK(_1224_ ), .Q(\myicache.data[3][6] ), .QN(_1379_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\rdata [5] ), .CK(_1224_ ), .Q(\myicache.data[3][5] ), .QN(_1380_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\rdata [4] ), .CK(_1224_ ), .Q(\myicache.data[3][4] ), .QN(_1381_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\rdata [3] ), .CK(_1224_ ), .Q(\myicache.data[3][3] ), .QN(_1382_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\rdata [2] ), .CK(_1224_ ), .Q(\myicache.data[3][2] ), .QN(_1383_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\rdata [28] ), .CK(_1224_ ), .Q(\myicache.data[3][28] ), .QN(_1384_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\rdata [1] ), .CK(_1224_ ), .Q(\myicache.data[3][1] ), .QN(_1385_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\rdata [0] ), .CK(_1224_ ), .Q(\myicache.data[3][0] ), .QN(_1386_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\rdata [27] ), .CK(_1224_ ), .Q(\myicache.data[3][27] ), .QN(_1387_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\rdata [26] ), .CK(_1224_ ), .Q(\myicache.data[3][26] ), .QN(_1388_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\rdata [25] ), .CK(_1224_ ), .Q(\myicache.data[3][25] ), .QN(_1389_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\rdata [24] ), .CK(_1224_ ), .Q(\myicache.data[3][24] ), .QN(_1390_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\rdata [23] ), .CK(_1224_ ), .Q(\myicache.data[3][23] ), .QN(_1391_ ) );
DFF_X1 \myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\rdata [22] ), .CK(_1224_ ), .Q(\myicache.data[3][22] ), .QN(_1392_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q ( .D(\rdata [31] ), .CK(_1223_ ), .Q(\myicache.data[4][31] ), .QN(_1393_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_1 ( .D(\rdata [30] ), .CK(_1223_ ), .Q(\myicache.data[4][30] ), .QN(_1394_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_10 ( .D(\rdata [21] ), .CK(_1223_ ), .Q(\myicache.data[4][21] ), .QN(_1395_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_11 ( .D(\rdata [20] ), .CK(_1223_ ), .Q(\myicache.data[4][20] ), .QN(_1396_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_12 ( .D(\rdata [19] ), .CK(_1223_ ), .Q(\myicache.data[4][19] ), .QN(_1397_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_13 ( .D(\rdata [18] ), .CK(_1223_ ), .Q(\myicache.data[4][18] ), .QN(_1398_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_14 ( .D(\rdata [17] ), .CK(_1223_ ), .Q(\myicache.data[4][17] ), .QN(_1399_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_15 ( .D(\rdata [16] ), .CK(_1223_ ), .Q(\myicache.data[4][16] ), .QN(_1400_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_16 ( .D(\rdata [15] ), .CK(_1223_ ), .Q(\myicache.data[4][15] ), .QN(_1401_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_17 ( .D(\rdata [14] ), .CK(_1223_ ), .Q(\myicache.data[4][14] ), .QN(_1402_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_18 ( .D(\rdata [13] ), .CK(_1223_ ), .Q(\myicache.data[4][13] ), .QN(_1403_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_19 ( .D(\rdata [12] ), .CK(_1223_ ), .Q(\myicache.data[4][12] ), .QN(_1404_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_2 ( .D(\rdata [29] ), .CK(_1223_ ), .Q(\myicache.data[4][29] ), .QN(_1405_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_20 ( .D(\rdata [11] ), .CK(_1223_ ), .Q(\myicache.data[4][11] ), .QN(_1406_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_21 ( .D(\rdata [10] ), .CK(_1223_ ), .Q(\myicache.data[4][10] ), .QN(_1407_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_22 ( .D(\rdata [9] ), .CK(_1223_ ), .Q(\myicache.data[4][9] ), .QN(_1408_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_23 ( .D(\rdata [8] ), .CK(_1223_ ), .Q(\myicache.data[4][8] ), .QN(_1409_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_24 ( .D(\rdata [7] ), .CK(_1223_ ), .Q(\myicache.data[4][7] ), .QN(_1410_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_25 ( .D(\rdata [6] ), .CK(_1223_ ), .Q(\myicache.data[4][6] ), .QN(_1411_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_26 ( .D(\rdata [5] ), .CK(_1223_ ), .Q(\myicache.data[4][5] ), .QN(_1412_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_27 ( .D(\rdata [4] ), .CK(_1223_ ), .Q(\myicache.data[4][4] ), .QN(_1413_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_28 ( .D(\rdata [3] ), .CK(_1223_ ), .Q(\myicache.data[4][3] ), .QN(_1414_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_29 ( .D(\rdata [2] ), .CK(_1223_ ), .Q(\myicache.data[4][2] ), .QN(_1415_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_3 ( .D(\rdata [28] ), .CK(_1223_ ), .Q(\myicache.data[4][28] ), .QN(_1416_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_30 ( .D(\rdata [1] ), .CK(_1223_ ), .Q(\myicache.data[4][1] ), .QN(_1417_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_31 ( .D(\rdata [0] ), .CK(_1223_ ), .Q(\myicache.data[4][0] ), .QN(_1418_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_4 ( .D(\rdata [27] ), .CK(_1223_ ), .Q(\myicache.data[4][27] ), .QN(_1419_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_5 ( .D(\rdata [26] ), .CK(_1223_ ), .Q(\myicache.data[4][26] ), .QN(_1420_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_6 ( .D(\rdata [25] ), .CK(_1223_ ), .Q(\myicache.data[4][25] ), .QN(_1421_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_7 ( .D(\rdata [24] ), .CK(_1223_ ), .Q(\myicache.data[4][24] ), .QN(_1422_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_8 ( .D(\rdata [23] ), .CK(_1223_ ), .Q(\myicache.data[4][23] ), .QN(_1423_ ) );
DFF_X1 \myicache.data[4]_$_DFFE_PP__Q_9 ( .D(\rdata [22] ), .CK(_1223_ ), .Q(\myicache.data[4][22] ), .QN(_1424_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q ( .D(\rdata [31] ), .CK(_1222_ ), .Q(\myicache.data[5][31] ), .QN(_1425_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_1 ( .D(\rdata [30] ), .CK(_1222_ ), .Q(\myicache.data[5][30] ), .QN(_1426_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_10 ( .D(\rdata [21] ), .CK(_1222_ ), .Q(\myicache.data[5][21] ), .QN(_1427_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_11 ( .D(\rdata [20] ), .CK(_1222_ ), .Q(\myicache.data[5][20] ), .QN(_1428_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_12 ( .D(\rdata [19] ), .CK(_1222_ ), .Q(\myicache.data[5][19] ), .QN(_1429_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_13 ( .D(\rdata [18] ), .CK(_1222_ ), .Q(\myicache.data[5][18] ), .QN(_1430_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_14 ( .D(\rdata [17] ), .CK(_1222_ ), .Q(\myicache.data[5][17] ), .QN(_1431_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_15 ( .D(\rdata [16] ), .CK(_1222_ ), .Q(\myicache.data[5][16] ), .QN(_1432_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_16 ( .D(\rdata [15] ), .CK(_1222_ ), .Q(\myicache.data[5][15] ), .QN(_1433_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_17 ( .D(\rdata [14] ), .CK(_1222_ ), .Q(\myicache.data[5][14] ), .QN(_1434_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_18 ( .D(\rdata [13] ), .CK(_1222_ ), .Q(\myicache.data[5][13] ), .QN(_1435_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_19 ( .D(\rdata [12] ), .CK(_1222_ ), .Q(\myicache.data[5][12] ), .QN(_1436_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_2 ( .D(\rdata [29] ), .CK(_1222_ ), .Q(\myicache.data[5][29] ), .QN(_1437_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_20 ( .D(\rdata [11] ), .CK(_1222_ ), .Q(\myicache.data[5][11] ), .QN(_1438_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_21 ( .D(\rdata [10] ), .CK(_1222_ ), .Q(\myicache.data[5][10] ), .QN(_1439_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_22 ( .D(\rdata [9] ), .CK(_1222_ ), .Q(\myicache.data[5][9] ), .QN(_1440_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_23 ( .D(\rdata [8] ), .CK(_1222_ ), .Q(\myicache.data[5][8] ), .QN(_1441_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_24 ( .D(\rdata [7] ), .CK(_1222_ ), .Q(\myicache.data[5][7] ), .QN(_1442_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_25 ( .D(\rdata [6] ), .CK(_1222_ ), .Q(\myicache.data[5][6] ), .QN(_1443_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_26 ( .D(\rdata [5] ), .CK(_1222_ ), .Q(\myicache.data[5][5] ), .QN(_1444_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_27 ( .D(\rdata [4] ), .CK(_1222_ ), .Q(\myicache.data[5][4] ), .QN(_1445_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_28 ( .D(\rdata [3] ), .CK(_1222_ ), .Q(\myicache.data[5][3] ), .QN(_1446_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_29 ( .D(\rdata [2] ), .CK(_1222_ ), .Q(\myicache.data[5][2] ), .QN(_1447_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_3 ( .D(\rdata [28] ), .CK(_1222_ ), .Q(\myicache.data[5][28] ), .QN(_1448_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_30 ( .D(\rdata [1] ), .CK(_1222_ ), .Q(\myicache.data[5][1] ), .QN(_1449_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_31 ( .D(\rdata [0] ), .CK(_1222_ ), .Q(\myicache.data[5][0] ), .QN(_1450_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_4 ( .D(\rdata [27] ), .CK(_1222_ ), .Q(\myicache.data[5][27] ), .QN(_1451_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_5 ( .D(\rdata [26] ), .CK(_1222_ ), .Q(\myicache.data[5][26] ), .QN(_1452_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_6 ( .D(\rdata [25] ), .CK(_1222_ ), .Q(\myicache.data[5][25] ), .QN(_1453_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_7 ( .D(\rdata [24] ), .CK(_1222_ ), .Q(\myicache.data[5][24] ), .QN(_1454_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_8 ( .D(\rdata [23] ), .CK(_1222_ ), .Q(\myicache.data[5][23] ), .QN(_1455_ ) );
DFF_X1 \myicache.data[5]_$_DFFE_PP__Q_9 ( .D(\rdata [22] ), .CK(_1222_ ), .Q(\myicache.data[5][22] ), .QN(_1456_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q ( .D(\rdata [31] ), .CK(_1221_ ), .Q(\myicache.data[6][31] ), .QN(_1457_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_1 ( .D(\rdata [30] ), .CK(_1221_ ), .Q(\myicache.data[6][30] ), .QN(_1458_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_10 ( .D(\rdata [21] ), .CK(_1221_ ), .Q(\myicache.data[6][21] ), .QN(_1459_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_11 ( .D(\rdata [20] ), .CK(_1221_ ), .Q(\myicache.data[6][20] ), .QN(_1460_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_12 ( .D(\rdata [19] ), .CK(_1221_ ), .Q(\myicache.data[6][19] ), .QN(_1461_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_13 ( .D(\rdata [18] ), .CK(_1221_ ), .Q(\myicache.data[6][18] ), .QN(_1462_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_14 ( .D(\rdata [17] ), .CK(_1221_ ), .Q(\myicache.data[6][17] ), .QN(_1463_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_15 ( .D(\rdata [16] ), .CK(_1221_ ), .Q(\myicache.data[6][16] ), .QN(_1464_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_16 ( .D(\rdata [15] ), .CK(_1221_ ), .Q(\myicache.data[6][15] ), .QN(_1465_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_17 ( .D(\rdata [14] ), .CK(_1221_ ), .Q(\myicache.data[6][14] ), .QN(_1466_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_18 ( .D(\rdata [13] ), .CK(_1221_ ), .Q(\myicache.data[6][13] ), .QN(_1467_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_19 ( .D(\rdata [12] ), .CK(_1221_ ), .Q(\myicache.data[6][12] ), .QN(_1468_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_2 ( .D(\rdata [29] ), .CK(_1221_ ), .Q(\myicache.data[6][29] ), .QN(_1469_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_20 ( .D(\rdata [11] ), .CK(_1221_ ), .Q(\myicache.data[6][11] ), .QN(_1470_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_21 ( .D(\rdata [10] ), .CK(_1221_ ), .Q(\myicache.data[6][10] ), .QN(_1471_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_22 ( .D(\rdata [9] ), .CK(_1221_ ), .Q(\myicache.data[6][9] ), .QN(_1472_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_23 ( .D(\rdata [8] ), .CK(_1221_ ), .Q(\myicache.data[6][8] ), .QN(_1473_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_24 ( .D(\rdata [7] ), .CK(_1221_ ), .Q(\myicache.data[6][7] ), .QN(_1474_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_25 ( .D(\rdata [6] ), .CK(_1221_ ), .Q(\myicache.data[6][6] ), .QN(_1475_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_26 ( .D(\rdata [5] ), .CK(_1221_ ), .Q(\myicache.data[6][5] ), .QN(_1476_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_27 ( .D(\rdata [4] ), .CK(_1221_ ), .Q(\myicache.data[6][4] ), .QN(_1477_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_28 ( .D(\rdata [3] ), .CK(_1221_ ), .Q(\myicache.data[6][3] ), .QN(_1478_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_29 ( .D(\rdata [2] ), .CK(_1221_ ), .Q(\myicache.data[6][2] ), .QN(_1479_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_3 ( .D(\rdata [28] ), .CK(_1221_ ), .Q(\myicache.data[6][28] ), .QN(_1480_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_30 ( .D(\rdata [1] ), .CK(_1221_ ), .Q(\myicache.data[6][1] ), .QN(_1481_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_31 ( .D(\rdata [0] ), .CK(_1221_ ), .Q(\myicache.data[6][0] ), .QN(_1482_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_4 ( .D(\rdata [27] ), .CK(_1221_ ), .Q(\myicache.data[6][27] ), .QN(_1483_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_5 ( .D(\rdata [26] ), .CK(_1221_ ), .Q(\myicache.data[6][26] ), .QN(_1484_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_6 ( .D(\rdata [25] ), .CK(_1221_ ), .Q(\myicache.data[6][25] ), .QN(_1485_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_7 ( .D(\rdata [24] ), .CK(_1221_ ), .Q(\myicache.data[6][24] ), .QN(_1486_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_8 ( .D(\rdata [23] ), .CK(_1221_ ), .Q(\myicache.data[6][23] ), .QN(_1487_ ) );
DFF_X1 \myicache.data[6]_$_DFFE_PP__Q_9 ( .D(\rdata [22] ), .CK(_1221_ ), .Q(\myicache.data[6][22] ), .QN(_1488_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q ( .D(\rdata [31] ), .CK(_1220_ ), .Q(\myicache.data[7][31] ), .QN(_1489_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_1 ( .D(\rdata [30] ), .CK(_1220_ ), .Q(\myicache.data[7][30] ), .QN(_1490_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_10 ( .D(\rdata [21] ), .CK(_1220_ ), .Q(\myicache.data[7][21] ), .QN(_1491_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_11 ( .D(\rdata [20] ), .CK(_1220_ ), .Q(\myicache.data[7][20] ), .QN(_1492_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_12 ( .D(\rdata [19] ), .CK(_1220_ ), .Q(\myicache.data[7][19] ), .QN(_1493_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_13 ( .D(\rdata [18] ), .CK(_1220_ ), .Q(\myicache.data[7][18] ), .QN(_1494_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_14 ( .D(\rdata [17] ), .CK(_1220_ ), .Q(\myicache.data[7][17] ), .QN(_1495_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_15 ( .D(\rdata [16] ), .CK(_1220_ ), .Q(\myicache.data[7][16] ), .QN(_1496_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_16 ( .D(\rdata [15] ), .CK(_1220_ ), .Q(\myicache.data[7][15] ), .QN(_1497_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_17 ( .D(\rdata [14] ), .CK(_1220_ ), .Q(\myicache.data[7][14] ), .QN(_1498_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_18 ( .D(\rdata [13] ), .CK(_1220_ ), .Q(\myicache.data[7][13] ), .QN(_1499_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_19 ( .D(\rdata [12] ), .CK(_1220_ ), .Q(\myicache.data[7][12] ), .QN(_1500_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_2 ( .D(\rdata [29] ), .CK(_1220_ ), .Q(\myicache.data[7][29] ), .QN(_1501_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_20 ( .D(\rdata [11] ), .CK(_1220_ ), .Q(\myicache.data[7][11] ), .QN(_1502_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_21 ( .D(\rdata [10] ), .CK(_1220_ ), .Q(\myicache.data[7][10] ), .QN(_1503_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_22 ( .D(\rdata [9] ), .CK(_1220_ ), .Q(\myicache.data[7][9] ), .QN(_1504_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_23 ( .D(\rdata [8] ), .CK(_1220_ ), .Q(\myicache.data[7][8] ), .QN(_1505_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_24 ( .D(\rdata [7] ), .CK(_1220_ ), .Q(\myicache.data[7][7] ), .QN(_1506_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_25 ( .D(\rdata [6] ), .CK(_1220_ ), .Q(\myicache.data[7][6] ), .QN(_1507_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_26 ( .D(\rdata [5] ), .CK(_1220_ ), .Q(\myicache.data[7][5] ), .QN(_1508_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_27 ( .D(\rdata [4] ), .CK(_1220_ ), .Q(\myicache.data[7][4] ), .QN(_1509_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_28 ( .D(\rdata [3] ), .CK(_1220_ ), .Q(\myicache.data[7][3] ), .QN(_1510_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_29 ( .D(\rdata [2] ), .CK(_1220_ ), .Q(\myicache.data[7][2] ), .QN(_1511_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_3 ( .D(\rdata [28] ), .CK(_1220_ ), .Q(\myicache.data[7][28] ), .QN(_1512_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_30 ( .D(\rdata [1] ), .CK(_1220_ ), .Q(\myicache.data[7][1] ), .QN(_1513_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_31 ( .D(\rdata [0] ), .CK(_1220_ ), .Q(\myicache.data[7][0] ), .QN(_1514_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_4 ( .D(\rdata [27] ), .CK(_1220_ ), .Q(\myicache.data[7][27] ), .QN(_1515_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_5 ( .D(\rdata [26] ), .CK(_1220_ ), .Q(\myicache.data[7][26] ), .QN(_1516_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_6 ( .D(\rdata [25] ), .CK(_1220_ ), .Q(\myicache.data[7][25] ), .QN(_1517_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_7 ( .D(\rdata [24] ), .CK(_1220_ ), .Q(\myicache.data[7][24] ), .QN(_1518_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_8 ( .D(\rdata [23] ), .CK(_1220_ ), .Q(\myicache.data[7][23] ), .QN(_1519_ ) );
DFF_X1 \myicache.data[7]_$_DFFE_PP__Q_9 ( .D(\rdata [22] ), .CK(_1220_ ), .Q(\myicache.data[7][22] ), .QN(_1520_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q ( .D(\araddr [31] ), .CK(_1219_ ), .Q(\myicache.tag[0][26] ), .QN(_1521_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\araddr [30] ), .CK(_1219_ ), .Q(\myicache.tag[0][25] ), .QN(_1522_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\araddr [21] ), .CK(_1219_ ), .Q(\myicache.tag[0][16] ), .QN(_1523_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\araddr [20] ), .CK(_1219_ ), .Q(\myicache.tag[0][15] ), .QN(_1524_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\araddr [19] ), .CK(_1219_ ), .Q(\myicache.tag[0][14] ), .QN(_1525_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\araddr [18] ), .CK(_1219_ ), .Q(\myicache.tag[0][13] ), .QN(_1526_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\araddr [17] ), .CK(_1219_ ), .Q(\myicache.tag[0][12] ), .QN(_1527_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\araddr [16] ), .CK(_1219_ ), .Q(\myicache.tag[0][11] ), .QN(_1528_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\araddr [15] ), .CK(_1219_ ), .Q(\myicache.tag[0][10] ), .QN(_1529_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\araddr [14] ), .CK(_1219_ ), .Q(\myicache.tag[0][9] ), .QN(_1530_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\araddr [13] ), .CK(_1219_ ), .Q(\myicache.tag[0][8] ), .QN(_1531_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\araddr [12] ), .CK(_1219_ ), .Q(\myicache.tag[0][7] ), .QN(_1532_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\araddr [29] ), .CK(_1219_ ), .Q(\myicache.tag[0][24] ), .QN(_1533_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\araddr [11] ), .CK(_1219_ ), .Q(\myicache.tag[0][6] ), .QN(_1534_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\araddr [10] ), .CK(_1219_ ), .Q(\myicache.tag[0][5] ), .QN(_1535_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\araddr [9] ), .CK(_1219_ ), .Q(\myicache.tag[0][4] ), .QN(_1536_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\araddr [8] ), .CK(_1219_ ), .Q(\myicache.tag[0][3] ), .QN(_1537_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\araddr [7] ), .CK(_1219_ ), .Q(\myicache.tag[0][2] ), .QN(_1538_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\araddr [6] ), .CK(_1219_ ), .Q(\myicache.tag[0][1] ), .QN(_1539_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\araddr [5] ), .CK(_1219_ ), .Q(\myicache.tag[0][0] ), .QN(_1540_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\araddr [28] ), .CK(_1219_ ), .Q(\myicache.tag[0][23] ), .QN(_1541_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\araddr [27] ), .CK(_1219_ ), .Q(\myicache.tag[0][22] ), .QN(_1542_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\araddr [26] ), .CK(_1219_ ), .Q(\myicache.tag[0][21] ), .QN(_1543_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\araddr [25] ), .CK(_1219_ ), .Q(\myicache.tag[0][20] ), .QN(_1544_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\araddr [24] ), .CK(_1219_ ), .Q(\myicache.tag[0][19] ), .QN(_1545_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\araddr [23] ), .CK(_1219_ ), .Q(\myicache.tag[0][18] ), .QN(_1546_ ) );
DFF_X1 \myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\araddr [22] ), .CK(_1219_ ), .Q(\myicache.tag[0][17] ), .QN(_1547_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q ( .D(\araddr [31] ), .CK(_1218_ ), .Q(\myicache.tag[1][26] ), .QN(_1548_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\araddr [30] ), .CK(_1218_ ), .Q(\myicache.tag[1][25] ), .QN(_1549_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\araddr [21] ), .CK(_1218_ ), .Q(\myicache.tag[1][16] ), .QN(_1550_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\araddr [20] ), .CK(_1218_ ), .Q(\myicache.tag[1][15] ), .QN(_1551_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\araddr [19] ), .CK(_1218_ ), .Q(\myicache.tag[1][14] ), .QN(_1552_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\araddr [18] ), .CK(_1218_ ), .Q(\myicache.tag[1][13] ), .QN(_1553_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\araddr [17] ), .CK(_1218_ ), .Q(\myicache.tag[1][12] ), .QN(_1554_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\araddr [16] ), .CK(_1218_ ), .Q(\myicache.tag[1][11] ), .QN(_1555_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\araddr [15] ), .CK(_1218_ ), .Q(\myicache.tag[1][10] ), .QN(_1556_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\araddr [14] ), .CK(_1218_ ), .Q(\myicache.tag[1][9] ), .QN(_1557_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\araddr [13] ), .CK(_1218_ ), .Q(\myicache.tag[1][8] ), .QN(_1558_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\araddr [12] ), .CK(_1218_ ), .Q(\myicache.tag[1][7] ), .QN(_1559_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\araddr [29] ), .CK(_1218_ ), .Q(\myicache.tag[1][24] ), .QN(_1560_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\araddr [11] ), .CK(_1218_ ), .Q(\myicache.tag[1][6] ), .QN(_1561_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\araddr [10] ), .CK(_1218_ ), .Q(\myicache.tag[1][5] ), .QN(_1562_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\araddr [9] ), .CK(_1218_ ), .Q(\myicache.tag[1][4] ), .QN(_1563_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\araddr [8] ), .CK(_1218_ ), .Q(\myicache.tag[1][3] ), .QN(_1564_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\araddr [7] ), .CK(_1218_ ), .Q(\myicache.tag[1][2] ), .QN(_1565_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\araddr [6] ), .CK(_1218_ ), .Q(\myicache.tag[1][1] ), .QN(_1566_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\araddr [5] ), .CK(_1218_ ), .Q(\myicache.tag[1][0] ), .QN(_1567_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\araddr [28] ), .CK(_1218_ ), .Q(\myicache.tag[1][23] ), .QN(_1568_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\araddr [27] ), .CK(_1218_ ), .Q(\myicache.tag[1][22] ), .QN(_1569_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\araddr [26] ), .CK(_1218_ ), .Q(\myicache.tag[1][21] ), .QN(_1570_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\araddr [25] ), .CK(_1218_ ), .Q(\myicache.tag[1][20] ), .QN(_1571_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\araddr [24] ), .CK(_1218_ ), .Q(\myicache.tag[1][19] ), .QN(_1572_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\araddr [23] ), .CK(_1218_ ), .Q(\myicache.tag[1][18] ), .QN(_1573_ ) );
DFF_X1 \myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\araddr [22] ), .CK(_1218_ ), .Q(\myicache.tag[1][17] ), .QN(_1574_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q ( .D(\araddr [31] ), .CK(_1217_ ), .Q(\myicache.tag[2][26] ), .QN(_1575_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\araddr [30] ), .CK(_1217_ ), .Q(\myicache.tag[2][25] ), .QN(_1576_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\araddr [21] ), .CK(_1217_ ), .Q(\myicache.tag[2][16] ), .QN(_1577_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\araddr [20] ), .CK(_1217_ ), .Q(\myicache.tag[2][15] ), .QN(_1578_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\araddr [19] ), .CK(_1217_ ), .Q(\myicache.tag[2][14] ), .QN(_1579_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\araddr [18] ), .CK(_1217_ ), .Q(\myicache.tag[2][13] ), .QN(_1580_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\araddr [17] ), .CK(_1217_ ), .Q(\myicache.tag[2][12] ), .QN(_1581_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\araddr [16] ), .CK(_1217_ ), .Q(\myicache.tag[2][11] ), .QN(_1582_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\araddr [15] ), .CK(_1217_ ), .Q(\myicache.tag[2][10] ), .QN(_1583_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\araddr [14] ), .CK(_1217_ ), .Q(\myicache.tag[2][9] ), .QN(_1584_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\araddr [13] ), .CK(_1217_ ), .Q(\myicache.tag[2][8] ), .QN(_1585_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\araddr [12] ), .CK(_1217_ ), .Q(\myicache.tag[2][7] ), .QN(_1586_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\araddr [29] ), .CK(_1217_ ), .Q(\myicache.tag[2][24] ), .QN(_1587_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\araddr [11] ), .CK(_1217_ ), .Q(\myicache.tag[2][6] ), .QN(_1588_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\araddr [10] ), .CK(_1217_ ), .Q(\myicache.tag[2][5] ), .QN(_1589_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\araddr [9] ), .CK(_1217_ ), .Q(\myicache.tag[2][4] ), .QN(_1590_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\araddr [8] ), .CK(_1217_ ), .Q(\myicache.tag[2][3] ), .QN(_1591_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\araddr [7] ), .CK(_1217_ ), .Q(\myicache.tag[2][2] ), .QN(_1592_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\araddr [6] ), .CK(_1217_ ), .Q(\myicache.tag[2][1] ), .QN(_1593_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\araddr [5] ), .CK(_1217_ ), .Q(\myicache.tag[2][0] ), .QN(_1594_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\araddr [28] ), .CK(_1217_ ), .Q(\myicache.tag[2][23] ), .QN(_1595_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\araddr [27] ), .CK(_1217_ ), .Q(\myicache.tag[2][22] ), .QN(_1596_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\araddr [26] ), .CK(_1217_ ), .Q(\myicache.tag[2][21] ), .QN(_1597_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\araddr [25] ), .CK(_1217_ ), .Q(\myicache.tag[2][20] ), .QN(_1598_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\araddr [24] ), .CK(_1217_ ), .Q(\myicache.tag[2][19] ), .QN(_1599_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\araddr [23] ), .CK(_1217_ ), .Q(\myicache.tag[2][18] ), .QN(_1600_ ) );
DFF_X1 \myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\araddr [22] ), .CK(_1217_ ), .Q(\myicache.tag[2][17] ), .QN(_1601_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q ( .D(\araddr [31] ), .CK(_1216_ ), .Q(\myicache.tag[3][26] ), .QN(_1602_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\araddr [30] ), .CK(_1216_ ), .Q(\myicache.tag[3][25] ), .QN(_1603_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\araddr [21] ), .CK(_1216_ ), .Q(\myicache.tag[3][16] ), .QN(_1604_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\araddr [20] ), .CK(_1216_ ), .Q(\myicache.tag[3][15] ), .QN(_1605_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\araddr [19] ), .CK(_1216_ ), .Q(\myicache.tag[3][14] ), .QN(_1606_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\araddr [18] ), .CK(_1216_ ), .Q(\myicache.tag[3][13] ), .QN(_1607_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\araddr [17] ), .CK(_1216_ ), .Q(\myicache.tag[3][12] ), .QN(_1608_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\araddr [16] ), .CK(_1216_ ), .Q(\myicache.tag[3][11] ), .QN(_1609_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\araddr [15] ), .CK(_1216_ ), .Q(\myicache.tag[3][10] ), .QN(_1610_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\araddr [14] ), .CK(_1216_ ), .Q(\myicache.tag[3][9] ), .QN(_1611_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\araddr [13] ), .CK(_1216_ ), .Q(\myicache.tag[3][8] ), .QN(_1612_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\araddr [12] ), .CK(_1216_ ), .Q(\myicache.tag[3][7] ), .QN(_1613_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\araddr [29] ), .CK(_1216_ ), .Q(\myicache.tag[3][24] ), .QN(_1614_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\araddr [11] ), .CK(_1216_ ), .Q(\myicache.tag[3][6] ), .QN(_1615_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\araddr [10] ), .CK(_1216_ ), .Q(\myicache.tag[3][5] ), .QN(_1616_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\araddr [9] ), .CK(_1216_ ), .Q(\myicache.tag[3][4] ), .QN(_1617_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\araddr [8] ), .CK(_1216_ ), .Q(\myicache.tag[3][3] ), .QN(_1618_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\araddr [7] ), .CK(_1216_ ), .Q(\myicache.tag[3][2] ), .QN(_1619_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\araddr [6] ), .CK(_1216_ ), .Q(\myicache.tag[3][1] ), .QN(_1620_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\araddr [5] ), .CK(_1216_ ), .Q(\myicache.tag[3][0] ), .QN(_1621_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\araddr [28] ), .CK(_1216_ ), .Q(\myicache.tag[3][23] ), .QN(_1622_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\araddr [27] ), .CK(_1216_ ), .Q(\myicache.tag[3][22] ), .QN(_1623_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\araddr [26] ), .CK(_1216_ ), .Q(\myicache.tag[3][21] ), .QN(_1624_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\araddr [25] ), .CK(_1216_ ), .Q(\myicache.tag[3][20] ), .QN(_1625_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\araddr [24] ), .CK(_1216_ ), .Q(\myicache.tag[3][19] ), .QN(_1626_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\araddr [23] ), .CK(_1216_ ), .Q(\myicache.tag[3][18] ), .QN(_1627_ ) );
DFF_X1 \myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\araddr [22] ), .CK(_1216_ ), .Q(\myicache.tag[3][17] ), .QN(_1263_ ) );
DFF_X1 \myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_0000_ ), .CK(_1215_ ), .Q(\myicache.valid [0] ), .QN(_1262_ ) );
DFF_X1 \myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_0001_ ), .CK(_1214_ ), .Q(\myicache.valid [1] ), .QN(_1261_ ) );
DFF_X1 \myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_0002_ ), .CK(_1213_ ), .Q(\myicache.valid [2] ), .QN(_1628_ ) );
DFF_X1 \myicache.valid[3]_$_DFFE_PP__Q ( .D(wen_$_ANDNOT__A_Y ), .CK(_1212_ ), .Q(\myicache.valid [3] ), .QN(_1260_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q ( .D(_0003_ ), .CK(_1211_ ), .Q(\araddr [30] ), .QN(_1259_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_1 ( .D(_0004_ ), .CK(_1211_ ), .Q(\araddr [29] ), .QN(_1258_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_10 ( .D(_0005_ ), .CK(_1211_ ), .Q(\araddr [20] ), .QN(_1257_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_11 ( .D(_0006_ ), .CK(_1211_ ), .Q(\araddr [19] ), .QN(_1256_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_12 ( .D(_0007_ ), .CK(_1211_ ), .Q(\araddr [18] ), .QN(pc_$_SDFFE_PP0P__Q_12_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_B ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_13 ( .D(_0008_ ), .CK(_1211_ ), .Q(\araddr [17] ), .QN(_1255_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_14 ( .D(_0009_ ), .CK(_1211_ ), .Q(\araddr [16] ), .QN(_1254_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_15 ( .D(_0010_ ), .CK(_1211_ ), .Q(\araddr [15] ), .QN(_1253_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_16 ( .D(_0011_ ), .CK(_1211_ ), .Q(\araddr [14] ), .QN(_1252_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_17 ( .D(_0012_ ), .CK(_1211_ ), .Q(\araddr [13] ), .QN(_1251_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_18 ( .D(_0013_ ), .CK(_1211_ ), .Q(\araddr [12] ), .QN(_1250_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_19 ( .D(_0014_ ), .CK(_1211_ ), .Q(\araddr [11] ), .QN(_1249_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_2 ( .D(_0015_ ), .CK(_1211_ ), .Q(\araddr [28] ), .QN(_1248_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_20 ( .D(_0016_ ), .CK(_1211_ ), .Q(\araddr [10] ), .QN(_1247_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_21 ( .D(_0017_ ), .CK(_1211_ ), .Q(\araddr [9] ), .QN(_1246_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_22 ( .D(_0018_ ), .CK(_1211_ ), .Q(\araddr [8] ), .QN(_1245_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_23 ( .D(_0019_ ), .CK(_1211_ ), .Q(\araddr [7] ), .QN(_1244_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_24 ( .D(_0020_ ), .CK(_1211_ ), .Q(\araddr [6] ), .QN(_1243_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_25 ( .D(_0021_ ), .CK(_1211_ ), .Q(\araddr [5] ), .QN(pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_26 ( .D(_0022_ ), .CK(_1211_ ), .Q(fanout_net_6 ), .QN(_1242_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_26_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_0024_ ), .CK(clock ), .Q(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_1241_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_27 ( .D(_0023_ ), .CK(_1211_ ), .Q(fanout_net_2 ), .QN(pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_0026_ ), .CK(clock ), .Q(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_1239_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_28 ( .D(_0025_ ), .CK(_1211_ ), .Q(\pc [2] ), .QN(_1240_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_29 ( .D(_0027_ ), .CK(_1211_ ), .Q(\pc [1] ), .QN(pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_3 ( .D(_0028_ ), .CK(_1211_ ), .Q(\araddr [27] ), .QN(_1238_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_30 ( .D(_0029_ ), .CK(_1210_ ), .Q(\pc [0] ), .QN(tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_4 ( .D(_0030_ ), .CK(_1211_ ), .Q(\araddr [26] ), .QN(_1237_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_5 ( .D(_0031_ ), .CK(_1211_ ), .Q(\araddr [25] ), .QN(_1236_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_6 ( .D(_0032_ ), .CK(_1211_ ), .Q(\araddr [24] ), .QN(_1235_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_7 ( .D(_0033_ ), .CK(_1211_ ), .Q(\araddr [23] ), .QN(_1234_ ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_8 ( .D(_0034_ ), .CK(_1211_ ), .Q(\araddr [22] ), .QN(pc_$_SDFFE_PP0P__Q_8_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_B ) );
DFF_X1 pc_$_SDFFE_PP0P__Q_9 ( .D(_0035_ ), .CK(_1211_ ), .Q(\araddr [21] ), .QN(_1233_ ) );
DFF_X1 pc_$_SDFFE_PP1P__Q ( .D(_0036_ ), .CK(_1211_ ), .Q(\araddr [31] ), .QN(_1232_ ) );
DFF_X1 state_$_DFF_P__Q ( .D(state_$_DFF_P__Q_D ), .CK(clock ), .Q(\state [2] ), .QN(_1630_ ) );
DFF_X1 state_$_DFF_P__Q_1 ( .D(state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\state [1] ), .QN(_1631_ ) );
DFF_X1 state_$_DFF_P__Q_2 ( .D(state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\state [0] ), .QN(check_assert_$_DFFE_PP__Q_E_$_ANDNOT__Y_B_$_MUX__Y_A ) );
DFF_X1 tmp_offset_$_SDFFE_PP0P__Q ( .D(_0037_ ), .CK(_1209_ ), .Q(\tmp_offset [2] ), .QN(_1629_ ) );
DFF_X1 to_reset_$_SDFF_PP0__Q ( .D(_0039_ ), .CK(clock ), .Q(to_reset ), .QN(_1230_ ) );
DFF_X1 wen_$_SDFFE_PP0P__Q ( .D(_0038_ ), .CK(_1208_ ), .Q(\myicache.wen ), .QN(_1231_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(fanout_net_2 ), .Z(\araddr [3] ) );
BUF_X8 fanout_buf_3 ( .A(fanout_net_2 ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(fanout_net_2 ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(fanout_net_2 ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(fanout_net_6 ), .Z(\araddr [4] ) );
BUF_X8 fanout_buf_7 ( .A(fanout_net_6 ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(fanout_net_6 ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(fanout_net_6 ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(to_reset ), .Z(fanout_net_11 ) );

endmodule
