//Generate the verilog at 2025-11-14T20:46:19 by iSTA.
module ysyx_24110017 (
clock,
io_interrupt,
io_master_arready,
io_master_arvalid,
io_master_awready,
io_master_awvalid,
io_master_bready,
io_master_bvalid,
io_master_rlast,
io_master_rready,
io_master_rvalid,
io_master_wlast,
io_master_wready,
io_master_wvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_awready,
io_slave_awvalid,
io_slave_bready,
io_slave_bvalid,
io_slave_rlast,
io_slave_rready,
io_slave_rvalid,
io_slave_wlast,
io_slave_wready,
io_slave_wvalid,
reset,
io_master_araddr,
io_master_arburst,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_awaddr,
io_master_awburst,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_bid,
io_master_bresp,
io_master_rdata,
io_master_rid,
io_master_rresp,
io_master_wdata,
io_master_wstrb,
io_slave_araddr,
io_slave_arburst,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_awaddr,
io_slave_awburst,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_bid,
io_slave_bresp,
io_slave_rdata,
io_slave_rid,
io_slave_rresp,
io_slave_wdata,
io_slave_wstrb
);

input clock ;
input io_interrupt ;
input io_master_arready ;
output io_master_arvalid ;
input io_master_awready ;
output io_master_awvalid ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_rlast ;
output io_master_rready ;
input io_master_rvalid ;
output io_master_wlast ;
input io_master_wready ;
output io_master_wvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
output io_slave_awready ;
input io_slave_awvalid ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_rlast ;
input io_slave_rready ;
output io_slave_rvalid ;
input io_slave_wlast ;
output io_slave_wready ;
input io_slave_wvalid ;
input reset ;
output [31:0] io_master_araddr ;
output [1:0] io_master_arburst ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [31:0] io_master_awaddr ;
output [1:0] io_master_awburst ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
input [3:0] io_master_bid ;
input [1:0] io_master_bresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [1:0] io_master_rresp ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [31:0] io_slave_araddr ;
input [1:0] io_slave_arburst ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [31:0] io_slave_awaddr ;
input [1:0] io_slave_awburst ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
output [3:0] io_slave_bid ;
output [1:0] io_slave_bresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;
output [1:0] io_slave_rresp ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;

wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire _08922_ ;
wire _08923_ ;
wire _08924_ ;
wire _08925_ ;
wire _08926_ ;
wire _08927_ ;
wire _08928_ ;
wire _08929_ ;
wire _08930_ ;
wire _08931_ ;
wire _08932_ ;
wire _08933_ ;
wire _08934_ ;
wire _08935_ ;
wire _08936_ ;
wire _08937_ ;
wire _08938_ ;
wire _08939_ ;
wire _08940_ ;
wire _08941_ ;
wire _08942_ ;
wire _08943_ ;
wire _08944_ ;
wire _08945_ ;
wire _08946_ ;
wire _08947_ ;
wire _08948_ ;
wire _08949_ ;
wire _08950_ ;
wire _08951_ ;
wire _08952_ ;
wire _08953_ ;
wire _08954_ ;
wire _08955_ ;
wire _08956_ ;
wire _08957_ ;
wire _08958_ ;
wire _08959_ ;
wire _08960_ ;
wire _08961_ ;
wire _08962_ ;
wire _08963_ ;
wire _08964_ ;
wire _08965_ ;
wire _08966_ ;
wire _08967_ ;
wire _08968_ ;
wire _08969_ ;
wire _08970_ ;
wire _08971_ ;
wire _08972_ ;
wire _08973_ ;
wire _08974_ ;
wire _08975_ ;
wire _08976_ ;
wire _08977_ ;
wire _08978_ ;
wire _08979_ ;
wire _08980_ ;
wire _08981_ ;
wire _08982_ ;
wire _08983_ ;
wire _08984_ ;
wire _08985_ ;
wire _08986_ ;
wire _08987_ ;
wire _08988_ ;
wire _08989_ ;
wire _08990_ ;
wire _08991_ ;
wire _08992_ ;
wire _08993_ ;
wire _08994_ ;
wire _08995_ ;
wire _08996_ ;
wire _08997_ ;
wire _08998_ ;
wire _08999_ ;
wire _09000_ ;
wire _09001_ ;
wire _09002_ ;
wire _09003_ ;
wire _09004_ ;
wire _09005_ ;
wire _09006_ ;
wire _09007_ ;
wire _09008_ ;
wire _09009_ ;
wire _09010_ ;
wire _09011_ ;
wire _09012_ ;
wire _09013_ ;
wire _09014_ ;
wire _09015_ ;
wire _09016_ ;
wire _09017_ ;
wire _09018_ ;
wire _09019_ ;
wire _09020_ ;
wire _09021_ ;
wire _09022_ ;
wire _09023_ ;
wire _09024_ ;
wire _09025_ ;
wire _09026_ ;
wire _09027_ ;
wire _09028_ ;
wire _09029_ ;
wire _09030_ ;
wire _09031_ ;
wire _09032_ ;
wire _09033_ ;
wire _09034_ ;
wire _09035_ ;
wire _09036_ ;
wire _09037_ ;
wire _09038_ ;
wire _09039_ ;
wire _09040_ ;
wire _09041_ ;
wire _09042_ ;
wire _09043_ ;
wire _09044_ ;
wire _09045_ ;
wire _09046_ ;
wire _09047_ ;
wire _09048_ ;
wire _09049_ ;
wire _09050_ ;
wire _09051_ ;
wire _09052_ ;
wire _09053_ ;
wire _09054_ ;
wire _09055_ ;
wire _09056_ ;
wire _09057_ ;
wire _09058_ ;
wire _09059_ ;
wire _09060_ ;
wire _09061_ ;
wire _09062_ ;
wire _09063_ ;
wire _09064_ ;
wire _09065_ ;
wire _09066_ ;
wire _09067_ ;
wire _09068_ ;
wire _09069_ ;
wire _09070_ ;
wire _09071_ ;
wire _09072_ ;
wire _09073_ ;
wire _09074_ ;
wire _09075_ ;
wire _09076_ ;
wire _09077_ ;
wire _09078_ ;
wire _09079_ ;
wire _09080_ ;
wire _09081_ ;
wire _09082_ ;
wire _09083_ ;
wire _09084_ ;
wire _09085_ ;
wire _09086_ ;
wire _09087_ ;
wire _09088_ ;
wire _09089_ ;
wire _09090_ ;
wire _09091_ ;
wire _09092_ ;
wire _09093_ ;
wire _09094_ ;
wire _09095_ ;
wire _09096_ ;
wire _09097_ ;
wire _09098_ ;
wire _09099_ ;
wire _09100_ ;
wire _09101_ ;
wire _09102_ ;
wire _09103_ ;
wire _09104_ ;
wire _09105_ ;
wire _09106_ ;
wire _09107_ ;
wire _09108_ ;
wire _09109_ ;
wire _09110_ ;
wire _09111_ ;
wire _09112_ ;
wire _09113_ ;
wire _09114_ ;
wire _09115_ ;
wire _09116_ ;
wire _09117_ ;
wire _09118_ ;
wire _09119_ ;
wire _09120_ ;
wire _09121_ ;
wire _09122_ ;
wire _09123_ ;
wire _09124_ ;
wire _09125_ ;
wire _09126_ ;
wire _09127_ ;
wire _09128_ ;
wire _09129_ ;
wire _09130_ ;
wire _09131_ ;
wire _09132_ ;
wire _09133_ ;
wire _09134_ ;
wire _09135_ ;
wire _09136_ ;
wire _09137_ ;
wire _09138_ ;
wire _09139_ ;
wire _09140_ ;
wire _09141_ ;
wire _09142_ ;
wire _09143_ ;
wire _09144_ ;
wire _09145_ ;
wire _09146_ ;
wire _09147_ ;
wire _09148_ ;
wire _09149_ ;
wire _09150_ ;
wire _09151_ ;
wire _09152_ ;
wire _09153_ ;
wire _09154_ ;
wire _09155_ ;
wire _09156_ ;
wire _09157_ ;
wire _09158_ ;
wire _09159_ ;
wire _09160_ ;
wire _09161_ ;
wire _09162_ ;
wire _09163_ ;
wire _09164_ ;
wire _09165_ ;
wire _09166_ ;
wire _09167_ ;
wire _09168_ ;
wire _09169_ ;
wire _09170_ ;
wire _09171_ ;
wire _09172_ ;
wire _09173_ ;
wire _09174_ ;
wire _09175_ ;
wire _09176_ ;
wire _09177_ ;
wire _09178_ ;
wire _09179_ ;
wire _09180_ ;
wire _09181_ ;
wire _09182_ ;
wire _09183_ ;
wire _09184_ ;
wire _09185_ ;
wire _09186_ ;
wire _09187_ ;
wire _09188_ ;
wire _09189_ ;
wire _09190_ ;
wire _09191_ ;
wire _09192_ ;
wire _09193_ ;
wire _09194_ ;
wire _09195_ ;
wire _09196_ ;
wire _09197_ ;
wire _09198_ ;
wire _09199_ ;
wire _09200_ ;
wire _09201_ ;
wire _09202_ ;
wire _09203_ ;
wire _09204_ ;
wire _09205_ ;
wire _09206_ ;
wire _09207_ ;
wire _09208_ ;
wire _09209_ ;
wire _09210_ ;
wire _09211_ ;
wire _09212_ ;
wire _09213_ ;
wire _09214_ ;
wire _09215_ ;
wire _09216_ ;
wire _09217_ ;
wire _09218_ ;
wire _09219_ ;
wire _09220_ ;
wire _09221_ ;
wire _09222_ ;
wire _09223_ ;
wire _09224_ ;
wire _09225_ ;
wire _09226_ ;
wire _09227_ ;
wire _09228_ ;
wire _09229_ ;
wire _09230_ ;
wire _09231_ ;
wire _09232_ ;
wire _09233_ ;
wire _09234_ ;
wire _09235_ ;
wire _09236_ ;
wire _09237_ ;
wire _09238_ ;
wire _09239_ ;
wire _09240_ ;
wire _09241_ ;
wire _09242_ ;
wire _09243_ ;
wire _09244_ ;
wire _09245_ ;
wire _09246_ ;
wire _09247_ ;
wire _09248_ ;
wire _09249_ ;
wire _09250_ ;
wire _09251_ ;
wire _09252_ ;
wire _09253_ ;
wire _09254_ ;
wire _09255_ ;
wire _09256_ ;
wire _09257_ ;
wire _09258_ ;
wire _09259_ ;
wire _09260_ ;
wire _09261_ ;
wire _09262_ ;
wire _09263_ ;
wire _09264_ ;
wire _09265_ ;
wire _09266_ ;
wire _09267_ ;
wire _09268_ ;
wire _09269_ ;
wire _09270_ ;
wire _09271_ ;
wire _09272_ ;
wire _09273_ ;
wire _09274_ ;
wire _09275_ ;
wire _09276_ ;
wire _09277_ ;
wire _09278_ ;
wire _09279_ ;
wire _09280_ ;
wire _09281_ ;
wire _09282_ ;
wire _09283_ ;
wire _09284_ ;
wire _09285_ ;
wire _09286_ ;
wire _09287_ ;
wire _09288_ ;
wire _09289_ ;
wire _09290_ ;
wire _09291_ ;
wire _09292_ ;
wire _09293_ ;
wire _09294_ ;
wire _09295_ ;
wire _09296_ ;
wire _09297_ ;
wire _09298_ ;
wire _09299_ ;
wire _09300_ ;
wire _09301_ ;
wire _09302_ ;
wire _09303_ ;
wire _09304_ ;
wire _09305_ ;
wire _09306_ ;
wire _09307_ ;
wire _09308_ ;
wire _09309_ ;
wire _09310_ ;
wire _09311_ ;
wire _09312_ ;
wire _09313_ ;
wire _09314_ ;
wire _09315_ ;
wire _09316_ ;
wire _09317_ ;
wire _09318_ ;
wire _09319_ ;
wire _09320_ ;
wire _09321_ ;
wire _09322_ ;
wire _09323_ ;
wire _09324_ ;
wire _09325_ ;
wire _09326_ ;
wire _09327_ ;
wire _09328_ ;
wire _09329_ ;
wire _09330_ ;
wire _09331_ ;
wire _09332_ ;
wire _09333_ ;
wire _09334_ ;
wire _09335_ ;
wire _09336_ ;
wire _09337_ ;
wire _09338_ ;
wire _09339_ ;
wire _09340_ ;
wire _09341_ ;
wire _09342_ ;
wire _09343_ ;
wire _09344_ ;
wire _09345_ ;
wire _09346_ ;
wire _09347_ ;
wire _09348_ ;
wire _09349_ ;
wire _09350_ ;
wire _09351_ ;
wire _09352_ ;
wire _09353_ ;
wire _09354_ ;
wire _09355_ ;
wire _09356_ ;
wire _09357_ ;
wire _09358_ ;
wire _09359_ ;
wire _09360_ ;
wire _09361_ ;
wire _09362_ ;
wire _09363_ ;
wire _09364_ ;
wire _09365_ ;
wire _09366_ ;
wire _09367_ ;
wire _09368_ ;
wire _09369_ ;
wire _09370_ ;
wire _09371_ ;
wire _09372_ ;
wire _09373_ ;
wire _09374_ ;
wire _09375_ ;
wire _09376_ ;
wire _09377_ ;
wire _09378_ ;
wire _09379_ ;
wire _09380_ ;
wire _09381_ ;
wire _09382_ ;
wire _09383_ ;
wire _09384_ ;
wire _09385_ ;
wire _09386_ ;
wire _09387_ ;
wire _09388_ ;
wire _09389_ ;
wire _09390_ ;
wire _09391_ ;
wire _09392_ ;
wire _09393_ ;
wire _09394_ ;
wire _09395_ ;
wire _09396_ ;
wire _09397_ ;
wire _09398_ ;
wire _09399_ ;
wire _09400_ ;
wire _09401_ ;
wire _09402_ ;
wire _09403_ ;
wire _09404_ ;
wire _09405_ ;
wire _09406_ ;
wire _09407_ ;
wire _09408_ ;
wire _09409_ ;
wire _09410_ ;
wire _09411_ ;
wire _09412_ ;
wire _09413_ ;
wire _09414_ ;
wire _09415_ ;
wire _09416_ ;
wire _09417_ ;
wire _09418_ ;
wire _09419_ ;
wire _09420_ ;
wire _09421_ ;
wire _09422_ ;
wire _09423_ ;
wire _09424_ ;
wire _09425_ ;
wire _09426_ ;
wire _09427_ ;
wire _09428_ ;
wire _09429_ ;
wire _09430_ ;
wire _09431_ ;
wire _09432_ ;
wire _09433_ ;
wire _09434_ ;
wire _09435_ ;
wire _09436_ ;
wire _09437_ ;
wire _09438_ ;
wire _09439_ ;
wire _09440_ ;
wire _09441_ ;
wire _09442_ ;
wire _09443_ ;
wire _09444_ ;
wire _09445_ ;
wire _09446_ ;
wire _09447_ ;
wire _09448_ ;
wire _09449_ ;
wire _09450_ ;
wire _09451_ ;
wire _09452_ ;
wire _09453_ ;
wire _09454_ ;
wire _09455_ ;
wire _09456_ ;
wire _09457_ ;
wire _09458_ ;
wire _09459_ ;
wire _09460_ ;
wire _09461_ ;
wire _09462_ ;
wire _09463_ ;
wire _09464_ ;
wire _09465_ ;
wire _09466_ ;
wire _09467_ ;
wire _09468_ ;
wire _09469_ ;
wire _09470_ ;
wire _09471_ ;
wire _09472_ ;
wire _09473_ ;
wire _09474_ ;
wire _09475_ ;
wire _09476_ ;
wire _09477_ ;
wire _09478_ ;
wire _09479_ ;
wire _09480_ ;
wire _09481_ ;
wire _09482_ ;
wire _09483_ ;
wire _09484_ ;
wire _09485_ ;
wire _09486_ ;
wire _09487_ ;
wire _09488_ ;
wire _09489_ ;
wire _09490_ ;
wire _09491_ ;
wire _09492_ ;
wire _09493_ ;
wire _09494_ ;
wire _09495_ ;
wire _09496_ ;
wire _09497_ ;
wire _09498_ ;
wire _09499_ ;
wire _09500_ ;
wire _09501_ ;
wire _09502_ ;
wire _09503_ ;
wire _09504_ ;
wire _09505_ ;
wire _09506_ ;
wire _09507_ ;
wire _09508_ ;
wire _09509_ ;
wire _09510_ ;
wire _09511_ ;
wire _09512_ ;
wire _09513_ ;
wire _09514_ ;
wire _09515_ ;
wire _09516_ ;
wire _09517_ ;
wire _09518_ ;
wire _09519_ ;
wire _09520_ ;
wire _09521_ ;
wire _09522_ ;
wire _09523_ ;
wire _09524_ ;
wire _09525_ ;
wire _09526_ ;
wire _09527_ ;
wire _09528_ ;
wire _09529_ ;
wire _09530_ ;
wire _09531_ ;
wire _09532_ ;
wire _09533_ ;
wire _09534_ ;
wire _09535_ ;
wire _09536_ ;
wire _09537_ ;
wire _09538_ ;
wire _09539_ ;
wire _09540_ ;
wire _09541_ ;
wire _09542_ ;
wire _09543_ ;
wire _09544_ ;
wire _09545_ ;
wire _09546_ ;
wire _09547_ ;
wire _09548_ ;
wire _09549_ ;
wire _09550_ ;
wire _09551_ ;
wire _09552_ ;
wire _09553_ ;
wire _09554_ ;
wire _09555_ ;
wire _09556_ ;
wire _09557_ ;
wire _09558_ ;
wire _09559_ ;
wire _09560_ ;
wire _09561_ ;
wire _09562_ ;
wire _09563_ ;
wire _09564_ ;
wire _09565_ ;
wire _09566_ ;
wire _09567_ ;
wire _09568_ ;
wire _09569_ ;
wire _09570_ ;
wire _09571_ ;
wire _09572_ ;
wire _09573_ ;
wire _09574_ ;
wire _09575_ ;
wire _09576_ ;
wire _09577_ ;
wire _09578_ ;
wire _09579_ ;
wire _09580_ ;
wire _09581_ ;
wire _09582_ ;
wire _09583_ ;
wire _09584_ ;
wire _09585_ ;
wire _09586_ ;
wire _09587_ ;
wire _09588_ ;
wire _09589_ ;
wire _09590_ ;
wire _09591_ ;
wire _09592_ ;
wire _09593_ ;
wire _09594_ ;
wire _09595_ ;
wire _09596_ ;
wire _09597_ ;
wire _09598_ ;
wire _09599_ ;
wire _09600_ ;
wire _09601_ ;
wire _09602_ ;
wire _09603_ ;
wire _09604_ ;
wire _09605_ ;
wire _09606_ ;
wire _09607_ ;
wire _09608_ ;
wire _09609_ ;
wire _09610_ ;
wire _09611_ ;
wire _09612_ ;
wire _09613_ ;
wire _09614_ ;
wire _09615_ ;
wire _09616_ ;
wire _09617_ ;
wire _09618_ ;
wire _09619_ ;
wire _09620_ ;
wire _09621_ ;
wire _09622_ ;
wire _09623_ ;
wire _09624_ ;
wire _09625_ ;
wire _09626_ ;
wire _09627_ ;
wire _09628_ ;
wire _09629_ ;
wire _09630_ ;
wire _09631_ ;
wire _09632_ ;
wire _09633_ ;
wire _09634_ ;
wire _09635_ ;
wire _09636_ ;
wire _09637_ ;
wire _09638_ ;
wire _09639_ ;
wire _09640_ ;
wire _09641_ ;
wire _09642_ ;
wire _09643_ ;
wire _09644_ ;
wire _09645_ ;
wire _09646_ ;
wire _09647_ ;
wire _09648_ ;
wire _09649_ ;
wire _09650_ ;
wire _09651_ ;
wire _09652_ ;
wire _09653_ ;
wire _09654_ ;
wire _09655_ ;
wire _09656_ ;
wire _09657_ ;
wire _09658_ ;
wire _09659_ ;
wire _09660_ ;
wire _09661_ ;
wire _09662_ ;
wire _09663_ ;
wire _09664_ ;
wire _09665_ ;
wire _09666_ ;
wire _09667_ ;
wire _09668_ ;
wire _09669_ ;
wire _09670_ ;
wire _09671_ ;
wire _09672_ ;
wire _09673_ ;
wire _09674_ ;
wire _09675_ ;
wire _09676_ ;
wire _09677_ ;
wire _09678_ ;
wire _09679_ ;
wire _09680_ ;
wire _09681_ ;
wire _09682_ ;
wire _09683_ ;
wire _09684_ ;
wire _09685_ ;
wire _09686_ ;
wire _09687_ ;
wire _09688_ ;
wire _09689_ ;
wire _09690_ ;
wire _09691_ ;
wire _09692_ ;
wire _09693_ ;
wire _09694_ ;
wire _09695_ ;
wire _09696_ ;
wire _09697_ ;
wire _09698_ ;
wire _09699_ ;
wire _09700_ ;
wire _09701_ ;
wire _09702_ ;
wire _09703_ ;
wire _09704_ ;
wire _09705_ ;
wire _09706_ ;
wire _09707_ ;
wire _09708_ ;
wire _09709_ ;
wire _09710_ ;
wire _09711_ ;
wire _09712_ ;
wire _09713_ ;
wire _09714_ ;
wire _09715_ ;
wire _09716_ ;
wire _09717_ ;
wire _09718_ ;
wire _09719_ ;
wire _09720_ ;
wire _09721_ ;
wire _09722_ ;
wire _09723_ ;
wire _09724_ ;
wire _09725_ ;
wire _09726_ ;
wire _09727_ ;
wire _09728_ ;
wire _09729_ ;
wire _09730_ ;
wire _09731_ ;
wire _09732_ ;
wire _09733_ ;
wire _09734_ ;
wire _09735_ ;
wire _09736_ ;
wire _09737_ ;
wire _09738_ ;
wire _09739_ ;
wire _09740_ ;
wire _09741_ ;
wire _09742_ ;
wire _09743_ ;
wire _09744_ ;
wire _09745_ ;
wire _09746_ ;
wire _09747_ ;
wire _09748_ ;
wire _09749_ ;
wire _09750_ ;
wire _09751_ ;
wire _09752_ ;
wire _09753_ ;
wire _09754_ ;
wire _09755_ ;
wire _09756_ ;
wire _09757_ ;
wire _09758_ ;
wire _09759_ ;
wire _09760_ ;
wire _09761_ ;
wire _09762_ ;
wire _09763_ ;
wire _09764_ ;
wire _09765_ ;
wire _09766_ ;
wire _09767_ ;
wire _09768_ ;
wire _09769_ ;
wire _09770_ ;
wire _09771_ ;
wire _09772_ ;
wire _09773_ ;
wire _09774_ ;
wire _09775_ ;
wire _09776_ ;
wire _09777_ ;
wire _09778_ ;
wire _09779_ ;
wire _09780_ ;
wire _09781_ ;
wire _09782_ ;
wire _09783_ ;
wire _09784_ ;
wire _09785_ ;
wire _09786_ ;
wire _09787_ ;
wire _09788_ ;
wire _09789_ ;
wire _09790_ ;
wire _09791_ ;
wire _09792_ ;
wire _09793_ ;
wire _09794_ ;
wire _09795_ ;
wire _09796_ ;
wire _09797_ ;
wire _09798_ ;
wire _09799_ ;
wire _09800_ ;
wire _09801_ ;
wire _09802_ ;
wire _09803_ ;
wire _09804_ ;
wire _09805_ ;
wire _09806_ ;
wire _09807_ ;
wire _09808_ ;
wire _09809_ ;
wire _09810_ ;
wire _09811_ ;
wire _09812_ ;
wire _09813_ ;
wire _09814_ ;
wire _09815_ ;
wire _09816_ ;
wire _09817_ ;
wire _09818_ ;
wire _09819_ ;
wire _09820_ ;
wire _09821_ ;
wire _09822_ ;
wire _09823_ ;
wire _09824_ ;
wire _09825_ ;
wire _09826_ ;
wire _09827_ ;
wire _09828_ ;
wire _09829_ ;
wire _09830_ ;
wire _09831_ ;
wire _09832_ ;
wire _09833_ ;
wire _09834_ ;
wire _09835_ ;
wire _09836_ ;
wire _09837_ ;
wire _09838_ ;
wire _09839_ ;
wire _09840_ ;
wire _09841_ ;
wire _09842_ ;
wire _09843_ ;
wire _09844_ ;
wire _09845_ ;
wire _09846_ ;
wire _09847_ ;
wire _09848_ ;
wire _09849_ ;
wire _09850_ ;
wire _09851_ ;
wire _09852_ ;
wire _09853_ ;
wire _09854_ ;
wire _09855_ ;
wire _09856_ ;
wire _09857_ ;
wire _09858_ ;
wire _09859_ ;
wire _09860_ ;
wire _09861_ ;
wire _09862_ ;
wire _09863_ ;
wire _09864_ ;
wire _09865_ ;
wire _09866_ ;
wire _09867_ ;
wire _09868_ ;
wire _09869_ ;
wire _09870_ ;
wire _09871_ ;
wire _09872_ ;
wire _09873_ ;
wire _09874_ ;
wire _09875_ ;
wire _09876_ ;
wire _09877_ ;
wire _09878_ ;
wire _09879_ ;
wire _09880_ ;
wire _09881_ ;
wire _09882_ ;
wire _09883_ ;
wire _09884_ ;
wire _09885_ ;
wire _09886_ ;
wire _09887_ ;
wire _09888_ ;
wire _09889_ ;
wire _09890_ ;
wire _09891_ ;
wire _09892_ ;
wire _09893_ ;
wire _09894_ ;
wire _09895_ ;
wire _09896_ ;
wire _09897_ ;
wire _09898_ ;
wire _09899_ ;
wire _09900_ ;
wire _09901_ ;
wire _09902_ ;
wire _09903_ ;
wire _09904_ ;
wire _09905_ ;
wire _09906_ ;
wire _09907_ ;
wire _09908_ ;
wire _09909_ ;
wire _09910_ ;
wire _09911_ ;
wire _09912_ ;
wire _09913_ ;
wire _09914_ ;
wire _09915_ ;
wire _09916_ ;
wire _09917_ ;
wire _09918_ ;
wire _09919_ ;
wire _09920_ ;
wire _09921_ ;
wire _09922_ ;
wire _09923_ ;
wire _09924_ ;
wire _09925_ ;
wire _09926_ ;
wire _09927_ ;
wire _09928_ ;
wire _09929_ ;
wire _09930_ ;
wire _09931_ ;
wire _09932_ ;
wire _09933_ ;
wire _09934_ ;
wire _09935_ ;
wire _09936_ ;
wire _09937_ ;
wire _09938_ ;
wire _09939_ ;
wire _09940_ ;
wire _09941_ ;
wire _09942_ ;
wire _09943_ ;
wire _09944_ ;
wire _09945_ ;
wire _09946_ ;
wire _09947_ ;
wire _09948_ ;
wire _09949_ ;
wire _09950_ ;
wire _09951_ ;
wire _09952_ ;
wire _09953_ ;
wire _09954_ ;
wire _09955_ ;
wire _09956_ ;
wire _09957_ ;
wire _09958_ ;
wire _09959_ ;
wire _09960_ ;
wire _09961_ ;
wire _09962_ ;
wire _09963_ ;
wire _09964_ ;
wire _09965_ ;
wire _09966_ ;
wire _09967_ ;
wire _09968_ ;
wire _09969_ ;
wire _09970_ ;
wire _09971_ ;
wire _09972_ ;
wire _09973_ ;
wire _09974_ ;
wire _09975_ ;
wire _09976_ ;
wire _09977_ ;
wire _09978_ ;
wire _09979_ ;
wire _09980_ ;
wire _09981_ ;
wire _09982_ ;
wire _09983_ ;
wire _09984_ ;
wire _09985_ ;
wire _09986_ ;
wire _09987_ ;
wire _09988_ ;
wire _09989_ ;
wire _09990_ ;
wire _09991_ ;
wire _09992_ ;
wire _09993_ ;
wire _09994_ ;
wire _09995_ ;
wire _09996_ ;
wire _09997_ ;
wire _09998_ ;
wire _09999_ ;
wire _10000_ ;
wire _10001_ ;
wire _10002_ ;
wire _10003_ ;
wire _10004_ ;
wire _10005_ ;
wire _10006_ ;
wire _10007_ ;
wire _10008_ ;
wire _10009_ ;
wire _10010_ ;
wire _10011_ ;
wire _10012_ ;
wire _10013_ ;
wire _10014_ ;
wire _10015_ ;
wire _10016_ ;
wire _10017_ ;
wire _10018_ ;
wire _10019_ ;
wire _10020_ ;
wire _10021_ ;
wire _10022_ ;
wire _10023_ ;
wire _10024_ ;
wire _10025_ ;
wire _10026_ ;
wire _10027_ ;
wire _10028_ ;
wire _10029_ ;
wire _10030_ ;
wire _10031_ ;
wire _10032_ ;
wire _10033_ ;
wire _10034_ ;
wire _10035_ ;
wire _10036_ ;
wire _10037_ ;
wire _10038_ ;
wire _10039_ ;
wire _10040_ ;
wire _10041_ ;
wire _10042_ ;
wire _10043_ ;
wire _10044_ ;
wire _10045_ ;
wire _10046_ ;
wire _10047_ ;
wire _10048_ ;
wire _10049_ ;
wire _10050_ ;
wire _10051_ ;
wire _10052_ ;
wire _10053_ ;
wire _10054_ ;
wire _10055_ ;
wire _10056_ ;
wire _10057_ ;
wire _10058_ ;
wire _10059_ ;
wire _10060_ ;
wire _10061_ ;
wire _10062_ ;
wire _10063_ ;
wire _10064_ ;
wire _10065_ ;
wire _10066_ ;
wire _10067_ ;
wire _10068_ ;
wire _10069_ ;
wire _10070_ ;
wire _10071_ ;
wire _10072_ ;
wire _10073_ ;
wire _10074_ ;
wire _10075_ ;
wire _10076_ ;
wire _10077_ ;
wire _10078_ ;
wire _10079_ ;
wire _10080_ ;
wire _10081_ ;
wire _10082_ ;
wire _10083_ ;
wire _10084_ ;
wire _10085_ ;
wire _10086_ ;
wire _10087_ ;
wire _10088_ ;
wire _10089_ ;
wire _10090_ ;
wire _10091_ ;
wire _10092_ ;
wire _10093_ ;
wire _10094_ ;
wire _10095_ ;
wire _10096_ ;
wire _10097_ ;
wire _10098_ ;
wire _10099_ ;
wire _10100_ ;
wire _10101_ ;
wire _10102_ ;
wire _10103_ ;
wire _10104_ ;
wire _10105_ ;
wire _10106_ ;
wire _10107_ ;
wire _10108_ ;
wire _10109_ ;
wire _10110_ ;
wire _10111_ ;
wire _10112_ ;
wire _10113_ ;
wire _10114_ ;
wire _10115_ ;
wire _10116_ ;
wire _10117_ ;
wire _10118_ ;
wire _10119_ ;
wire _10120_ ;
wire _10121_ ;
wire _10122_ ;
wire _10123_ ;
wire _10124_ ;
wire _10125_ ;
wire _10126_ ;
wire _10127_ ;
wire _10128_ ;
wire _10129_ ;
wire _10130_ ;
wire _10131_ ;
wire _10132_ ;
wire _10133_ ;
wire _10134_ ;
wire _10135_ ;
wire _10136_ ;
wire _10137_ ;
wire _10138_ ;
wire _10139_ ;
wire _10140_ ;
wire _10141_ ;
wire _10142_ ;
wire _10143_ ;
wire _10144_ ;
wire _10145_ ;
wire _10146_ ;
wire _10147_ ;
wire _10148_ ;
wire _10149_ ;
wire _10150_ ;
wire _10151_ ;
wire _10152_ ;
wire _10153_ ;
wire _10154_ ;
wire _10155_ ;
wire _10156_ ;
wire _10157_ ;
wire _10158_ ;
wire _10159_ ;
wire _10160_ ;
wire _10161_ ;
wire _10162_ ;
wire _10163_ ;
wire _10164_ ;
wire _10165_ ;
wire _10166_ ;
wire _10167_ ;
wire _10168_ ;
wire _10169_ ;
wire _10170_ ;
wire _10171_ ;
wire _10172_ ;
wire _10173_ ;
wire _10174_ ;
wire _10175_ ;
wire _10176_ ;
wire _10177_ ;
wire _10178_ ;
wire _10179_ ;
wire _10180_ ;
wire _10181_ ;
wire _10182_ ;
wire _10183_ ;
wire _10184_ ;
wire _10185_ ;
wire _10186_ ;
wire _10187_ ;
wire _10188_ ;
wire _10189_ ;
wire _10190_ ;
wire _10191_ ;
wire _10192_ ;
wire _10193_ ;
wire _10194_ ;
wire _10195_ ;
wire _10196_ ;
wire _10197_ ;
wire _10198_ ;
wire _10199_ ;
wire _10200_ ;
wire _10201_ ;
wire _10202_ ;
wire _10203_ ;
wire _10204_ ;
wire _10205_ ;
wire _10206_ ;
wire _10207_ ;
wire _10208_ ;
wire _10209_ ;
wire _10210_ ;
wire _10211_ ;
wire _10212_ ;
wire _10213_ ;
wire _10214_ ;
wire _10215_ ;
wire _10216_ ;
wire _10217_ ;
wire _10218_ ;
wire _10219_ ;
wire _10220_ ;
wire _10221_ ;
wire _10222_ ;
wire _10223_ ;
wire _10224_ ;
wire _10225_ ;
wire _10226_ ;
wire _10227_ ;
wire _10228_ ;
wire _10229_ ;
wire _10230_ ;
wire _10231_ ;
wire _10232_ ;
wire _10233_ ;
wire _10234_ ;
wire _10235_ ;
wire _10236_ ;
wire _10237_ ;
wire _10238_ ;
wire _10239_ ;
wire _10240_ ;
wire _10241_ ;
wire _10242_ ;
wire _10243_ ;
wire _10244_ ;
wire _10245_ ;
wire _10246_ ;
wire _10247_ ;
wire _10248_ ;
wire _10249_ ;
wire _10250_ ;
wire _10251_ ;
wire _10252_ ;
wire _10253_ ;
wire _10254_ ;
wire _10255_ ;
wire _10256_ ;
wire _10257_ ;
wire _10258_ ;
wire _10259_ ;
wire _10260_ ;
wire _10261_ ;
wire _10262_ ;
wire _10263_ ;
wire _10264_ ;
wire _10265_ ;
wire _10266_ ;
wire _10267_ ;
wire _10268_ ;
wire _10269_ ;
wire _10270_ ;
wire _10271_ ;
wire _10272_ ;
wire _10273_ ;
wire _10274_ ;
wire _10275_ ;
wire _10276_ ;
wire _10277_ ;
wire _10278_ ;
wire _10279_ ;
wire _10280_ ;
wire _10281_ ;
wire _10282_ ;
wire _10283_ ;
wire _10284_ ;
wire _10285_ ;
wire _10286_ ;
wire _10287_ ;
wire _10288_ ;
wire _10289_ ;
wire _10290_ ;
wire _10291_ ;
wire _10292_ ;
wire _10293_ ;
wire _10294_ ;
wire _10295_ ;
wire _10296_ ;
wire _10297_ ;
wire _10298_ ;
wire _10299_ ;
wire _10300_ ;
wire _10301_ ;
wire _10302_ ;
wire _10303_ ;
wire _10304_ ;
wire _10305_ ;
wire _10306_ ;
wire _10307_ ;
wire _10308_ ;
wire _10309_ ;
wire _10310_ ;
wire _10311_ ;
wire _10312_ ;
wire _10313_ ;
wire _10314_ ;
wire _10315_ ;
wire _10316_ ;
wire _10317_ ;
wire _10318_ ;
wire _10319_ ;
wire _10320_ ;
wire _10321_ ;
wire _10322_ ;
wire _10323_ ;
wire _10324_ ;
wire _10325_ ;
wire _10326_ ;
wire _10327_ ;
wire _10328_ ;
wire _10329_ ;
wire _10330_ ;
wire _10331_ ;
wire _10332_ ;
wire _10333_ ;
wire _10334_ ;
wire _10335_ ;
wire _10336_ ;
wire _10337_ ;
wire _10338_ ;
wire _10339_ ;
wire _10340_ ;
wire _10341_ ;
wire _10342_ ;
wire _10343_ ;
wire _10344_ ;
wire _10345_ ;
wire _10346_ ;
wire _10347_ ;
wire _10348_ ;
wire _10349_ ;
wire _10350_ ;
wire _10351_ ;
wire _10352_ ;
wire _10353_ ;
wire _10354_ ;
wire _10355_ ;
wire _10356_ ;
wire _10357_ ;
wire _10358_ ;
wire _10359_ ;
wire _10360_ ;
wire _10361_ ;
wire _10362_ ;
wire _10363_ ;
wire _10364_ ;
wire _10365_ ;
wire _10366_ ;
wire _10367_ ;
wire _10368_ ;
wire _10369_ ;
wire _10370_ ;
wire _10371_ ;
wire _10372_ ;
wire _10373_ ;
wire _10374_ ;
wire _10375_ ;
wire _10376_ ;
wire _10377_ ;
wire _10378_ ;
wire _10379_ ;
wire _10380_ ;
wire _10381_ ;
wire _10382_ ;
wire _10383_ ;
wire _10384_ ;
wire _10385_ ;
wire _10386_ ;
wire _10387_ ;
wire _10388_ ;
wire _10389_ ;
wire _10390_ ;
wire _10391_ ;
wire _10392_ ;
wire _10393_ ;
wire _10394_ ;
wire _10395_ ;
wire _10396_ ;
wire _10397_ ;
wire _10398_ ;
wire _10399_ ;
wire _10400_ ;
wire _10401_ ;
wire _10402_ ;
wire _10403_ ;
wire _10404_ ;
wire _10405_ ;
wire _10406_ ;
wire _10407_ ;
wire _10408_ ;
wire _10409_ ;
wire _10410_ ;
wire _10411_ ;
wire _10412_ ;
wire _10413_ ;
wire _10414_ ;
wire _10415_ ;
wire _10416_ ;
wire _10417_ ;
wire _10418_ ;
wire _10419_ ;
wire _10420_ ;
wire _10421_ ;
wire _10422_ ;
wire _10423_ ;
wire _10424_ ;
wire _10425_ ;
wire _10426_ ;
wire _10427_ ;
wire _10428_ ;
wire _10429_ ;
wire _10430_ ;
wire _10431_ ;
wire _10432_ ;
wire _10433_ ;
wire _10434_ ;
wire _10435_ ;
wire _10436_ ;
wire _10437_ ;
wire _10438_ ;
wire _10439_ ;
wire _10440_ ;
wire _10441_ ;
wire _10442_ ;
wire _10443_ ;
wire _10444_ ;
wire _10445_ ;
wire _10446_ ;
wire _10447_ ;
wire _10448_ ;
wire _10449_ ;
wire _10450_ ;
wire _10451_ ;
wire _10452_ ;
wire _10453_ ;
wire _10454_ ;
wire _10455_ ;
wire _10456_ ;
wire _10457_ ;
wire _10458_ ;
wire _10459_ ;
wire _10460_ ;
wire _10461_ ;
wire _10462_ ;
wire _10463_ ;
wire _10464_ ;
wire _10465_ ;
wire _10466_ ;
wire _10467_ ;
wire _10468_ ;
wire _10469_ ;
wire _10470_ ;
wire _10471_ ;
wire _10472_ ;
wire _10473_ ;
wire _10474_ ;
wire _10475_ ;
wire _10476_ ;
wire _10477_ ;
wire _10478_ ;
wire _10479_ ;
wire _10480_ ;
wire _10481_ ;
wire _10482_ ;
wire _10483_ ;
wire _10484_ ;
wire _10485_ ;
wire _10486_ ;
wire _10487_ ;
wire _10488_ ;
wire _10489_ ;
wire _10490_ ;
wire _10491_ ;
wire _10492_ ;
wire _10493_ ;
wire _10494_ ;
wire _10495_ ;
wire _10496_ ;
wire _10497_ ;
wire _10498_ ;
wire _10499_ ;
wire _10500_ ;
wire _10501_ ;
wire _10502_ ;
wire _10503_ ;
wire _10504_ ;
wire _10505_ ;
wire _10506_ ;
wire _10507_ ;
wire _10508_ ;
wire _10509_ ;
wire _10510_ ;
wire _10511_ ;
wire _10512_ ;
wire _10513_ ;
wire _10514_ ;
wire _10515_ ;
wire _10516_ ;
wire _10517_ ;
wire _10518_ ;
wire _10519_ ;
wire _10520_ ;
wire _10521_ ;
wire _10522_ ;
wire _10523_ ;
wire _10524_ ;
wire _10525_ ;
wire _10526_ ;
wire _10527_ ;
wire _10528_ ;
wire _10529_ ;
wire _10530_ ;
wire _10531_ ;
wire _10532_ ;
wire _10533_ ;
wire _10534_ ;
wire _10535_ ;
wire _10536_ ;
wire _10537_ ;
wire _10538_ ;
wire _10539_ ;
wire _10540_ ;
wire _10541_ ;
wire _10542_ ;
wire _10543_ ;
wire _10544_ ;
wire _10545_ ;
wire _10546_ ;
wire _10547_ ;
wire _10548_ ;
wire _10549_ ;
wire _10550_ ;
wire _10551_ ;
wire _10552_ ;
wire _10553_ ;
wire _10554_ ;
wire _10555_ ;
wire _10556_ ;
wire _10557_ ;
wire _10558_ ;
wire _10559_ ;
wire _10560_ ;
wire _10561_ ;
wire _10562_ ;
wire _10563_ ;
wire _10564_ ;
wire _10565_ ;
wire _10566_ ;
wire _10567_ ;
wire _10568_ ;
wire _10569_ ;
wire _10570_ ;
wire _10571_ ;
wire _10572_ ;
wire _10573_ ;
wire _10574_ ;
wire _10575_ ;
wire _10576_ ;
wire _10577_ ;
wire _10578_ ;
wire _10579_ ;
wire _10580_ ;
wire _10581_ ;
wire _10582_ ;
wire _10583_ ;
wire _10584_ ;
wire _10585_ ;
wire _10586_ ;
wire _10587_ ;
wire _10588_ ;
wire _10589_ ;
wire _10590_ ;
wire _10591_ ;
wire _10592_ ;
wire _10593_ ;
wire _10594_ ;
wire _10595_ ;
wire _10596_ ;
wire _10597_ ;
wire _10598_ ;
wire _10599_ ;
wire _10600_ ;
wire _10601_ ;
wire _10602_ ;
wire _10603_ ;
wire _10604_ ;
wire _10605_ ;
wire _10606_ ;
wire _10607_ ;
wire _10608_ ;
wire _10609_ ;
wire _10610_ ;
wire _10611_ ;
wire _10612_ ;
wire _10613_ ;
wire _10614_ ;
wire _10615_ ;
wire _10616_ ;
wire _10617_ ;
wire _10618_ ;
wire _10619_ ;
wire _10620_ ;
wire _10621_ ;
wire _10622_ ;
wire _10623_ ;
wire _10624_ ;
wire _10625_ ;
wire _10626_ ;
wire _10627_ ;
wire _10628_ ;
wire _10629_ ;
wire _10630_ ;
wire _10631_ ;
wire _10632_ ;
wire _10633_ ;
wire _10634_ ;
wire _10635_ ;
wire _10636_ ;
wire _10637_ ;
wire _10638_ ;
wire _10639_ ;
wire _10640_ ;
wire _10641_ ;
wire _10642_ ;
wire _10643_ ;
wire _10644_ ;
wire _10645_ ;
wire _10646_ ;
wire _10647_ ;
wire _10648_ ;
wire _10649_ ;
wire _10650_ ;
wire _10651_ ;
wire _10652_ ;
wire _10653_ ;
wire _10654_ ;
wire _10655_ ;
wire _10656_ ;
wire _10657_ ;
wire _10658_ ;
wire _10659_ ;
wire _10660_ ;
wire _10661_ ;
wire _10662_ ;
wire _10663_ ;
wire _10664_ ;
wire _10665_ ;
wire _10666_ ;
wire _10667_ ;
wire _10668_ ;
wire _10669_ ;
wire _10670_ ;
wire _10671_ ;
wire _10672_ ;
wire _10673_ ;
wire _10674_ ;
wire _10675_ ;
wire _10676_ ;
wire _10677_ ;
wire _10678_ ;
wire _10679_ ;
wire _10680_ ;
wire _10681_ ;
wire _10682_ ;
wire _10683_ ;
wire _10684_ ;
wire _10685_ ;
wire _10686_ ;
wire _10687_ ;
wire _10688_ ;
wire _10689_ ;
wire _10690_ ;
wire _10691_ ;
wire _10692_ ;
wire _10693_ ;
wire _10694_ ;
wire _10695_ ;
wire _10696_ ;
wire _10697_ ;
wire _10698_ ;
wire _10699_ ;
wire _10700_ ;
wire _10701_ ;
wire _10702_ ;
wire _10703_ ;
wire _10704_ ;
wire _10705_ ;
wire _10706_ ;
wire _10707_ ;
wire _10708_ ;
wire _10709_ ;
wire _10710_ ;
wire _10711_ ;
wire _10712_ ;
wire _10713_ ;
wire _10714_ ;
wire _10715_ ;
wire _10716_ ;
wire _10717_ ;
wire _10718_ ;
wire _10719_ ;
wire _10720_ ;
wire _10721_ ;
wire _10722_ ;
wire _10723_ ;
wire _10724_ ;
wire _10725_ ;
wire _10726_ ;
wire _10727_ ;
wire _10728_ ;
wire _10729_ ;
wire _10730_ ;
wire _10731_ ;
wire _10732_ ;
wire _10733_ ;
wire _10734_ ;
wire _10735_ ;
wire _10736_ ;
wire _10737_ ;
wire _10738_ ;
wire _10739_ ;
wire _10740_ ;
wire _10741_ ;
wire _10742_ ;
wire _10743_ ;
wire _10744_ ;
wire _10745_ ;
wire _10746_ ;
wire _10747_ ;
wire _10748_ ;
wire _10749_ ;
wire _10750_ ;
wire _10751_ ;
wire _10752_ ;
wire _10753_ ;
wire _10754_ ;
wire _10755_ ;
wire _10756_ ;
wire _10757_ ;
wire _10758_ ;
wire _10759_ ;
wire _10760_ ;
wire _10761_ ;
wire _10762_ ;
wire _10763_ ;
wire _10764_ ;
wire _10765_ ;
wire _10766_ ;
wire _10767_ ;
wire _10768_ ;
wire _10769_ ;
wire _10770_ ;
wire _10771_ ;
wire _10772_ ;
wire _10773_ ;
wire _10774_ ;
wire _10775_ ;
wire _10776_ ;
wire _10777_ ;
wire _10778_ ;
wire _10779_ ;
wire _10780_ ;
wire _10781_ ;
wire _10782_ ;
wire _10783_ ;
wire _10784_ ;
wire _10785_ ;
wire _10786_ ;
wire _10787_ ;
wire _10788_ ;
wire _10789_ ;
wire _10790_ ;
wire _10791_ ;
wire _10792_ ;
wire _10793_ ;
wire _10794_ ;
wire _10795_ ;
wire _10796_ ;
wire _10797_ ;
wire _10798_ ;
wire _10799_ ;
wire \BTB.bindex ;
wire \BTB.bindex_pre ;
wire \BTB.bsnpc_reg[0][0] ;
wire \BTB.bsnpc_reg[0][1] ;
wire \BTB.bsnpc_reg[0][2] ;
wire \BTB.bsnpc_reg[0][3] ;
wire \BTB.bsnpc_reg[0][4] ;
wire \BTB.bsnpc_reg[0][5] ;
wire \BTB.bsnpc_reg[0][6] ;
wire \BTB.bsnpc_reg[0][7] ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_1_Y ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_1_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_1_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_2_Y ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_2_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_2_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_3_Y ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_3_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_3_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_4_Y ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_4_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_4_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_5_Y ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_5_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_5_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_Y ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ;
wire \BTB.bsnpc_reg[0]_$_NOT__A_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ;
wire \BTB.bsnpc_reg[1][0] ;
wire \BTB.bsnpc_reg[1][1] ;
wire \BTB.bsnpc_reg[1][2] ;
wire \BTB.bsnpc_reg[1][3] ;
wire \BTB.bsnpc_reg[1][4] ;
wire \BTB.bsnpc_reg[1][5] ;
wire \BTB.bsnpc_reg[1][6] ;
wire \BTB.bsnpc_reg[1][7] ;
wire \BTB.bsnpc_reg[1]_$_NOT__A_1_Y ;
wire \BTB.bsnpc_reg[1]_$_NOT__A_2_Y ;
wire \BTB.bsnpc_reg[1]_$_NOT__A_3_Y ;
wire \BTB.bsnpc_reg[1]_$_NOT__A_4_Y ;
wire \BTB.bsnpc_reg[1]_$_NOT__A_5_Y ;
wire \BTB.bsnpc_reg[1]_$_NOT__A_Y ;
wire \BTB.btag_reg[0][0] ;
wire \BTB.btag_reg[0][10] ;
wire \BTB.btag_reg[0][11] ;
wire \BTB.btag_reg[0][12] ;
wire \BTB.btag_reg[0][1] ;
wire \BTB.btag_reg[0][2] ;
wire \BTB.btag_reg[0][3] ;
wire \BTB.btag_reg[0][4] ;
wire \BTB.btag_reg[0][5] ;
wire \BTB.btag_reg[0][6] ;
wire \BTB.btag_reg[0][7] ;
wire \BTB.btag_reg[0][8] ;
wire \BTB.btag_reg[0][9] ;
wire \BTB.btag_reg[1][0] ;
wire \BTB.btag_reg[1][10] ;
wire \BTB.btag_reg[1][11] ;
wire \BTB.btag_reg[1][12] ;
wire \BTB.btag_reg[1][1] ;
wire \BTB.btag_reg[1][2] ;
wire \BTB.btag_reg[1][3] ;
wire \BTB.btag_reg[1][4] ;
wire \BTB.btag_reg[1][5] ;
wire \BTB.btag_reg[1][6] ;
wire \BTB.btag_reg[1][7] ;
wire \BTB.btag_reg[1][8] ;
wire \BTB.btag_reg[1][9] ;
wire \BTB.jsnpc_reg[0][0] ;
wire \BTB.jsnpc_reg[0][10] ;
wire \BTB.jsnpc_reg[0][11] ;
wire \BTB.jsnpc_reg[0][12] ;
wire \BTB.jsnpc_reg[0][13] ;
wire \BTB.jsnpc_reg[0][14] ;
wire \BTB.jsnpc_reg[0][15] ;
wire \BTB.jsnpc_reg[0][1] ;
wire \BTB.jsnpc_reg[0][2] ;
wire \BTB.jsnpc_reg[0][3] ;
wire \BTB.jsnpc_reg[0][4] ;
wire \BTB.jsnpc_reg[0][5] ;
wire \BTB.jsnpc_reg[0][6] ;
wire \BTB.jsnpc_reg[0][7] ;
wire \BTB.jsnpc_reg[0][8] ;
wire \BTB.jsnpc_reg[0][9] ;
wire \BTB.jsnpc_reg[1][0] ;
wire \BTB.jsnpc_reg[1][10] ;
wire \BTB.jsnpc_reg[1][11] ;
wire \BTB.jsnpc_reg[1][12] ;
wire \BTB.jsnpc_reg[1][13] ;
wire \BTB.jsnpc_reg[1][14] ;
wire \BTB.jsnpc_reg[1][15] ;
wire \BTB.jsnpc_reg[1][1] ;
wire \BTB.jsnpc_reg[1][2] ;
wire \BTB.jsnpc_reg[1][3] ;
wire \BTB.jsnpc_reg[1][4] ;
wire \BTB.jsnpc_reg[1][5] ;
wire \BTB.jsnpc_reg[1][6] ;
wire \BTB.jsnpc_reg[1][7] ;
wire \BTB.jsnpc_reg[1][8] ;
wire \BTB.jsnpc_reg[1][9] ;
wire \BTB.jtag_reg[0][0] ;
wire \BTB.jtag_reg[0][10] ;
wire \BTB.jtag_reg[0][11] ;
wire \BTB.jtag_reg[0][12] ;
wire \BTB.jtag_reg[0][1] ;
wire \BTB.jtag_reg[0][2] ;
wire \BTB.jtag_reg[0][3] ;
wire \BTB.jtag_reg[0][4] ;
wire \BTB.jtag_reg[0][5] ;
wire \BTB.jtag_reg[0][6] ;
wire \BTB.jtag_reg[0][7] ;
wire \BTB.jtag_reg[0][8] ;
wire \BTB.jtag_reg[0][9] ;
wire \BTB.jtag_reg[1][0] ;
wire \BTB.jtag_reg[1][10] ;
wire \BTB.jtag_reg[1][11] ;
wire \BTB.jtag_reg[1][12] ;
wire \BTB.jtag_reg[1][1] ;
wire \BTB.jtag_reg[1][2] ;
wire \BTB.jtag_reg[1][3] ;
wire \BTB.jtag_reg[1][4] ;
wire \BTB.jtag_reg[1][5] ;
wire \BTB.jtag_reg[1][6] ;
wire \BTB.jtag_reg[1][7] ;
wire \BTB.jtag_reg[1][8] ;
wire \BTB.jtag_reg[1][9] ;
wire CHazarden ;
wire \CLINT.c_axi_arready ;
wire \CLINT.c_axi_arready_$_DFF_P__Q_D ;
wire \CLINT.c_axi_arready_$_NOT__A_Y ;
wire \CLINT.c_axi_rvalid ;
wire \CLINT.c_axi_rvalid_$_NOT__A_Y ;
wire \EXU.dnpc_$_MUX__Y_31_B_$_MUX__B_Y_$_MUX__B_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.dnpc_$_MUX__Y_31_B_$_MUX__B_Y_$_MUX__B_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.funct7_i ;
wire \EXU.gpr_wen_o ;
wire \EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B ;
wire \EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ;
wire \EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_A ;
wire \EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_B ;
wire \EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_B_$_MUX__A_B ;
wire \EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_A ;
wire \EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \EXU.state ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_10_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_10_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_10_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_10_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_11_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_12_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_13_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_14_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_14_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_14_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_14_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_15_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_15_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_15_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_15_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_16_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_17_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_17_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_17_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_17_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_18_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_18_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_18_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_18_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_19_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_20_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_21_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_22_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_23_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_23_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_23_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_23_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_24_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_25_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_25_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_25_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_25_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_26_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_27_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_2_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_3_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_4_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_5_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_6_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_8_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B ;
wire \ICACHE.axi_rvalid ;
wire \ICACHE.axi_rvalid_enable ;
wire \ICACHE.burst_counter_$_DFFE_PP__Q_1_D_$_MUX__Y_B ;
wire \ICACHE.burst_counter_$_DFFE_PP__Q_E_$_ANDNOT__Y_B_$_MUX__Y_A ;
wire \ICACHE.cache_reg[0][10] ;
wire \ICACHE.cache_reg[0][11] ;
wire \ICACHE.cache_reg[0][12] ;
wire \ICACHE.cache_reg[0][13] ;
wire \ICACHE.cache_reg[0][14] ;
wire \ICACHE.cache_reg[0][15] ;
wire \ICACHE.cache_reg[0][16] ;
wire \ICACHE.cache_reg[0][17] ;
wire \ICACHE.cache_reg[0][18] ;
wire \ICACHE.cache_reg[0][19] ;
wire \ICACHE.cache_reg[0][20] ;
wire \ICACHE.cache_reg[0][21] ;
wire \ICACHE.cache_reg[0][22] ;
wire \ICACHE.cache_reg[0][23] ;
wire \ICACHE.cache_reg[0][24] ;
wire \ICACHE.cache_reg[0][25] ;
wire \ICACHE.cache_reg[0][26] ;
wire \ICACHE.cache_reg[0][27] ;
wire \ICACHE.cache_reg[0][28] ;
wire \ICACHE.cache_reg[0][29] ;
wire \ICACHE.cache_reg[0][2] ;
wire \ICACHE.cache_reg[0][30] ;
wire \ICACHE.cache_reg[0][31] ;
wire \ICACHE.cache_reg[0][3] ;
wire \ICACHE.cache_reg[0][4] ;
wire \ICACHE.cache_reg[0][5] ;
wire \ICACHE.cache_reg[0][6] ;
wire \ICACHE.cache_reg[0][7] ;
wire \ICACHE.cache_reg[0][8] ;
wire \ICACHE.cache_reg[0][9] ;
wire \ICACHE.cache_reg[1][10] ;
wire \ICACHE.cache_reg[1][11] ;
wire \ICACHE.cache_reg[1][12] ;
wire \ICACHE.cache_reg[1][13] ;
wire \ICACHE.cache_reg[1][14] ;
wire \ICACHE.cache_reg[1][15] ;
wire \ICACHE.cache_reg[1][16] ;
wire \ICACHE.cache_reg[1][17] ;
wire \ICACHE.cache_reg[1][18] ;
wire \ICACHE.cache_reg[1][19] ;
wire \ICACHE.cache_reg[1][20] ;
wire \ICACHE.cache_reg[1][21] ;
wire \ICACHE.cache_reg[1][22] ;
wire \ICACHE.cache_reg[1][23] ;
wire \ICACHE.cache_reg[1][24] ;
wire \ICACHE.cache_reg[1][25] ;
wire \ICACHE.cache_reg[1][26] ;
wire \ICACHE.cache_reg[1][27] ;
wire \ICACHE.cache_reg[1][28] ;
wire \ICACHE.cache_reg[1][29] ;
wire \ICACHE.cache_reg[1][2] ;
wire \ICACHE.cache_reg[1][30] ;
wire \ICACHE.cache_reg[1][31] ;
wire \ICACHE.cache_reg[1][3] ;
wire \ICACHE.cache_reg[1][4] ;
wire \ICACHE.cache_reg[1][5] ;
wire \ICACHE.cache_reg[1][6] ;
wire \ICACHE.cache_reg[1][7] ;
wire \ICACHE.cache_reg[1][8] ;
wire \ICACHE.cache_reg[1][9] ;
wire \ICACHE.cache_reg[2][10] ;
wire \ICACHE.cache_reg[2][11] ;
wire \ICACHE.cache_reg[2][12] ;
wire \ICACHE.cache_reg[2][13] ;
wire \ICACHE.cache_reg[2][14] ;
wire \ICACHE.cache_reg[2][15] ;
wire \ICACHE.cache_reg[2][16] ;
wire \ICACHE.cache_reg[2][17] ;
wire \ICACHE.cache_reg[2][18] ;
wire \ICACHE.cache_reg[2][19] ;
wire \ICACHE.cache_reg[2][20] ;
wire \ICACHE.cache_reg[2][21] ;
wire \ICACHE.cache_reg[2][22] ;
wire \ICACHE.cache_reg[2][23] ;
wire \ICACHE.cache_reg[2][24] ;
wire \ICACHE.cache_reg[2][25] ;
wire \ICACHE.cache_reg[2][26] ;
wire \ICACHE.cache_reg[2][27] ;
wire \ICACHE.cache_reg[2][28] ;
wire \ICACHE.cache_reg[2][29] ;
wire \ICACHE.cache_reg[2][2] ;
wire \ICACHE.cache_reg[2][30] ;
wire \ICACHE.cache_reg[2][31] ;
wire \ICACHE.cache_reg[2][3] ;
wire \ICACHE.cache_reg[2][4] ;
wire \ICACHE.cache_reg[2][5] ;
wire \ICACHE.cache_reg[2][6] ;
wire \ICACHE.cache_reg[2][7] ;
wire \ICACHE.cache_reg[2][8] ;
wire \ICACHE.cache_reg[2][9] ;
wire \ICACHE.cache_reg[3][10] ;
wire \ICACHE.cache_reg[3][11] ;
wire \ICACHE.cache_reg[3][12] ;
wire \ICACHE.cache_reg[3][13] ;
wire \ICACHE.cache_reg[3][14] ;
wire \ICACHE.cache_reg[3][15] ;
wire \ICACHE.cache_reg[3][16] ;
wire \ICACHE.cache_reg[3][17] ;
wire \ICACHE.cache_reg[3][18] ;
wire \ICACHE.cache_reg[3][19] ;
wire \ICACHE.cache_reg[3][20] ;
wire \ICACHE.cache_reg[3][21] ;
wire \ICACHE.cache_reg[3][22] ;
wire \ICACHE.cache_reg[3][23] ;
wire \ICACHE.cache_reg[3][24] ;
wire \ICACHE.cache_reg[3][25] ;
wire \ICACHE.cache_reg[3][26] ;
wire \ICACHE.cache_reg[3][27] ;
wire \ICACHE.cache_reg[3][28] ;
wire \ICACHE.cache_reg[3][29] ;
wire \ICACHE.cache_reg[3][2] ;
wire \ICACHE.cache_reg[3][30] ;
wire \ICACHE.cache_reg[3][31] ;
wire \ICACHE.cache_reg[3][3] ;
wire \ICACHE.cache_reg[3][4] ;
wire \ICACHE.cache_reg[3][5] ;
wire \ICACHE.cache_reg[3][6] ;
wire \ICACHE.cache_reg[3][7] ;
wire \ICACHE.cache_reg[3][8] ;
wire \ICACHE.cache_reg[3][9] ;
wire \ICACHE.cache_reg[4][10] ;
wire \ICACHE.cache_reg[4][11] ;
wire \ICACHE.cache_reg[4][12] ;
wire \ICACHE.cache_reg[4][13] ;
wire \ICACHE.cache_reg[4][14] ;
wire \ICACHE.cache_reg[4][15] ;
wire \ICACHE.cache_reg[4][16] ;
wire \ICACHE.cache_reg[4][17] ;
wire \ICACHE.cache_reg[4][18] ;
wire \ICACHE.cache_reg[4][19] ;
wire \ICACHE.cache_reg[4][20] ;
wire \ICACHE.cache_reg[4][21] ;
wire \ICACHE.cache_reg[4][22] ;
wire \ICACHE.cache_reg[4][23] ;
wire \ICACHE.cache_reg[4][24] ;
wire \ICACHE.cache_reg[4][25] ;
wire \ICACHE.cache_reg[4][26] ;
wire \ICACHE.cache_reg[4][27] ;
wire \ICACHE.cache_reg[4][28] ;
wire \ICACHE.cache_reg[4][29] ;
wire \ICACHE.cache_reg[4][2] ;
wire \ICACHE.cache_reg[4][30] ;
wire \ICACHE.cache_reg[4][31] ;
wire \ICACHE.cache_reg[4][3] ;
wire \ICACHE.cache_reg[4][4] ;
wire \ICACHE.cache_reg[4][5] ;
wire \ICACHE.cache_reg[4][6] ;
wire \ICACHE.cache_reg[4][7] ;
wire \ICACHE.cache_reg[4][8] ;
wire \ICACHE.cache_reg[4][9] ;
wire \ICACHE.cache_reg[5][10] ;
wire \ICACHE.cache_reg[5][11] ;
wire \ICACHE.cache_reg[5][12] ;
wire \ICACHE.cache_reg[5][13] ;
wire \ICACHE.cache_reg[5][14] ;
wire \ICACHE.cache_reg[5][15] ;
wire \ICACHE.cache_reg[5][16] ;
wire \ICACHE.cache_reg[5][17] ;
wire \ICACHE.cache_reg[5][18] ;
wire \ICACHE.cache_reg[5][19] ;
wire \ICACHE.cache_reg[5][20] ;
wire \ICACHE.cache_reg[5][21] ;
wire \ICACHE.cache_reg[5][22] ;
wire \ICACHE.cache_reg[5][23] ;
wire \ICACHE.cache_reg[5][24] ;
wire \ICACHE.cache_reg[5][25] ;
wire \ICACHE.cache_reg[5][26] ;
wire \ICACHE.cache_reg[5][27] ;
wire \ICACHE.cache_reg[5][28] ;
wire \ICACHE.cache_reg[5][29] ;
wire \ICACHE.cache_reg[5][2] ;
wire \ICACHE.cache_reg[5][30] ;
wire \ICACHE.cache_reg[5][31] ;
wire \ICACHE.cache_reg[5][3] ;
wire \ICACHE.cache_reg[5][4] ;
wire \ICACHE.cache_reg[5][5] ;
wire \ICACHE.cache_reg[5][6] ;
wire \ICACHE.cache_reg[5][7] ;
wire \ICACHE.cache_reg[5][8] ;
wire \ICACHE.cache_reg[5][9] ;
wire \ICACHE.cache_reg[6][10] ;
wire \ICACHE.cache_reg[6][11] ;
wire \ICACHE.cache_reg[6][12] ;
wire \ICACHE.cache_reg[6][13] ;
wire \ICACHE.cache_reg[6][14] ;
wire \ICACHE.cache_reg[6][15] ;
wire \ICACHE.cache_reg[6][16] ;
wire \ICACHE.cache_reg[6][17] ;
wire \ICACHE.cache_reg[6][18] ;
wire \ICACHE.cache_reg[6][19] ;
wire \ICACHE.cache_reg[6][20] ;
wire \ICACHE.cache_reg[6][21] ;
wire \ICACHE.cache_reg[6][22] ;
wire \ICACHE.cache_reg[6][23] ;
wire \ICACHE.cache_reg[6][24] ;
wire \ICACHE.cache_reg[6][25] ;
wire \ICACHE.cache_reg[6][26] ;
wire \ICACHE.cache_reg[6][27] ;
wire \ICACHE.cache_reg[6][28] ;
wire \ICACHE.cache_reg[6][29] ;
wire \ICACHE.cache_reg[6][2] ;
wire \ICACHE.cache_reg[6][30] ;
wire \ICACHE.cache_reg[6][31] ;
wire \ICACHE.cache_reg[6][3] ;
wire \ICACHE.cache_reg[6][4] ;
wire \ICACHE.cache_reg[6][5] ;
wire \ICACHE.cache_reg[6][6] ;
wire \ICACHE.cache_reg[6][7] ;
wire \ICACHE.cache_reg[6][8] ;
wire \ICACHE.cache_reg[6][9] ;
wire \ICACHE.cache_reg[7][10] ;
wire \ICACHE.cache_reg[7][11] ;
wire \ICACHE.cache_reg[7][12] ;
wire \ICACHE.cache_reg[7][13] ;
wire \ICACHE.cache_reg[7][14] ;
wire \ICACHE.cache_reg[7][15] ;
wire \ICACHE.cache_reg[7][16] ;
wire \ICACHE.cache_reg[7][17] ;
wire \ICACHE.cache_reg[7][18] ;
wire \ICACHE.cache_reg[7][19] ;
wire \ICACHE.cache_reg[7][20] ;
wire \ICACHE.cache_reg[7][21] ;
wire \ICACHE.cache_reg[7][22] ;
wire \ICACHE.cache_reg[7][23] ;
wire \ICACHE.cache_reg[7][24] ;
wire \ICACHE.cache_reg[7][25] ;
wire \ICACHE.cache_reg[7][26] ;
wire \ICACHE.cache_reg[7][27] ;
wire \ICACHE.cache_reg[7][28] ;
wire \ICACHE.cache_reg[7][29] ;
wire \ICACHE.cache_reg[7][2] ;
wire \ICACHE.cache_reg[7][30] ;
wire \ICACHE.cache_reg[7][31] ;
wire \ICACHE.cache_reg[7][3] ;
wire \ICACHE.cache_reg[7][4] ;
wire \ICACHE.cache_reg[7][5] ;
wire \ICACHE.cache_reg[7][6] ;
wire \ICACHE.cache_reg[7][7] ;
wire \ICACHE.cache_reg[7][8] ;
wire \ICACHE.cache_reg[7][9] ;
wire \ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \ICACHE.m_axi_arready ;
wire \ICACHE.m_axi_arvalid ;
wire \ICACHE.m_axi_rready ;
wire \ICACHE.s_axi_arvalid ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_10_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_11_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_12_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_13_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_14_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_15_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_16_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_17_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_18_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_19_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_1_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_20_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_21_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_22_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_23_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_24_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_25_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_26_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_27_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_28_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_29_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_2_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_3_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_4_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_5_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_6_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_7_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_8_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_9_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rdata_$_ANDNOT__Y_B_$_MUX__Y_A ;
wire \ICACHE.s_axi_rready ;
wire \ICACHE.state_$_MUX__S_A ;
wire \ICACHE.state_$_MUX__S_B ;
wire \ICACHE.tag_reg[0][0] ;
wire \ICACHE.tag_reg[0][10] ;
wire \ICACHE.tag_reg[0][1] ;
wire \ICACHE.tag_reg[0][2] ;
wire \ICACHE.tag_reg[0][3] ;
wire \ICACHE.tag_reg[0][4] ;
wire \ICACHE.tag_reg[0][5] ;
wire \ICACHE.tag_reg[0][6] ;
wire \ICACHE.tag_reg[0][7] ;
wire \ICACHE.tag_reg[0][8] ;
wire \ICACHE.tag_reg[0][9] ;
wire \ICACHE.tag_reg[1][0] ;
wire \ICACHE.tag_reg[1][10] ;
wire \ICACHE.tag_reg[1][1] ;
wire \ICACHE.tag_reg[1][2] ;
wire \ICACHE.tag_reg[1][3] ;
wire \ICACHE.tag_reg[1][4] ;
wire \ICACHE.tag_reg[1][5] ;
wire \ICACHE.tag_reg[1][6] ;
wire \ICACHE.tag_reg[1][7] ;
wire \ICACHE.tag_reg[1][8] ;
wire \ICACHE.tag_reg[1][9] ;
wire \ICACHE.valid_reg[0][0] ;
wire \ICACHE.valid_reg[0][1] ;
wire \ICACHE.valid_reg[0][2] ;
wire \ICACHE.valid_reg[0][3] ;
wire \ICACHE.valid_reg[1][0] ;
wire \ICACHE.valid_reg[1][1] ;
wire \ICACHE.valid_reg[1][2] ;
wire \ICACHE.valid_reg[1][3] ;
wire \IDU.if_valid_i ;
wire \IDU.imm_$_NOR__Y_10_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_10_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_1_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_2_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_3_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_4_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_5_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_6_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_7_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_7_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_8_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_8_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_9_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_9_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \IDU.imm_$_NOR__Y_A_$_MUX__Y_B ;
wire \IDU.ls_valid_o ;
wire \IDU.ls_valid_o_$_DFFE_PP__Q_D_$_ANDNOT__Y_B_$_NOR__Y_B_$_ANDNOT__Y_A ;
wire \IDU.ls_valid_o_$_DFFE_PP__Q_E_$_OR__Y_B ;
wire \IDU.prevalid ;
wire \IDU.prevalid_$_NAND__B_A_$_ANDNOT__Y_B ;
wire \IDU.state ;
wire \IDU.updata ;
wire \IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y ;
wire \IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ;
wire \IFU.state ;
wire \IFU.state_$_NOT__A_Y ;
wire \IFU.updata ;
wire \LSU.axi_state_$_DFF_P__Q_1_D ;
wire \LSU.axi_state_$_DFF_P__Q_2_D ;
wire \LSU.axi_state_$_DFF_P__Q_D ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_10_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_10_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_11_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_11_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_14_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_14_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_15_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_15_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_16_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_16_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_17_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_18_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_19_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_20_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_21_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_B_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_B_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_2_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_2_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_4_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_4_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_5_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_5_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_7_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_7_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_8_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_8_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A ;
wire \LSU.ls_addr_i_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \LSU.ls_axi_arvalid ;
wire \LSU.ls_axi_arvalid_$_SDFFE_PP0P__Q_D ;
wire \LSU.ls_axi_awvalid ;
wire \LSU.ls_axi_awvalid_$_NOT__A_Y ;
wire \LSU.ls_axi_bready ;
wire \LSU.ls_axi_rready ;
wire \LSU.ls_axi_rready_$_ANDNOT__A_Y ;
wire \LSU.ls_axi_rready_$_NOT__A_Y ;
wire \LSU.ls_axi_wlast ;
wire \LSU.ls_axi_wlast_$_DFFE_PP__Q_D ;
wire \LSU.ls_axi_wvalid ;
wire \LSU.ls_axi_wvalid_$_NOT__A_Y ;
wire \LSU.ls_read_done ;
wire \LSU.ls_read_done_$_OR__B_Y_$_ORNOT__A_Y_$_ANDNOT__A_Y_$_OR__A_1_B ;
wire \LSU.ls_wdata_i_$_MUX__Y_16_A_$_ANDNOT__Y_B ;
wire \LSU.ls_wdata_i_$_MUX__Y_17_A_$_ANDNOT__Y_B ;
wire \LSU.ls_wdata_i_$_MUX__Y_18_A_$_ANDNOT__Y_B ;
wire \LSU.ls_wdata_i_$_MUX__Y_19_A_$_ANDNOT__Y_B ;
wire \LSU.ls_wdata_i_$_MUX__Y_20_A_$_ANDNOT__Y_B ;
wire \LSU.ls_wdata_i_$_MUX__Y_21_A_$_ANDNOT__Y_B ;
wire \LSU.ls_wdata_i_$_MUX__Y_22_A_$_ANDNOT__Y_B ;
wire \LSU.ls_wdata_i_$_MUX__Y_23_A_$_ANDNOT__Y_B ;
wire \RFU.rf[10][0] ;
wire \RFU.rf[10][10] ;
wire \RFU.rf[10][11] ;
wire \RFU.rf[10][12] ;
wire \RFU.rf[10][13] ;
wire \RFU.rf[10][14] ;
wire \RFU.rf[10][15] ;
wire \RFU.rf[10][16] ;
wire \RFU.rf[10][17] ;
wire \RFU.rf[10][18] ;
wire \RFU.rf[10][19] ;
wire \RFU.rf[10][1] ;
wire \RFU.rf[10][20] ;
wire \RFU.rf[10][21] ;
wire \RFU.rf[10][22] ;
wire \RFU.rf[10][23] ;
wire \RFU.rf[10][24] ;
wire \RFU.rf[10][25] ;
wire \RFU.rf[10][26] ;
wire \RFU.rf[10][27] ;
wire \RFU.rf[10][28] ;
wire \RFU.rf[10][29] ;
wire \RFU.rf[10][2] ;
wire \RFU.rf[10][30] ;
wire \RFU.rf[10][31] ;
wire \RFU.rf[10][3] ;
wire \RFU.rf[10][4] ;
wire \RFU.rf[10][5] ;
wire \RFU.rf[10][6] ;
wire \RFU.rf[10][7] ;
wire \RFU.rf[10][8] ;
wire \RFU.rf[10][9] ;
wire \RFU.rf[11][0] ;
wire \RFU.rf[11][10] ;
wire \RFU.rf[11][11] ;
wire \RFU.rf[11][12] ;
wire \RFU.rf[11][13] ;
wire \RFU.rf[11][14] ;
wire \RFU.rf[11][15] ;
wire \RFU.rf[11][16] ;
wire \RFU.rf[11][17] ;
wire \RFU.rf[11][18] ;
wire \RFU.rf[11][19] ;
wire \RFU.rf[11][1] ;
wire \RFU.rf[11][20] ;
wire \RFU.rf[11][21] ;
wire \RFU.rf[11][22] ;
wire \RFU.rf[11][23] ;
wire \RFU.rf[11][24] ;
wire \RFU.rf[11][25] ;
wire \RFU.rf[11][26] ;
wire \RFU.rf[11][27] ;
wire \RFU.rf[11][28] ;
wire \RFU.rf[11][29] ;
wire \RFU.rf[11][2] ;
wire \RFU.rf[11][30] ;
wire \RFU.rf[11][31] ;
wire \RFU.rf[11][3] ;
wire \RFU.rf[11][4] ;
wire \RFU.rf[11][5] ;
wire \RFU.rf[11][6] ;
wire \RFU.rf[11][7] ;
wire \RFU.rf[11][8] ;
wire \RFU.rf[11][9] ;
wire \RFU.rf[12][0] ;
wire \RFU.rf[12][10] ;
wire \RFU.rf[12][11] ;
wire \RFU.rf[12][12] ;
wire \RFU.rf[12][13] ;
wire \RFU.rf[12][14] ;
wire \RFU.rf[12][15] ;
wire \RFU.rf[12][16] ;
wire \RFU.rf[12][17] ;
wire \RFU.rf[12][18] ;
wire \RFU.rf[12][19] ;
wire \RFU.rf[12][1] ;
wire \RFU.rf[12][20] ;
wire \RFU.rf[12][21] ;
wire \RFU.rf[12][22] ;
wire \RFU.rf[12][23] ;
wire \RFU.rf[12][24] ;
wire \RFU.rf[12][25] ;
wire \RFU.rf[12][26] ;
wire \RFU.rf[12][27] ;
wire \RFU.rf[12][28] ;
wire \RFU.rf[12][29] ;
wire \RFU.rf[12][2] ;
wire \RFU.rf[12][30] ;
wire \RFU.rf[12][31] ;
wire \RFU.rf[12][3] ;
wire \RFU.rf[12][4] ;
wire \RFU.rf[12][5] ;
wire \RFU.rf[12][6] ;
wire \RFU.rf[12][7] ;
wire \RFU.rf[12][8] ;
wire \RFU.rf[12][9] ;
wire \RFU.rf[13][0] ;
wire \RFU.rf[13][10] ;
wire \RFU.rf[13][11] ;
wire \RFU.rf[13][12] ;
wire \RFU.rf[13][13] ;
wire \RFU.rf[13][14] ;
wire \RFU.rf[13][15] ;
wire \RFU.rf[13][16] ;
wire \RFU.rf[13][17] ;
wire \RFU.rf[13][18] ;
wire \RFU.rf[13][19] ;
wire \RFU.rf[13][1] ;
wire \RFU.rf[13][20] ;
wire \RFU.rf[13][21] ;
wire \RFU.rf[13][22] ;
wire \RFU.rf[13][23] ;
wire \RFU.rf[13][24] ;
wire \RFU.rf[13][25] ;
wire \RFU.rf[13][26] ;
wire \RFU.rf[13][27] ;
wire \RFU.rf[13][28] ;
wire \RFU.rf[13][29] ;
wire \RFU.rf[13][2] ;
wire \RFU.rf[13][30] ;
wire \RFU.rf[13][31] ;
wire \RFU.rf[13][3] ;
wire \RFU.rf[13][4] ;
wire \RFU.rf[13][5] ;
wire \RFU.rf[13][6] ;
wire \RFU.rf[13][7] ;
wire \RFU.rf[13][8] ;
wire \RFU.rf[13][9] ;
wire \RFU.rf[14][0] ;
wire \RFU.rf[14][10] ;
wire \RFU.rf[14][11] ;
wire \RFU.rf[14][12] ;
wire \RFU.rf[14][13] ;
wire \RFU.rf[14][14] ;
wire \RFU.rf[14][15] ;
wire \RFU.rf[14][16] ;
wire \RFU.rf[14][17] ;
wire \RFU.rf[14][18] ;
wire \RFU.rf[14][19] ;
wire \RFU.rf[14][1] ;
wire \RFU.rf[14][20] ;
wire \RFU.rf[14][21] ;
wire \RFU.rf[14][22] ;
wire \RFU.rf[14][23] ;
wire \RFU.rf[14][24] ;
wire \RFU.rf[14][25] ;
wire \RFU.rf[14][26] ;
wire \RFU.rf[14][27] ;
wire \RFU.rf[14][28] ;
wire \RFU.rf[14][29] ;
wire \RFU.rf[14][2] ;
wire \RFU.rf[14][30] ;
wire \RFU.rf[14][31] ;
wire \RFU.rf[14][3] ;
wire \RFU.rf[14][4] ;
wire \RFU.rf[14][5] ;
wire \RFU.rf[14][6] ;
wire \RFU.rf[14][7] ;
wire \RFU.rf[14][8] ;
wire \RFU.rf[14][9] ;
wire \RFU.rf[15][0] ;
wire \RFU.rf[15][10] ;
wire \RFU.rf[15][11] ;
wire \RFU.rf[15][12] ;
wire \RFU.rf[15][13] ;
wire \RFU.rf[15][14] ;
wire \RFU.rf[15][15] ;
wire \RFU.rf[15][16] ;
wire \RFU.rf[15][17] ;
wire \RFU.rf[15][18] ;
wire \RFU.rf[15][19] ;
wire \RFU.rf[15][1] ;
wire \RFU.rf[15][20] ;
wire \RFU.rf[15][21] ;
wire \RFU.rf[15][22] ;
wire \RFU.rf[15][23] ;
wire \RFU.rf[15][24] ;
wire \RFU.rf[15][25] ;
wire \RFU.rf[15][26] ;
wire \RFU.rf[15][27] ;
wire \RFU.rf[15][28] ;
wire \RFU.rf[15][29] ;
wire \RFU.rf[15][2] ;
wire \RFU.rf[15][30] ;
wire \RFU.rf[15][31] ;
wire \RFU.rf[15][3] ;
wire \RFU.rf[15][4] ;
wire \RFU.rf[15][5] ;
wire \RFU.rf[15][6] ;
wire \RFU.rf[15][7] ;
wire \RFU.rf[15][8] ;
wire \RFU.rf[15][9] ;
wire \RFU.rf[1][0] ;
wire \RFU.rf[1][10] ;
wire \RFU.rf[1][11] ;
wire \RFU.rf[1][12] ;
wire \RFU.rf[1][13] ;
wire \RFU.rf[1][14] ;
wire \RFU.rf[1][15] ;
wire \RFU.rf[1][16] ;
wire \RFU.rf[1][17] ;
wire \RFU.rf[1][18] ;
wire \RFU.rf[1][19] ;
wire \RFU.rf[1][1] ;
wire \RFU.rf[1][20] ;
wire \RFU.rf[1][21] ;
wire \RFU.rf[1][22] ;
wire \RFU.rf[1][23] ;
wire \RFU.rf[1][24] ;
wire \RFU.rf[1][25] ;
wire \RFU.rf[1][26] ;
wire \RFU.rf[1][27] ;
wire \RFU.rf[1][28] ;
wire \RFU.rf[1][29] ;
wire \RFU.rf[1][2] ;
wire \RFU.rf[1][30] ;
wire \RFU.rf[1][31] ;
wire \RFU.rf[1][3] ;
wire \RFU.rf[1][4] ;
wire \RFU.rf[1][5] ;
wire \RFU.rf[1][6] ;
wire \RFU.rf[1][7] ;
wire \RFU.rf[1][8] ;
wire \RFU.rf[1][9] ;
wire \RFU.rf[2][0] ;
wire \RFU.rf[2][10] ;
wire \RFU.rf[2][11] ;
wire \RFU.rf[2][12] ;
wire \RFU.rf[2][13] ;
wire \RFU.rf[2][14] ;
wire \RFU.rf[2][15] ;
wire \RFU.rf[2][16] ;
wire \RFU.rf[2][17] ;
wire \RFU.rf[2][18] ;
wire \RFU.rf[2][19] ;
wire \RFU.rf[2][1] ;
wire \RFU.rf[2][20] ;
wire \RFU.rf[2][21] ;
wire \RFU.rf[2][22] ;
wire \RFU.rf[2][23] ;
wire \RFU.rf[2][24] ;
wire \RFU.rf[2][25] ;
wire \RFU.rf[2][26] ;
wire \RFU.rf[2][27] ;
wire \RFU.rf[2][28] ;
wire \RFU.rf[2][29] ;
wire \RFU.rf[2][2] ;
wire \RFU.rf[2][30] ;
wire \RFU.rf[2][31] ;
wire \RFU.rf[2][3] ;
wire \RFU.rf[2][4] ;
wire \RFU.rf[2][5] ;
wire \RFU.rf[2][6] ;
wire \RFU.rf[2][7] ;
wire \RFU.rf[2][8] ;
wire \RFU.rf[2][9] ;
wire \RFU.rf[3][0] ;
wire \RFU.rf[3][10] ;
wire \RFU.rf[3][11] ;
wire \RFU.rf[3][12] ;
wire \RFU.rf[3][13] ;
wire \RFU.rf[3][14] ;
wire \RFU.rf[3][15] ;
wire \RFU.rf[3][16] ;
wire \RFU.rf[3][17] ;
wire \RFU.rf[3][18] ;
wire \RFU.rf[3][19] ;
wire \RFU.rf[3][1] ;
wire \RFU.rf[3][20] ;
wire \RFU.rf[3][21] ;
wire \RFU.rf[3][22] ;
wire \RFU.rf[3][23] ;
wire \RFU.rf[3][24] ;
wire \RFU.rf[3][25] ;
wire \RFU.rf[3][26] ;
wire \RFU.rf[3][27] ;
wire \RFU.rf[3][28] ;
wire \RFU.rf[3][29] ;
wire \RFU.rf[3][2] ;
wire \RFU.rf[3][30] ;
wire \RFU.rf[3][31] ;
wire \RFU.rf[3][3] ;
wire \RFU.rf[3][4] ;
wire \RFU.rf[3][5] ;
wire \RFU.rf[3][6] ;
wire \RFU.rf[3][7] ;
wire \RFU.rf[3][8] ;
wire \RFU.rf[3][9] ;
wire \RFU.rf[4][0] ;
wire \RFU.rf[4][10] ;
wire \RFU.rf[4][11] ;
wire \RFU.rf[4][12] ;
wire \RFU.rf[4][13] ;
wire \RFU.rf[4][14] ;
wire \RFU.rf[4][15] ;
wire \RFU.rf[4][16] ;
wire \RFU.rf[4][17] ;
wire \RFU.rf[4][18] ;
wire \RFU.rf[4][19] ;
wire \RFU.rf[4][1] ;
wire \RFU.rf[4][20] ;
wire \RFU.rf[4][21] ;
wire \RFU.rf[4][22] ;
wire \RFU.rf[4][23] ;
wire \RFU.rf[4][24] ;
wire \RFU.rf[4][25] ;
wire \RFU.rf[4][26] ;
wire \RFU.rf[4][27] ;
wire \RFU.rf[4][28] ;
wire \RFU.rf[4][29] ;
wire \RFU.rf[4][2] ;
wire \RFU.rf[4][30] ;
wire \RFU.rf[4][31] ;
wire \RFU.rf[4][3] ;
wire \RFU.rf[4][4] ;
wire \RFU.rf[4][5] ;
wire \RFU.rf[4][6] ;
wire \RFU.rf[4][7] ;
wire \RFU.rf[4][8] ;
wire \RFU.rf[4][9] ;
wire \RFU.rf[5][0] ;
wire \RFU.rf[5][10] ;
wire \RFU.rf[5][11] ;
wire \RFU.rf[5][12] ;
wire \RFU.rf[5][13] ;
wire \RFU.rf[5][14] ;
wire \RFU.rf[5][15] ;
wire \RFU.rf[5][16] ;
wire \RFU.rf[5][17] ;
wire \RFU.rf[5][18] ;
wire \RFU.rf[5][19] ;
wire \RFU.rf[5][1] ;
wire \RFU.rf[5][20] ;
wire \RFU.rf[5][21] ;
wire \RFU.rf[5][22] ;
wire \RFU.rf[5][23] ;
wire \RFU.rf[5][24] ;
wire \RFU.rf[5][25] ;
wire \RFU.rf[5][26] ;
wire \RFU.rf[5][27] ;
wire \RFU.rf[5][28] ;
wire \RFU.rf[5][29] ;
wire \RFU.rf[5][2] ;
wire \RFU.rf[5][30] ;
wire \RFU.rf[5][31] ;
wire \RFU.rf[5][3] ;
wire \RFU.rf[5][4] ;
wire \RFU.rf[5][5] ;
wire \RFU.rf[5][6] ;
wire \RFU.rf[5][7] ;
wire \RFU.rf[5][8] ;
wire \RFU.rf[5][9] ;
wire \RFU.rf[6][0] ;
wire \RFU.rf[6][10] ;
wire \RFU.rf[6][11] ;
wire \RFU.rf[6][12] ;
wire \RFU.rf[6][13] ;
wire \RFU.rf[6][14] ;
wire \RFU.rf[6][15] ;
wire \RFU.rf[6][16] ;
wire \RFU.rf[6][17] ;
wire \RFU.rf[6][18] ;
wire \RFU.rf[6][19] ;
wire \RFU.rf[6][1] ;
wire \RFU.rf[6][20] ;
wire \RFU.rf[6][21] ;
wire \RFU.rf[6][22] ;
wire \RFU.rf[6][23] ;
wire \RFU.rf[6][24] ;
wire \RFU.rf[6][25] ;
wire \RFU.rf[6][26] ;
wire \RFU.rf[6][27] ;
wire \RFU.rf[6][28] ;
wire \RFU.rf[6][29] ;
wire \RFU.rf[6][2] ;
wire \RFU.rf[6][30] ;
wire \RFU.rf[6][31] ;
wire \RFU.rf[6][3] ;
wire \RFU.rf[6][4] ;
wire \RFU.rf[6][5] ;
wire \RFU.rf[6][6] ;
wire \RFU.rf[6][7] ;
wire \RFU.rf[6][8] ;
wire \RFU.rf[6][9] ;
wire \RFU.rf[7][0] ;
wire \RFU.rf[7][10] ;
wire \RFU.rf[7][11] ;
wire \RFU.rf[7][12] ;
wire \RFU.rf[7][13] ;
wire \RFU.rf[7][14] ;
wire \RFU.rf[7][15] ;
wire \RFU.rf[7][16] ;
wire \RFU.rf[7][17] ;
wire \RFU.rf[7][18] ;
wire \RFU.rf[7][19] ;
wire \RFU.rf[7][1] ;
wire \RFU.rf[7][20] ;
wire \RFU.rf[7][21] ;
wire \RFU.rf[7][22] ;
wire \RFU.rf[7][23] ;
wire \RFU.rf[7][24] ;
wire \RFU.rf[7][25] ;
wire \RFU.rf[7][26] ;
wire \RFU.rf[7][27] ;
wire \RFU.rf[7][28] ;
wire \RFU.rf[7][29] ;
wire \RFU.rf[7][2] ;
wire \RFU.rf[7][30] ;
wire \RFU.rf[7][31] ;
wire \RFU.rf[7][3] ;
wire \RFU.rf[7][4] ;
wire \RFU.rf[7][5] ;
wire \RFU.rf[7][6] ;
wire \RFU.rf[7][7] ;
wire \RFU.rf[7][8] ;
wire \RFU.rf[7][9] ;
wire \RFU.rf[8][0] ;
wire \RFU.rf[8][10] ;
wire \RFU.rf[8][11] ;
wire \RFU.rf[8][12] ;
wire \RFU.rf[8][13] ;
wire \RFU.rf[8][14] ;
wire \RFU.rf[8][15] ;
wire \RFU.rf[8][16] ;
wire \RFU.rf[8][17] ;
wire \RFU.rf[8][18] ;
wire \RFU.rf[8][19] ;
wire \RFU.rf[8][1] ;
wire \RFU.rf[8][20] ;
wire \RFU.rf[8][21] ;
wire \RFU.rf[8][22] ;
wire \RFU.rf[8][23] ;
wire \RFU.rf[8][24] ;
wire \RFU.rf[8][25] ;
wire \RFU.rf[8][26] ;
wire \RFU.rf[8][27] ;
wire \RFU.rf[8][28] ;
wire \RFU.rf[8][29] ;
wire \RFU.rf[8][2] ;
wire \RFU.rf[8][30] ;
wire \RFU.rf[8][31] ;
wire \RFU.rf[8][3] ;
wire \RFU.rf[8][4] ;
wire \RFU.rf[8][5] ;
wire \RFU.rf[8][6] ;
wire \RFU.rf[8][7] ;
wire \RFU.rf[8][8] ;
wire \RFU.rf[8][9] ;
wire \RFU.rf[9][0] ;
wire \RFU.rf[9][10] ;
wire \RFU.rf[9][11] ;
wire \RFU.rf[9][12] ;
wire \RFU.rf[9][13] ;
wire \RFU.rf[9][14] ;
wire \RFU.rf[9][15] ;
wire \RFU.rf[9][16] ;
wire \RFU.rf[9][17] ;
wire \RFU.rf[9][18] ;
wire \RFU.rf[9][19] ;
wire \RFU.rf[9][1] ;
wire \RFU.rf[9][20] ;
wire \RFU.rf[9][21] ;
wire \RFU.rf[9][22] ;
wire \RFU.rf[9][23] ;
wire \RFU.rf[9][24] ;
wire \RFU.rf[9][25] ;
wire \RFU.rf[9][26] ;
wire \RFU.rf[9][27] ;
wire \RFU.rf[9][28] ;
wire \RFU.rf[9][29] ;
wire \RFU.rf[9][2] ;
wire \RFU.rf[9][30] ;
wire \RFU.rf[9][31] ;
wire \RFU.rf[9][3] ;
wire \RFU.rf[9][4] ;
wire \RFU.rf[9][5] ;
wire \RFU.rf[9][6] ;
wire \RFU.rf[9][7] ;
wire \RFU.rf[9][8] ;
wire \RFU.rf[9][9] ;
wire \Xbar.state_$_DFF_P__Q_1_D ;
wire \Xbar.state_$_DFF_P__Q_2_D ;
wire \Xbar.state_$_DFF_P__Q_D ;
wire clock ;
wire io_interrupt ;
wire io_master_arready ;
wire io_master_arsize_$_ANDNOT__Y_1_B_$_OR__Y_A_$_OR__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_AND__Y_B_$_OR__Y_B ;
wire io_master_arvalid ;
wire io_master_arvalid_$_ANDNOT__Y_B_$_MUX__Y_A ;
wire io_master_arvalid_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_rlast ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_wlast ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_rlast ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_wlast ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire prepc_$_ANDNOT__Y_10_B_$_XOR__Y_B_$_XOR__Y_B ;
wire prepc_$_ANDNOT__Y_12_B_$_XOR__Y_B_$_XOR__Y_B ;
wire prepc_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_B ;
wire prepc_$_ANDNOT__Y_6_B_$_XOR__Y_B_$_XOR__Y_B ;
wire prepc_$_ANDNOT__Y_8_B_$_XOR__Y_B_$_XOR__Y_B ;
wire reset ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire [12:0] \BTB.btag ;
wire [12:0] \BTB.btag_pre ;
wire [31:0] \BTB.pc_i ;
wire [31:0] \BTB.prepc_tag_i ;
wire [31:0] \CLINT.c_axi_rdata ;
wire [63:0] \CLINT.mtime ;
wire [0:0] \CLINT.mtime_$_SDFF_PP0__Q_63_D ;
wire [1:0] \EXU.add_pc_4 ;
wire [1:0] \EXU.counter ;
wire [0:0] \EXU.counter_$_SDFFE_PP0N__Q_1_D ;
wire [3:0] \EXU.csrs_wen_o ;
wire [31:0] \EXU.dnpc_o ;
wire [2:0] \EXU.funct3_i ;
wire [31:0] \EXU.imm_i ;
wire [31:0] \EXU.ls_rdata_i ;
wire [31:0] \EXU.mcause_i ;
wire [31:0] \EXU.mepc_i ;
wire [31:0] \EXU.mstatus_i ;
wire [31:0] \EXU.mtvec_i ;
wire [4:0] \EXU.op_i ;
wire [31:0] \EXU.pc_i ;
wire [31:0] \EXU.r1_i ;
wire [31:0] \EXU.r2_i ;
wire [3:0] \EXU.rd_i ;
wire [3:0] \EXU.rd_o ;
wire [31:0] \EXU.xrd_o ;
wire [1:0] \ICACHE.burst_counter ;
wire [31:0] \ICACHE.s_axi_araddr ;
wire [3:0] \ICACHE.s_axi_arlen ;
wire [15:0] \ICACHE.tag_check ;
wire [2:0] \IDU.funct3 ;
wire [6:0] \IDU.funct7 ;
wire [11:0] \IDU.immB ;
wire [4:0] \IDU.immI ;
wire [19:0] \IDU.immJ ;
wire [6:0] \IDU.inst_i ;
wire [2:0] \LSU.axi_state ;
wire [31:0] \LSU.ls_axi_araddr ;
wire [31:0] \LSU.ls_axi_awaddr ;
wire [31:0] \LSU.ls_axi_wdata ;
wire [2:0] \Xbar.state ;
wire [31:0] io_master_araddr ;
wire [1:0] io_master_arburst ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [31:0] io_master_awaddr ;
wire [1:0] io_master_awburst ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [3:0] io_master_bid ;
wire [1:0] io_master_bresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [31:0] io_slave_araddr ;
wire [1:0] io_slave_arburst ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [31:0] io_slave_awaddr ;
wire [1:0] io_slave_awburst ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [3:0] io_slave_bid ;
wire [1:0] io_slave_bresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;

assign \io_master_arid [0] = \io_master_arburst [1] ;
assign \io_master_arid [1] = \io_master_arburst [1] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arlen [3] ;
assign \io_master_arlen [5] = \io_master_arlen [3] ;
assign \io_master_arlen [6] = \io_master_arlen [3] ;
assign \io_master_arlen [7] = \io_master_arlen [3] ;
assign \io_master_arsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign \io_master_awid [0] = \io_master_arburst [1] ;
assign \io_master_awid [1] = \io_master_arburst [1] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;

NOR2_X4 _10800_ ( .A1(\IDU.inst_i [3] ), .A2(\IDU.inst_i [2] ), .ZN(_03721_ ) );
INV_X2 _10801_ ( .A(\IDU.inst_i [4] ), .ZN(_03722_ ) );
AND3_X1 _10802_ ( .A1(_03721_ ), .A2(\IDU.inst_i [5] ), .A3(_03722_ ), .ZN(_03723_ ) );
AND2_X1 _10803_ ( .A1(_03723_ ), .A2(\IDU.inst_i [6] ), .ZN(_03724_ ) );
AND2_X1 _10804_ ( .A1(_03723_ ), .A2(\IDU.ls_valid_o_$_DFFE_PP__Q_D_$_ANDNOT__Y_B_$_NOR__Y_B_$_ANDNOT__Y_A ), .ZN(_03725_ ) );
NOR2_X2 _10805_ ( .A1(_03724_ ), .A2(_03725_ ), .ZN(_03726_ ) );
INV_X1 _10806_ ( .A(_03726_ ), .ZN(_03727_ ) );
AND3_X1 _10807_ ( .A1(_03722_ ), .A2(\IDU.inst_i [6] ), .A3(\IDU.inst_i [5] ), .ZN(_03728_ ) );
INV_X1 _10808_ ( .A(\IDU.inst_i [2] ), .ZN(_03729_ ) );
NOR2_X1 _10809_ ( .A1(_03729_ ), .A2(\IDU.inst_i [3] ), .ZN(_03730_ ) );
AND2_X1 _10810_ ( .A1(_03728_ ), .A2(_03730_ ), .ZN(_03731_ ) );
INV_X1 _10811_ ( .A(\IDU.inst_i [6] ), .ZN(_03732_ ) );
INV_X1 _10812_ ( .A(\IDU.inst_i [5] ), .ZN(_03733_ ) );
AND4_X1 _10813_ ( .A1(_03732_ ), .A2(_03721_ ), .A3(_03733_ ), .A4(_03722_ ), .ZN(_03734_ ) );
AND2_X4 _10814_ ( .A1(\IDU.inst_i [4] ), .A2(\IDU.ls_valid_o_$_DFFE_PP__Q_D_$_ANDNOT__Y_B_$_NOR__Y_B_$_ANDNOT__Y_A ), .ZN(_03735_ ) );
AND3_X1 _10815_ ( .A1(_03735_ ), .A2(_03733_ ), .A3(_03721_ ), .ZN(_03736_ ) );
OR3_X1 _10816_ ( .A1(_03731_ ), .A2(_03734_ ), .A3(_03736_ ), .ZN(_03737_ ) );
AND2_X1 _10817_ ( .A1(\IDU.inst_i [5] ), .A2(\IDU.inst_i [4] ), .ZN(_03738_ ) );
AND2_X1 _10818_ ( .A1(_03738_ ), .A2(_03721_ ), .ZN(_03739_ ) );
AND2_X1 _10819_ ( .A1(_03739_ ), .A2(\IDU.inst_i [6] ), .ZN(_03740_ ) );
NOR3_X4 _10820_ ( .A1(_03727_ ), .A2(_03737_ ), .A3(_03740_ ), .ZN(_03741_ ) );
AND2_X1 _10821_ ( .A1(_03739_ ), .A2(_03732_ ), .ZN(_03742_ ) );
INV_X1 _10822_ ( .A(_03742_ ), .ZN(_03743_ ) );
AND2_X2 _10823_ ( .A1(_03741_ ), .A2(_03743_ ), .ZN(_03744_ ) );
AND2_X1 _10824_ ( .A1(\IDU.inst_i [3] ), .A2(\IDU.inst_i [2] ), .ZN(_03745_ ) );
AND2_X1 _10825_ ( .A1(_03728_ ), .A2(_03745_ ), .ZN(_03746_ ) );
INV_X1 _10826_ ( .A(_03746_ ), .ZN(_03747_ ) );
AND2_X4 _10827_ ( .A1(_03744_ ), .A2(_03747_ ), .ZN(_03748_ ) );
BUF_X2 _10828_ ( .A(_03748_ ), .Z(_03749_ ) );
INV_X1 _10829_ ( .A(\BTB.btag_pre [3] ), .ZN(_03750_ ) );
OR3_X1 _10830_ ( .A1(_03749_ ), .A2(_03750_ ), .A3(\IDU.imm_$_NOR__Y_5_A_$_MUX__Y_B ), .ZN(_03751_ ) );
NOR3_X1 _10831_ ( .A1(_03749_ ), .A2(\IDU.imm_$_NOR__Y_6_A_$_MUX__Y_B ), .A3(prepc_$_ANDNOT__Y_10_B_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_03752_ ) );
NOR2_X4 _10832_ ( .A1(_03737_ ), .A2(_03740_ ), .ZN(_03753_ ) );
AOI21_X1 _10833_ ( .A(\IDU.imm_$_NOR__Y_7_A_$_MUX__Y_B ), .B1(_03753_ ), .B2(_03747_ ), .ZN(_03754_ ) );
BUF_X2 _10834_ ( .A(_03746_ ), .Z(_03755_ ) );
NOR3_X1 _10835_ ( .A1(_03726_ ), .A2(\IDU.imm_$_NOR__Y_7_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03755_ ), .ZN(_03756_ ) );
OAI21_X1 _10836_ ( .A(\BTB.btag_pre [1] ), .B1(_03754_ ), .B2(_03756_ ), .ZN(_03757_ ) );
AOI21_X1 _10837_ ( .A(\IDU.imm_$_NOR__Y_9_A_$_MUX__Y_B ), .B1(_03753_ ), .B2(_03747_ ), .ZN(_03758_ ) );
NOR3_X1 _10838_ ( .A1(_03726_ ), .A2(\IDU.imm_$_NOR__Y_9_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03755_ ), .ZN(_03759_ ) );
OAI21_X1 _10839_ ( .A(\BTB.bindex_pre ), .B1(_03758_ ), .B2(_03759_ ), .ZN(_03760_ ) );
AOI21_X1 _10840_ ( .A(\IDU.imm_$_NOR__Y_10_A_$_MUX__Y_B ), .B1(_03753_ ), .B2(_03747_ ), .ZN(_03761_ ) );
NOR3_X1 _10841_ ( .A1(_03726_ ), .A2(\IDU.imm_$_NOR__Y_10_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03755_ ), .ZN(_03762_ ) );
NOR2_X1 _10842_ ( .A1(_03761_ ), .A2(_03762_ ), .ZN(_03763_ ) );
XNOR2_X1 _10843_ ( .A(_03763_ ), .B(\BTB.prepc_tag_i [1] ), .ZN(_03764_ ) );
INV_X1 _10844_ ( .A(_03725_ ), .ZN(_03765_ ) );
OAI21_X1 _10845_ ( .A(_03765_ ), .B1(_03753_ ), .B2(\IDU.imm_$_NOR__Y_A_$_MUX__Y_B ), .ZN(_03766_ ) );
AOI22_X1 _10846_ ( .A1(_03725_ ), .A2(\IDU.imm_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B1(\IDU.inst_i [6] ), .B2(_03723_ ), .ZN(_03767_ ) );
AND3_X1 _10847_ ( .A1(_03766_ ), .A2(\BTB.prepc_tag_i [0] ), .A3(_03767_ ), .ZN(_03768_ ) );
AND2_X1 _10848_ ( .A1(_03764_ ), .A2(_03768_ ), .ZN(_03769_ ) );
INV_X1 _10849_ ( .A(_03763_ ), .ZN(_03770_ ) );
AOI21_X1 _10850_ ( .A(_03769_ ), .B1(\BTB.prepc_tag_i [1] ), .B2(_03770_ ), .ZN(_03771_ ) );
OR2_X1 _10851_ ( .A1(_03758_ ), .A2(_03759_ ), .ZN(_03772_ ) );
XOR2_X1 _10852_ ( .A(_03772_ ), .B(prepc_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .Z(_03773_ ) );
OAI21_X2 _10853_ ( .A(_03760_ ), .B1(_03771_ ), .B2(_03773_ ), .ZN(_03774_ ) );
AOI21_X1 _10854_ ( .A(\IDU.imm_$_NOR__Y_8_A_$_MUX__Y_B ), .B1(_03753_ ), .B2(_03747_ ), .ZN(_03775_ ) );
NOR3_X1 _10855_ ( .A1(_03726_ ), .A2(\IDU.imm_$_NOR__Y_8_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03755_ ), .ZN(_03776_ ) );
OR2_X1 _10856_ ( .A1(_03775_ ), .A2(_03776_ ), .ZN(_03777_ ) );
XNOR2_X1 _10857_ ( .A(_03777_ ), .B(prepc_$_ANDNOT__Y_12_B_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_03778_ ) );
NAND2_X1 _10858_ ( .A1(_03774_ ), .A2(_03778_ ), .ZN(_03779_ ) );
INV_X1 _10859_ ( .A(prepc_$_ANDNOT__Y_12_B_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_03780_ ) );
OAI21_X1 _10860_ ( .A(_03780_ ), .B1(_03775_ ), .B2(_03776_ ), .ZN(_03781_ ) );
AND2_X2 _10861_ ( .A1(_03779_ ), .A2(_03781_ ), .ZN(_03782_ ) );
NOR3_X1 _10862_ ( .A1(_03754_ ), .A2(\BTB.btag_pre [1] ), .A3(_03756_ ), .ZN(_03783_ ) );
OAI21_X1 _10863_ ( .A(_03757_ ), .B1(_03782_ ), .B2(_03783_ ), .ZN(_03784_ ) );
NOR2_X1 _10864_ ( .A1(_03748_ ), .A2(\IDU.imm_$_NOR__Y_6_A_$_MUX__Y_B ), .ZN(_03785_ ) );
XNOR2_X1 _10865_ ( .A(_03785_ ), .B(prepc_$_ANDNOT__Y_10_B_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_03786_ ) );
AOI21_X2 _10866_ ( .A(_03752_ ), .B1(_03784_ ), .B2(_03786_ ), .ZN(_03787_ ) );
NOR2_X4 _10867_ ( .A1(_03749_ ), .A2(\IDU.imm_$_NOR__Y_5_A_$_MUX__Y_B ), .ZN(_03788_ ) );
XNOR2_X1 _10868_ ( .A(_03788_ ), .B(_03750_ ), .ZN(_03789_ ) );
INV_X1 _10869_ ( .A(_03789_ ), .ZN(_03790_ ) );
OAI21_X1 _10870_ ( .A(_03751_ ), .B1(_03787_ ), .B2(_03790_ ), .ZN(_03791_ ) );
NOR2_X1 _10871_ ( .A1(_03748_ ), .A2(\IDU.imm_$_NOR__Y_4_A_$_MUX__Y_B ), .ZN(_03792_ ) );
XNOR2_X1 _10872_ ( .A(_03792_ ), .B(prepc_$_ANDNOT__Y_8_B_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_03793_ ) );
INV_X1 _10873_ ( .A(_03793_ ), .ZN(_03794_ ) );
XNOR2_X1 _10874_ ( .A(_03791_ ), .B(_03794_ ), .ZN(_03795_ ) );
INV_X1 _10875_ ( .A(_03724_ ), .ZN(_03796_ ) );
NOR2_X1 _10876_ ( .A1(_03796_ ), .A2(\IDU.prevalid_$_NAND__B_A_$_ANDNOT__Y_B ), .ZN(_03797_ ) );
INV_X1 _10877_ ( .A(fanout_net_11 ), .ZN(_03798_ ) );
AND3_X1 _10878_ ( .A1(_03797_ ), .A2(_03798_ ), .A3(\IDU.prevalid ), .ZN(_03799_ ) );
OR2_X2 _10879_ ( .A1(_03797_ ), .A2(_03755_ ), .ZN(_03800_ ) );
BUF_X4 _10880_ ( .A(_03800_ ), .Z(_03801_ ) );
NAND4_X1 _10881_ ( .A1(_03795_ ), .A2(prepc_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .A3(_03799_ ), .A4(_03801_ ), .ZN(_03802_ ) );
NAND2_X1 _10882_ ( .A1(_03799_ ), .A2(prepc_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_03803_ ) );
BUF_X4 _10883_ ( .A(_03803_ ), .Z(_03804_ ) );
BUF_X4 _10884_ ( .A(_03798_ ), .Z(_03805_ ) );
BUF_X2 _10885_ ( .A(_03805_ ), .Z(_03806_ ) );
NAND3_X1 _10886_ ( .A1(_03804_ ), .A2(\BTB.bsnpc_reg[0][7] ), .A3(_03806_ ), .ZN(_03807_ ) );
NAND2_X1 _10887_ ( .A1(_03802_ ), .A2(_03807_ ), .ZN(_00000_ ) );
BUF_X8 _10888_ ( .A(_03805_ ), .Z(_03808_ ) );
BUF_X4 _10889_ ( .A(_03808_ ), .Z(_03809_ ) );
NAND3_X1 _10890_ ( .A1(_03804_ ), .A2(\BTB.bsnpc_reg[0][6] ), .A3(_03809_ ), .ZN(_03810_ ) );
XNOR2_X1 _10891_ ( .A(_03787_ ), .B(_03789_ ), .ZN(_03811_ ) );
NAND2_X1 _10892_ ( .A1(_03811_ ), .A2(_03801_ ), .ZN(_03812_ ) );
BUF_X4 _10893_ ( .A(_03803_ ), .Z(_03813_ ) );
BUF_X4 _10894_ ( .A(_03813_ ), .Z(_03814_ ) );
OAI21_X1 _10895_ ( .A(_03810_ ), .B1(_03812_ ), .B2(_03814_ ), .ZN(_00001_ ) );
NAND3_X1 _10896_ ( .A1(_03804_ ), .A2(\BTB.bsnpc_reg[0][5] ), .A3(_03809_ ), .ZN(_03815_ ) );
XOR2_X1 _10897_ ( .A(_03784_ ), .B(_03786_ ), .Z(_03816_ ) );
NAND2_X1 _10898_ ( .A1(_03816_ ), .A2(_03801_ ), .ZN(_03817_ ) );
OAI21_X1 _10899_ ( .A(_03815_ ), .B1(_03817_ ), .B2(_03814_ ), .ZN(_00002_ ) );
NAND3_X1 _10900_ ( .A1(_03804_ ), .A2(\BTB.bsnpc_reg[0][4] ), .A3(_03809_ ), .ZN(_03818_ ) );
NOR2_X1 _10901_ ( .A1(_03754_ ), .A2(_03756_ ), .ZN(_03819_ ) );
XNOR2_X1 _10902_ ( .A(_03819_ ), .B(\BTB.btag_pre [1] ), .ZN(_03820_ ) );
XNOR2_X1 _10903_ ( .A(_03782_ ), .B(_03820_ ), .ZN(_03821_ ) );
NAND2_X1 _10904_ ( .A1(_03821_ ), .A2(_03801_ ), .ZN(_03822_ ) );
OAI21_X1 _10905_ ( .A(_03818_ ), .B1(_03822_ ), .B2(_03814_ ), .ZN(_00003_ ) );
NAND3_X1 _10906_ ( .A1(_03804_ ), .A2(\BTB.bsnpc_reg[0][3] ), .A3(_03809_ ), .ZN(_03823_ ) );
XOR2_X1 _10907_ ( .A(_03774_ ), .B(_03778_ ), .Z(_03824_ ) );
NAND2_X1 _10908_ ( .A1(_03824_ ), .A2(_03801_ ), .ZN(_03825_ ) );
OAI21_X1 _10909_ ( .A(_03823_ ), .B1(_03825_ ), .B2(_03814_ ), .ZN(_00004_ ) );
NAND3_X1 _10910_ ( .A1(_03804_ ), .A2(\BTB.bsnpc_reg[0][2] ), .A3(_03809_ ), .ZN(_03826_ ) );
XOR2_X1 _10911_ ( .A(_03771_ ), .B(_03773_ ), .Z(_03827_ ) );
NAND2_X1 _10912_ ( .A1(_03827_ ), .A2(_03801_ ), .ZN(_03828_ ) );
OAI21_X1 _10913_ ( .A(_03826_ ), .B1(_03828_ ), .B2(_03814_ ), .ZN(_00005_ ) );
OR2_X1 _10914_ ( .A1(_03764_ ), .A2(_03768_ ), .ZN(_03829_ ) );
NAND2_X1 _10915_ ( .A1(_03829_ ), .A2(_03800_ ), .ZN(_03830_ ) );
BUF_X4 _10916_ ( .A(_03803_ ), .Z(_03831_ ) );
INV_X1 _10917_ ( .A(\BTB.bsnpc_reg[0][1] ), .ZN(_03832_ ) );
BUF_X4 _10918_ ( .A(_03805_ ), .Z(_03833_ ) );
NAND2_X1 _10919_ ( .A1(_03813_ ), .A2(_03833_ ), .ZN(_03834_ ) );
OAI22_X1 _10920_ ( .A1(_03830_ ), .A2(_03831_ ), .B1(_03832_ ), .B2(_03834_ ), .ZN(_00006_ ) );
AND2_X1 _10921_ ( .A1(_03766_ ), .A2(_03767_ ), .ZN(_03835_ ) );
OR2_X1 _10922_ ( .A1(_03835_ ), .A2(\BTB.prepc_tag_i [0] ), .ZN(_03836_ ) );
NAND2_X1 _10923_ ( .A1(_03836_ ), .A2(_03800_ ), .ZN(_03837_ ) );
INV_X1 _10924_ ( .A(\BTB.bsnpc_reg[0][0] ), .ZN(_03838_ ) );
OAI22_X1 _10925_ ( .A1(_03837_ ), .A2(_03831_ ), .B1(_03838_ ), .B2(_03834_ ), .ZN(_00007_ ) );
NAND2_X2 _10926_ ( .A1(_03799_ ), .A2(\BTB.bindex_pre ), .ZN(_03839_ ) );
BUF_X4 _10927_ ( .A(_03839_ ), .Z(_03840_ ) );
NAND3_X1 _10928_ ( .A1(_03840_ ), .A2(\BTB.bsnpc_reg[1][7] ), .A3(_03809_ ), .ZN(_03841_ ) );
NAND2_X1 _10929_ ( .A1(_03795_ ), .A2(_03801_ ), .ZN(_03842_ ) );
BUF_X4 _10930_ ( .A(_03839_ ), .Z(_03843_ ) );
OAI21_X1 _10931_ ( .A(_03841_ ), .B1(_03842_ ), .B2(_03843_ ), .ZN(_00008_ ) );
BUF_X4 _10932_ ( .A(_03805_ ), .Z(_03844_ ) );
BUF_X4 _10933_ ( .A(_03844_ ), .Z(_03845_ ) );
NAND3_X1 _10934_ ( .A1(_03840_ ), .A2(\BTB.bsnpc_reg[1][6] ), .A3(_03845_ ), .ZN(_03846_ ) );
OAI21_X1 _10935_ ( .A(_03846_ ), .B1(_03812_ ), .B2(_03843_ ), .ZN(_00009_ ) );
NAND3_X1 _10936_ ( .A1(_03840_ ), .A2(\BTB.bsnpc_reg[1][5] ), .A3(_03845_ ), .ZN(_03847_ ) );
OAI21_X1 _10937_ ( .A(_03847_ ), .B1(_03817_ ), .B2(_03843_ ), .ZN(_00010_ ) );
NAND3_X1 _10938_ ( .A1(_03840_ ), .A2(\BTB.bsnpc_reg[1][4] ), .A3(_03845_ ), .ZN(_03848_ ) );
OAI21_X1 _10939_ ( .A(_03848_ ), .B1(_03822_ ), .B2(_03843_ ), .ZN(_00011_ ) );
NAND3_X1 _10940_ ( .A1(_03840_ ), .A2(\BTB.bsnpc_reg[1][3] ), .A3(_03845_ ), .ZN(_03849_ ) );
OAI21_X1 _10941_ ( .A(_03849_ ), .B1(_03825_ ), .B2(_03843_ ), .ZN(_00012_ ) );
NAND3_X1 _10942_ ( .A1(_03840_ ), .A2(\BTB.bsnpc_reg[1][2] ), .A3(_03845_ ), .ZN(_03850_ ) );
OAI21_X1 _10943_ ( .A(_03850_ ), .B1(_03828_ ), .B2(_03843_ ), .ZN(_00013_ ) );
BUF_X4 _10944_ ( .A(_03839_ ), .Z(_03851_ ) );
INV_X1 _10945_ ( .A(\BTB.bsnpc_reg[1][1] ), .ZN(_03852_ ) );
NAND2_X1 _10946_ ( .A1(_03839_ ), .A2(_03833_ ), .ZN(_03853_ ) );
OAI22_X1 _10947_ ( .A1(_03830_ ), .A2(_03851_ ), .B1(_03852_ ), .B2(_03853_ ), .ZN(_00014_ ) );
INV_X1 _10948_ ( .A(\BTB.bsnpc_reg[1][0] ), .ZN(_03854_ ) );
OAI22_X1 _10949_ ( .A1(_03837_ ), .A2(_03840_ ), .B1(_03854_ ), .B2(_03853_ ), .ZN(_00015_ ) );
NAND3_X1 _10950_ ( .A1(_03804_ ), .A2(\BTB.btag_reg[0][12] ), .A3(_03845_ ), .ZN(_03855_ ) );
INV_X1 _10951_ ( .A(\BTB.btag_pre [12] ), .ZN(_03856_ ) );
OAI21_X1 _10952_ ( .A(_03855_ ), .B1(_03856_ ), .B2(_03814_ ), .ZN(_00016_ ) );
NAND3_X1 _10953_ ( .A1(_03804_ ), .A2(\BTB.btag_reg[0][11] ), .A3(_03845_ ), .ZN(_03857_ ) );
INV_X1 _10954_ ( .A(\BTB.btag_pre [11] ), .ZN(_03858_ ) );
OAI21_X1 _10955_ ( .A(_03857_ ), .B1(_03858_ ), .B2(_03814_ ), .ZN(_00017_ ) );
NAND3_X1 _10956_ ( .A1(_03804_ ), .A2(\BTB.btag_reg[0][2] ), .A3(_03845_ ), .ZN(_03859_ ) );
INV_X1 _10957_ ( .A(\BTB.btag_pre [2] ), .ZN(_03860_ ) );
OAI21_X1 _10958_ ( .A(_03859_ ), .B1(_03860_ ), .B2(_03814_ ), .ZN(_00018_ ) );
NAND3_X1 _10959_ ( .A1(_03804_ ), .A2(\BTB.btag_reg[0][1] ), .A3(_03845_ ), .ZN(_03861_ ) );
INV_X1 _10960_ ( .A(\BTB.btag_pre [1] ), .ZN(_03862_ ) );
OAI21_X1 _10961_ ( .A(_03861_ ), .B1(_03862_ ), .B2(_03814_ ), .ZN(_00019_ ) );
NAND3_X1 _10962_ ( .A1(_03813_ ), .A2(\BTB.btag_reg[0][0] ), .A3(_03845_ ), .ZN(_03863_ ) );
INV_X1 _10963_ ( .A(\BTB.btag_pre [0] ), .ZN(_03864_ ) );
OAI21_X1 _10964_ ( .A(_03863_ ), .B1(_03864_ ), .B2(_03814_ ), .ZN(_00020_ ) );
BUF_X4 _10965_ ( .A(_03808_ ), .Z(_03865_ ) );
NAND3_X1 _10966_ ( .A1(_03813_ ), .A2(\BTB.btag_reg[0][10] ), .A3(_03865_ ), .ZN(_03866_ ) );
INV_X1 _10967_ ( .A(\BTB.btag_pre [10] ), .ZN(_03867_ ) );
OAI21_X1 _10968_ ( .A(_03866_ ), .B1(_03867_ ), .B2(_03831_ ), .ZN(_00021_ ) );
NAND3_X1 _10969_ ( .A1(_03813_ ), .A2(\BTB.btag_reg[0][9] ), .A3(_03865_ ), .ZN(_03868_ ) );
INV_X1 _10970_ ( .A(\BTB.btag_pre [9] ), .ZN(_03869_ ) );
OAI21_X1 _10971_ ( .A(_03868_ ), .B1(_03869_ ), .B2(_03831_ ), .ZN(_00022_ ) );
NAND3_X1 _10972_ ( .A1(_03813_ ), .A2(\BTB.btag_reg[0][8] ), .A3(_03865_ ), .ZN(_03870_ ) );
INV_X1 _10973_ ( .A(\BTB.btag_pre [8] ), .ZN(_03871_ ) );
OAI21_X1 _10974_ ( .A(_03870_ ), .B1(_03871_ ), .B2(_03831_ ), .ZN(_00023_ ) );
NAND3_X1 _10975_ ( .A1(_03813_ ), .A2(\BTB.btag_reg[0][7] ), .A3(_03865_ ), .ZN(_03872_ ) );
INV_X1 _10976_ ( .A(\BTB.btag_pre [7] ), .ZN(_03873_ ) );
OAI21_X1 _10977_ ( .A(_03872_ ), .B1(_03873_ ), .B2(_03831_ ), .ZN(_00024_ ) );
NAND3_X1 _10978_ ( .A1(_03813_ ), .A2(\BTB.btag_reg[0][6] ), .A3(_03865_ ), .ZN(_03874_ ) );
INV_X1 _10979_ ( .A(\BTB.btag_pre [6] ), .ZN(_03875_ ) );
OAI21_X1 _10980_ ( .A(_03874_ ), .B1(_03875_ ), .B2(_03831_ ), .ZN(_00025_ ) );
NAND3_X1 _10981_ ( .A1(_03813_ ), .A2(\BTB.btag_reg[0][5] ), .A3(_03865_ ), .ZN(_03876_ ) );
INV_X1 _10982_ ( .A(\BTB.btag_pre [5] ), .ZN(_03877_ ) );
OAI21_X1 _10983_ ( .A(_03876_ ), .B1(_03877_ ), .B2(_03831_ ), .ZN(_00026_ ) );
NAND3_X1 _10984_ ( .A1(_03831_ ), .A2(\BTB.btag_reg[0][4] ), .A3(_03806_ ), .ZN(_03878_ ) );
NAND3_X1 _10985_ ( .A1(_03799_ ), .A2(\BTB.btag_pre [4] ), .A3(prepc_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_03879_ ) );
NAND2_X1 _10986_ ( .A1(_03878_ ), .A2(_03879_ ), .ZN(_00027_ ) );
NAND3_X1 _10987_ ( .A1(_03813_ ), .A2(\BTB.btag_reg[0][3] ), .A3(_03865_ ), .ZN(_03880_ ) );
OAI21_X1 _10988_ ( .A(_03880_ ), .B1(_03750_ ), .B2(_03831_ ), .ZN(_00028_ ) );
NAND3_X1 _10989_ ( .A1(_03840_ ), .A2(\BTB.btag_reg[1][12] ), .A3(_03865_ ), .ZN(_03881_ ) );
OAI21_X1 _10990_ ( .A(_03881_ ), .B1(_03856_ ), .B2(_03843_ ), .ZN(_00029_ ) );
NAND3_X1 _10991_ ( .A1(_03840_ ), .A2(\BTB.btag_reg[1][11] ), .A3(_03865_ ), .ZN(_03882_ ) );
OAI21_X1 _10992_ ( .A(_03882_ ), .B1(_03858_ ), .B2(_03843_ ), .ZN(_00030_ ) );
NAND3_X1 _10993_ ( .A1(_03840_ ), .A2(\BTB.btag_reg[1][2] ), .A3(_03865_ ), .ZN(_03883_ ) );
OAI21_X1 _10994_ ( .A(_03883_ ), .B1(_03860_ ), .B2(_03843_ ), .ZN(_00031_ ) );
BUF_X4 _10995_ ( .A(_03839_ ), .Z(_03884_ ) );
BUF_X4 _10996_ ( .A(_03808_ ), .Z(_03885_ ) );
NAND3_X1 _10997_ ( .A1(_03884_ ), .A2(\BTB.btag_reg[1][1] ), .A3(_03885_ ), .ZN(_03886_ ) );
OAI21_X1 _10998_ ( .A(_03886_ ), .B1(_03862_ ), .B2(_03843_ ), .ZN(_00032_ ) );
NAND3_X1 _10999_ ( .A1(_03884_ ), .A2(\BTB.btag_reg[1][0] ), .A3(_03885_ ), .ZN(_03887_ ) );
OAI21_X1 _11000_ ( .A(_03887_ ), .B1(_03864_ ), .B2(_03851_ ), .ZN(_00033_ ) );
NAND3_X1 _11001_ ( .A1(_03884_ ), .A2(\BTB.btag_reg[1][10] ), .A3(_03885_ ), .ZN(_03888_ ) );
OAI21_X1 _11002_ ( .A(_03888_ ), .B1(_03867_ ), .B2(_03851_ ), .ZN(_00034_ ) );
NAND3_X1 _11003_ ( .A1(_03884_ ), .A2(\BTB.btag_reg[1][9] ), .A3(_03885_ ), .ZN(_03889_ ) );
OAI21_X1 _11004_ ( .A(_03889_ ), .B1(_03869_ ), .B2(_03851_ ), .ZN(_00035_ ) );
NAND3_X1 _11005_ ( .A1(_03884_ ), .A2(\BTB.btag_reg[1][8] ), .A3(_03885_ ), .ZN(_03890_ ) );
OAI21_X1 _11006_ ( .A(_03890_ ), .B1(_03871_ ), .B2(_03851_ ), .ZN(_00036_ ) );
NAND3_X1 _11007_ ( .A1(_03884_ ), .A2(\BTB.btag_reg[1][7] ), .A3(_03885_ ), .ZN(_03891_ ) );
OAI21_X1 _11008_ ( .A(_03891_ ), .B1(_03873_ ), .B2(_03851_ ), .ZN(_00037_ ) );
NAND3_X1 _11009_ ( .A1(_03884_ ), .A2(\BTB.btag_reg[1][6] ), .A3(_03885_ ), .ZN(_03892_ ) );
OAI21_X1 _11010_ ( .A(_03892_ ), .B1(_03875_ ), .B2(_03851_ ), .ZN(_00038_ ) );
NAND3_X1 _11011_ ( .A1(_03884_ ), .A2(\BTB.btag_reg[1][5] ), .A3(_03885_ ), .ZN(_03893_ ) );
OAI21_X1 _11012_ ( .A(_03893_ ), .B1(_03877_ ), .B2(_03851_ ), .ZN(_00039_ ) );
NAND3_X1 _11013_ ( .A1(_03884_ ), .A2(\BTB.btag_reg[1][4] ), .A3(_03885_ ), .ZN(_03894_ ) );
INV_X1 _11014_ ( .A(\BTB.btag_pre [4] ), .ZN(_03895_ ) );
OAI21_X1 _11015_ ( .A(_03894_ ), .B1(_03895_ ), .B2(_03851_ ), .ZN(_00040_ ) );
NAND3_X1 _11016_ ( .A1(_03884_ ), .A2(\BTB.btag_reg[1][3] ), .A3(_03885_ ), .ZN(_03896_ ) );
OAI21_X1 _11017_ ( .A(_03896_ ), .B1(_03750_ ), .B2(_03851_ ), .ZN(_00041_ ) );
NAND3_X1 _11018_ ( .A1(_03723_ ), .A2(\IDU.prevalid_$_NAND__B_A_$_ANDNOT__Y_B ), .A3(\IDU.ls_valid_o_$_DFFE_PP__Q_D_$_ANDNOT__Y_B_$_NOR__Y_B_$_ANDNOT__Y_A ), .ZN(_03897_ ) );
AOI21_X1 _11019_ ( .A(\IDU.prevalid_$_NAND__B_A_$_ANDNOT__Y_B ), .B1(_03753_ ), .B2(_03743_ ), .ZN(_03898_ ) );
OAI21_X1 _11020_ ( .A(_03897_ ), .B1(_03898_ ), .B2(_03725_ ), .ZN(_03899_ ) );
MUX2_X1 _11021_ ( .A(\IDU.imm_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_03899_ ), .S(_03796_ ), .Z(_03900_ ) );
OR2_X1 _11022_ ( .A1(_03747_ ), .A2(\IDU.imm_$_NOR__Y_A_$_MUX__Y_B ), .ZN(_03901_ ) );
AOI21_X1 _11023_ ( .A(_03871_ ), .B1(_03900_ ), .B2(_03901_ ), .ZN(_03902_ ) );
INV_X1 _11024_ ( .A(_03902_ ), .ZN(_03903_ ) );
NOR3_X1 _11025_ ( .A1(_03749_ ), .A2(\IDU.imm_$_NOR__Y_2_A_$_MUX__Y_B ), .A3(prepc_$_ANDNOT__Y_6_B_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_03904_ ) );
INV_X1 _11026_ ( .A(_03904_ ), .ZN(_03905_ ) );
NOR2_X1 _11027_ ( .A1(_03749_ ), .A2(\IDU.imm_$_NOR__Y_3_A_$_MUX__Y_B ), .ZN(_03906_ ) );
XNOR2_X1 _11028_ ( .A(_03906_ ), .B(_03877_ ), .ZN(_03907_ ) );
NOR3_X1 _11029_ ( .A1(_03787_ ), .A2(_03790_ ), .A3(_03794_ ), .ZN(_03908_ ) );
NAND3_X1 _11030_ ( .A1(_03793_ ), .A2(\BTB.btag_pre [3] ), .A3(_03788_ ), .ZN(_03909_ ) );
INV_X1 _11031_ ( .A(_03792_ ), .ZN(_03910_ ) );
OAI21_X1 _11032_ ( .A(_03909_ ), .B1(prepc_$_ANDNOT__Y_8_B_$_XOR__Y_B_$_XOR__Y_B ), .B2(_03910_ ), .ZN(_03911_ ) );
OAI21_X1 _11033_ ( .A(_03907_ ), .B1(_03908_ ), .B2(_03911_ ), .ZN(_03912_ ) );
OR3_X1 _11034_ ( .A1(_03749_ ), .A2(_03877_ ), .A3(\IDU.imm_$_NOR__Y_3_A_$_MUX__Y_B ), .ZN(_03913_ ) );
AND2_X1 _11035_ ( .A1(_03912_ ), .A2(_03913_ ), .ZN(_03914_ ) );
NOR2_X1 _11036_ ( .A1(_03749_ ), .A2(\IDU.imm_$_NOR__Y_2_A_$_MUX__Y_B ), .ZN(_03915_ ) );
INV_X1 _11037_ ( .A(_03915_ ), .ZN(_03916_ ) );
AND2_X1 _11038_ ( .A1(_03916_ ), .A2(prepc_$_ANDNOT__Y_6_B_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_03917_ ) );
OAI21_X2 _11039_ ( .A(_03905_ ), .B1(_03914_ ), .B2(_03917_ ), .ZN(_03918_ ) );
NOR2_X1 _11040_ ( .A1(_03749_ ), .A2(\IDU.imm_$_NOR__Y_1_A_$_MUX__Y_B ), .ZN(_03919_ ) );
XNOR2_X1 _11041_ ( .A(_03919_ ), .B(_03873_ ), .ZN(_03920_ ) );
NAND2_X1 _11042_ ( .A1(_03918_ ), .A2(_03920_ ), .ZN(_03921_ ) );
OR3_X1 _11043_ ( .A1(_03749_ ), .A2(_03873_ ), .A3(\IDU.imm_$_NOR__Y_1_A_$_MUX__Y_B ), .ZN(_03922_ ) );
AND2_X1 _11044_ ( .A1(_03921_ ), .A2(_03922_ ), .ZN(_03923_ ) );
AND3_X1 _11045_ ( .A1(_03900_ ), .A2(_03871_ ), .A3(_03901_ ), .ZN(_03924_ ) );
OAI21_X2 _11046_ ( .A(_03903_ ), .B1(_03923_ ), .B2(_03924_ ), .ZN(_03925_ ) );
INV_X1 _11047_ ( .A(\IDU.funct7 [6] ), .ZN(_03926_ ) );
NOR2_X1 _11048_ ( .A1(_03741_ ), .A2(_03926_ ), .ZN(_03927_ ) );
AND2_X1 _11049_ ( .A1(_03730_ ), .A2(_03735_ ), .ZN(_03928_ ) );
NOR2_X1 _11050_ ( .A1(_03755_ ), .A2(_03928_ ), .ZN(_03929_ ) );
INV_X1 _11051_ ( .A(_03929_ ), .ZN(_03930_ ) );
AND2_X1 _11052_ ( .A1(_03930_ ), .A2(\IDU.funct3 [0] ), .ZN(_03931_ ) );
NOR2_X1 _11053_ ( .A1(_03927_ ), .A2(_03931_ ), .ZN(_03932_ ) );
XNOR2_X1 _11054_ ( .A(_03932_ ), .B(\BTB.btag_pre [9] ), .ZN(_03933_ ) );
INV_X1 _11055_ ( .A(_03927_ ), .ZN(_03934_ ) );
OAI21_X1 _11056_ ( .A(\IDU.funct3 [1] ), .B1(_03755_ ), .B2(_03928_ ), .ZN(_03935_ ) );
AND3_X1 _11057_ ( .A1(_03934_ ), .A2(_03867_ ), .A3(_03935_ ), .ZN(_03936_ ) );
AOI21_X1 _11058_ ( .A(_03867_ ), .B1(_03934_ ), .B2(_03935_ ), .ZN(_03937_ ) );
NOR2_X1 _11059_ ( .A1(_03936_ ), .A2(_03937_ ), .ZN(_03938_ ) );
AND3_X1 _11060_ ( .A1(_03925_ ), .A2(_03933_ ), .A3(_03938_ ), .ZN(_03939_ ) );
NOR4_X1 _11061_ ( .A1(_03936_ ), .A2(_03937_ ), .A3(_03869_ ), .A4(_03932_ ), .ZN(_03940_ ) );
OR3_X4 _11062_ ( .A1(_03939_ ), .A2(_03937_ ), .A3(_03940_ ), .ZN(_03941_ ) );
OAI21_X1 _11063_ ( .A(\IDU.funct3 [2] ), .B1(_03755_ ), .B2(_03928_ ), .ZN(_03942_ ) );
AND2_X1 _11064_ ( .A1(_03934_ ), .A2(_03942_ ), .ZN(_03943_ ) );
XNOR2_X1 _11065_ ( .A(_03943_ ), .B(\BTB.btag_pre [11] ), .ZN(_03944_ ) );
AND2_X1 _11066_ ( .A1(_03941_ ), .A2(_03944_ ), .ZN(_03945_ ) );
INV_X1 _11067_ ( .A(_03943_ ), .ZN(_03946_ ) );
AOI21_X1 _11068_ ( .A(_03945_ ), .B1(\BTB.btag_pre [11] ), .B2(_03946_ ), .ZN(_03947_ ) );
INV_X1 _11069_ ( .A(_03947_ ), .ZN(_03948_ ) );
INV_X1 _11070_ ( .A(\IDU.immJ [15] ), .ZN(_03949_ ) );
NOR2_X1 _11071_ ( .A1(_03929_ ), .A2(_03949_ ), .ZN(_03950_ ) );
OR2_X1 _11072_ ( .A1(_03927_ ), .A2(_03950_ ), .ZN(_03951_ ) );
XNOR2_X1 _11073_ ( .A(_03951_ ), .B(_03856_ ), .ZN(_03952_ ) );
AND2_X1 _11074_ ( .A1(_03948_ ), .A2(_03952_ ), .ZN(_03953_ ) );
OAI21_X1 _11075_ ( .A(_03800_ ), .B1(_03948_ ), .B2(_03952_ ), .ZN(_03954_ ) );
OR2_X2 _11076_ ( .A1(_03953_ ), .A2(_03954_ ), .ZN(_03955_ ) );
AND3_X1 _11077_ ( .A1(_03755_ ), .A2(_03798_ ), .A3(\IDU.prevalid ), .ZN(_03956_ ) );
NAND2_X1 _11078_ ( .A1(_03956_ ), .A2(prepc_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_03957_ ) );
BUF_X4 _11079_ ( .A(_03957_ ), .Z(_03958_ ) );
BUF_X4 _11080_ ( .A(_03958_ ), .Z(_03959_ ) );
INV_X1 _11081_ ( .A(\BTB.jsnpc_reg[0][15] ), .ZN(_03960_ ) );
NAND2_X2 _11082_ ( .A1(_03957_ ), .A2(_03844_ ), .ZN(_03961_ ) );
OAI22_X1 _11083_ ( .A1(_03955_ ), .A2(_03959_ ), .B1(_03960_ ), .B2(_03961_ ), .ZN(_00042_ ) );
INV_X1 _11084_ ( .A(_03797_ ), .ZN(_03962_ ) );
AOI22_X1 _11085_ ( .A1(_03941_ ), .A2(_03944_ ), .B1(_03962_ ), .B2(_03747_ ), .ZN(_03963_ ) );
OAI21_X1 _11086_ ( .A(_03963_ ), .B1(_03941_ ), .B2(_03944_ ), .ZN(_03964_ ) );
BUF_X4 _11087_ ( .A(_03957_ ), .Z(_03965_ ) );
INV_X1 _11088_ ( .A(\BTB.jsnpc_reg[0][14] ), .ZN(_03966_ ) );
OAI22_X1 _11089_ ( .A1(_03964_ ), .A2(_03965_ ), .B1(_03966_ ), .B2(_03961_ ), .ZN(_00043_ ) );
BUF_X4 _11090_ ( .A(_03808_ ), .Z(_03967_ ) );
NAND3_X1 _11091_ ( .A1(_03965_ ), .A2(\BTB.jsnpc_reg[0][5] ), .A3(_03967_ ), .ZN(_03968_ ) );
BUF_X4 _11092_ ( .A(_03958_ ), .Z(_03969_ ) );
OAI21_X1 _11093_ ( .A(_03968_ ), .B1(_03817_ ), .B2(_03969_ ), .ZN(_00044_ ) );
BUF_X4 _11094_ ( .A(_03957_ ), .Z(_03970_ ) );
NAND3_X1 _11095_ ( .A1(_03970_ ), .A2(\BTB.jsnpc_reg[0][4] ), .A3(_03967_ ), .ZN(_03971_ ) );
OAI21_X1 _11096_ ( .A(_03971_ ), .B1(_03822_ ), .B2(_03969_ ), .ZN(_00045_ ) );
NAND3_X1 _11097_ ( .A1(_03970_ ), .A2(\BTB.jsnpc_reg[0][3] ), .A3(_03967_ ), .ZN(_03972_ ) );
OAI21_X1 _11098_ ( .A(_03972_ ), .B1(_03825_ ), .B2(_03969_ ), .ZN(_00046_ ) );
NAND3_X1 _11099_ ( .A1(_03970_ ), .A2(\BTB.jsnpc_reg[0][2] ), .A3(_03967_ ), .ZN(_03973_ ) );
OAI21_X1 _11100_ ( .A(_03973_ ), .B1(_03828_ ), .B2(_03969_ ), .ZN(_00047_ ) );
INV_X1 _11101_ ( .A(\BTB.jsnpc_reg[0][1] ), .ZN(_03974_ ) );
OAI22_X1 _11102_ ( .A1(_03830_ ), .A2(_03965_ ), .B1(_03974_ ), .B2(_03961_ ), .ZN(_00048_ ) );
INV_X1 _11103_ ( .A(\BTB.jsnpc_reg[0][0] ), .ZN(_03975_ ) );
OAI22_X1 _11104_ ( .A1(_03837_ ), .A2(_03965_ ), .B1(_03975_ ), .B2(_03961_ ), .ZN(_00049_ ) );
AND2_X1 _11105_ ( .A1(_03925_ ), .A2(_03933_ ), .ZN(_03976_ ) );
NOR2_X1 _11106_ ( .A1(_03932_ ), .A2(_03869_ ), .ZN(_03977_ ) );
OR3_X1 _11107_ ( .A1(_03976_ ), .A2(_03977_ ), .A3(_03938_ ), .ZN(_03978_ ) );
OAI21_X1 _11108_ ( .A(_03938_ ), .B1(_03976_ ), .B2(_03977_ ), .ZN(_03979_ ) );
NAND3_X1 _11109_ ( .A1(_03978_ ), .A2(_03801_ ), .A3(_03979_ ), .ZN(_03980_ ) );
INV_X1 _11110_ ( .A(\BTB.jsnpc_reg[0][13] ), .ZN(_03981_ ) );
OAI22_X1 _11111_ ( .A1(_03980_ ), .A2(_03965_ ), .B1(_03981_ ), .B2(_03961_ ), .ZN(_00050_ ) );
AOI22_X1 _11112_ ( .A1(_03925_ ), .A2(_03933_ ), .B1(_03962_ ), .B2(_03747_ ), .ZN(_03982_ ) );
OAI21_X1 _11113_ ( .A(_03982_ ), .B1(_03925_ ), .B2(_03933_ ), .ZN(_03983_ ) );
INV_X1 _11114_ ( .A(\BTB.jsnpc_reg[0][12] ), .ZN(_03984_ ) );
OAI22_X1 _11115_ ( .A1(_03983_ ), .A2(_03965_ ), .B1(_03984_ ), .B2(_03961_ ), .ZN(_00051_ ) );
OR3_X1 _11116_ ( .A1(_03923_ ), .A2(_03902_ ), .A3(_03924_ ), .ZN(_03985_ ) );
OAI21_X1 _11117_ ( .A(_03923_ ), .B1(_03902_ ), .B2(_03924_ ), .ZN(_03986_ ) );
NAND3_X1 _11118_ ( .A1(_03985_ ), .A2(_03801_ ), .A3(_03986_ ), .ZN(_03987_ ) );
INV_X1 _11119_ ( .A(\BTB.jsnpc_reg[0][11] ), .ZN(_03988_ ) );
OAI22_X1 _11120_ ( .A1(_03987_ ), .A2(_03965_ ), .B1(_03988_ ), .B2(_03961_ ), .ZN(_00052_ ) );
AOI22_X1 _11121_ ( .A1(_03918_ ), .A2(_03920_ ), .B1(_03962_ ), .B2(_03747_ ), .ZN(_03989_ ) );
OAI21_X1 _11122_ ( .A(_03989_ ), .B1(_03920_ ), .B2(_03918_ ), .ZN(_03990_ ) );
INV_X1 _11123_ ( .A(\BTB.jsnpc_reg[0][10] ), .ZN(_03991_ ) );
OAI22_X1 _11124_ ( .A1(_03990_ ), .A2(_03965_ ), .B1(_03991_ ), .B2(_03961_ ), .ZN(_00053_ ) );
OR3_X1 _11125_ ( .A1(_03914_ ), .A2(_03904_ ), .A3(_03917_ ), .ZN(_03992_ ) );
OAI21_X1 _11126_ ( .A(_03914_ ), .B1(_03904_ ), .B2(_03917_ ), .ZN(_03993_ ) );
NAND3_X1 _11127_ ( .A1(_03992_ ), .A2(_03801_ ), .A3(_03993_ ), .ZN(_03994_ ) );
INV_X1 _11128_ ( .A(\BTB.jsnpc_reg[0][9] ), .ZN(_03995_ ) );
OAI22_X1 _11129_ ( .A1(_03994_ ), .A2(_03965_ ), .B1(_03995_ ), .B2(_03961_ ), .ZN(_00054_ ) );
AND2_X1 _11130_ ( .A1(_03912_ ), .A2(_03800_ ), .ZN(_03996_ ) );
OR2_X1 _11131_ ( .A1(_03908_ ), .A2(_03911_ ), .ZN(_03997_ ) );
OAI21_X1 _11132_ ( .A(_03996_ ), .B1(_03997_ ), .B2(_03907_ ), .ZN(_03998_ ) );
INV_X1 _11133_ ( .A(\BTB.jsnpc_reg[0][8] ), .ZN(_03999_ ) );
OAI22_X1 _11134_ ( .A1(_03998_ ), .A2(_03965_ ), .B1(_03999_ ), .B2(_03961_ ), .ZN(_00055_ ) );
NAND3_X1 _11135_ ( .A1(_03970_ ), .A2(\BTB.jsnpc_reg[0][7] ), .A3(_03967_ ), .ZN(_04000_ ) );
OAI21_X1 _11136_ ( .A(_04000_ ), .B1(_03842_ ), .B2(_03969_ ), .ZN(_00056_ ) );
NAND3_X1 _11137_ ( .A1(_03970_ ), .A2(\BTB.jsnpc_reg[0][6] ), .A3(_03967_ ), .ZN(_04001_ ) );
OAI21_X1 _11138_ ( .A(_04001_ ), .B1(_03812_ ), .B2(_03969_ ), .ZN(_00057_ ) );
NAND2_X1 _11139_ ( .A1(_03956_ ), .A2(\BTB.bindex_pre ), .ZN(_04002_ ) );
BUF_X4 _11140_ ( .A(_04002_ ), .Z(_04003_ ) );
BUF_X4 _11141_ ( .A(_04003_ ), .Z(_04004_ ) );
INV_X1 _11142_ ( .A(\BTB.jsnpc_reg[1][15] ), .ZN(_04005_ ) );
NAND2_X2 _11143_ ( .A1(_04002_ ), .A2(_03844_ ), .ZN(_04006_ ) );
OAI22_X1 _11144_ ( .A1(_03955_ ), .A2(_04004_ ), .B1(_04005_ ), .B2(_04006_ ), .ZN(_00058_ ) );
BUF_X4 _11145_ ( .A(_04002_ ), .Z(_04007_ ) );
INV_X1 _11146_ ( .A(\BTB.jsnpc_reg[1][14] ), .ZN(_04008_ ) );
OAI22_X1 _11147_ ( .A1(_03964_ ), .A2(_04007_ ), .B1(_04008_ ), .B2(_04006_ ), .ZN(_00059_ ) );
NAND3_X1 _11148_ ( .A1(_04007_ ), .A2(\BTB.jsnpc_reg[1][5] ), .A3(_03967_ ), .ZN(_04009_ ) );
BUF_X4 _11149_ ( .A(_04003_ ), .Z(_04010_ ) );
OAI21_X1 _11150_ ( .A(_04009_ ), .B1(_03817_ ), .B2(_04010_ ), .ZN(_00060_ ) );
BUF_X4 _11151_ ( .A(_04002_ ), .Z(_04011_ ) );
NAND3_X1 _11152_ ( .A1(_04011_ ), .A2(\BTB.jsnpc_reg[1][4] ), .A3(_03967_ ), .ZN(_04012_ ) );
OAI21_X1 _11153_ ( .A(_04012_ ), .B1(_03822_ ), .B2(_04010_ ), .ZN(_00061_ ) );
NAND3_X1 _11154_ ( .A1(_04011_ ), .A2(\BTB.jsnpc_reg[1][3] ), .A3(_03967_ ), .ZN(_04013_ ) );
OAI21_X1 _11155_ ( .A(_04013_ ), .B1(_03825_ ), .B2(_04010_ ), .ZN(_00062_ ) );
NAND3_X1 _11156_ ( .A1(_04011_ ), .A2(\BTB.jsnpc_reg[1][2] ), .A3(_03967_ ), .ZN(_04014_ ) );
OAI21_X1 _11157_ ( .A(_04014_ ), .B1(_03828_ ), .B2(_04010_ ), .ZN(_00063_ ) );
INV_X1 _11158_ ( .A(\BTB.jsnpc_reg[1][1] ), .ZN(_04015_ ) );
OAI22_X1 _11159_ ( .A1(_03830_ ), .A2(_04007_ ), .B1(_04015_ ), .B2(_04006_ ), .ZN(_00064_ ) );
INV_X1 _11160_ ( .A(\BTB.jsnpc_reg[1][0] ), .ZN(_04016_ ) );
OAI22_X1 _11161_ ( .A1(_03837_ ), .A2(_04007_ ), .B1(_04016_ ), .B2(_04006_ ), .ZN(_00065_ ) );
INV_X1 _11162_ ( .A(\BTB.jsnpc_reg[1][13] ), .ZN(_04017_ ) );
OAI22_X1 _11163_ ( .A1(_03980_ ), .A2(_04007_ ), .B1(_04017_ ), .B2(_04006_ ), .ZN(_00066_ ) );
INV_X1 _11164_ ( .A(\BTB.jsnpc_reg[1][12] ), .ZN(_04018_ ) );
OAI22_X1 _11165_ ( .A1(_03983_ ), .A2(_04007_ ), .B1(_04018_ ), .B2(_04006_ ), .ZN(_00067_ ) );
INV_X1 _11166_ ( .A(\BTB.jsnpc_reg[1][11] ), .ZN(_04019_ ) );
OAI22_X1 _11167_ ( .A1(_03987_ ), .A2(_04007_ ), .B1(_04019_ ), .B2(_04006_ ), .ZN(_00068_ ) );
INV_X1 _11168_ ( .A(\BTB.jsnpc_reg[1][10] ), .ZN(_04020_ ) );
OAI22_X1 _11169_ ( .A1(_03990_ ), .A2(_04007_ ), .B1(_04020_ ), .B2(_04006_ ), .ZN(_00069_ ) );
INV_X1 _11170_ ( .A(\BTB.jsnpc_reg[1][9] ), .ZN(_04021_ ) );
OAI22_X1 _11171_ ( .A1(_03994_ ), .A2(_04007_ ), .B1(_04021_ ), .B2(_04006_ ), .ZN(_00070_ ) );
INV_X1 _11172_ ( .A(\BTB.jsnpc_reg[1][8] ), .ZN(_04022_ ) );
OAI22_X1 _11173_ ( .A1(_03998_ ), .A2(_04007_ ), .B1(_04022_ ), .B2(_04006_ ), .ZN(_00071_ ) );
BUF_X4 _11174_ ( .A(_03808_ ), .Z(_04023_ ) );
NAND3_X1 _11175_ ( .A1(_04011_ ), .A2(\BTB.jsnpc_reg[1][7] ), .A3(_04023_ ), .ZN(_04024_ ) );
OAI21_X1 _11176_ ( .A(_04024_ ), .B1(_03842_ ), .B2(_04010_ ), .ZN(_00072_ ) );
NAND3_X1 _11177_ ( .A1(_04011_ ), .A2(\BTB.jsnpc_reg[1][6] ), .A3(_04023_ ), .ZN(_04025_ ) );
OAI21_X1 _11178_ ( .A(_04025_ ), .B1(_03812_ ), .B2(_04010_ ), .ZN(_00073_ ) );
NAND3_X1 _11179_ ( .A1(_03970_ ), .A2(\BTB.jtag_reg[0][12] ), .A3(_04023_ ), .ZN(_04026_ ) );
OAI21_X1 _11180_ ( .A(_04026_ ), .B1(_03856_ ), .B2(_03969_ ), .ZN(_00074_ ) );
NAND3_X1 _11181_ ( .A1(_03970_ ), .A2(\BTB.jtag_reg[0][11] ), .A3(_04023_ ), .ZN(_04027_ ) );
OAI21_X1 _11182_ ( .A(_04027_ ), .B1(_03858_ ), .B2(_03969_ ), .ZN(_00075_ ) );
NAND3_X1 _11183_ ( .A1(_03970_ ), .A2(\BTB.jtag_reg[0][2] ), .A3(_04023_ ), .ZN(_04028_ ) );
OAI21_X1 _11184_ ( .A(_04028_ ), .B1(_03860_ ), .B2(_03969_ ), .ZN(_00076_ ) );
NAND3_X1 _11185_ ( .A1(_03970_ ), .A2(\BTB.jtag_reg[0][1] ), .A3(_04023_ ), .ZN(_04029_ ) );
OAI21_X1 _11186_ ( .A(_04029_ ), .B1(_03862_ ), .B2(_03969_ ), .ZN(_00077_ ) );
NAND3_X1 _11187_ ( .A1(_03970_ ), .A2(\BTB.jtag_reg[0][0] ), .A3(_04023_ ), .ZN(_04030_ ) );
OAI21_X1 _11188_ ( .A(_04030_ ), .B1(_03864_ ), .B2(_03959_ ), .ZN(_00078_ ) );
NAND3_X1 _11189_ ( .A1(_03958_ ), .A2(\BTB.jtag_reg[0][10] ), .A3(_04023_ ), .ZN(_04031_ ) );
OAI21_X1 _11190_ ( .A(_04031_ ), .B1(_03867_ ), .B2(_03959_ ), .ZN(_00079_ ) );
NAND3_X1 _11191_ ( .A1(_03958_ ), .A2(\BTB.jtag_reg[0][9] ), .A3(_04023_ ), .ZN(_04032_ ) );
OAI21_X1 _11192_ ( .A(_04032_ ), .B1(_03869_ ), .B2(_03959_ ), .ZN(_00080_ ) );
NAND3_X1 _11193_ ( .A1(_03958_ ), .A2(\BTB.jtag_reg[0][8] ), .A3(_04023_ ), .ZN(_04033_ ) );
OAI21_X1 _11194_ ( .A(_04033_ ), .B1(_03871_ ), .B2(_03959_ ), .ZN(_00081_ ) );
BUF_X4 _11195_ ( .A(_03808_ ), .Z(_04034_ ) );
NAND3_X1 _11196_ ( .A1(_03958_ ), .A2(\BTB.jtag_reg[0][7] ), .A3(_04034_ ), .ZN(_04035_ ) );
OAI21_X1 _11197_ ( .A(_04035_ ), .B1(_03873_ ), .B2(_03959_ ), .ZN(_00082_ ) );
NAND3_X1 _11198_ ( .A1(_03958_ ), .A2(\BTB.jtag_reg[0][6] ), .A3(_04034_ ), .ZN(_04036_ ) );
OAI21_X1 _11199_ ( .A(_04036_ ), .B1(_03875_ ), .B2(_03959_ ), .ZN(_00083_ ) );
NAND3_X1 _11200_ ( .A1(_03958_ ), .A2(\BTB.jtag_reg[0][5] ), .A3(_04034_ ), .ZN(_04037_ ) );
OAI21_X1 _11201_ ( .A(_04037_ ), .B1(_03877_ ), .B2(_03959_ ), .ZN(_00084_ ) );
NAND3_X1 _11202_ ( .A1(_03958_ ), .A2(\BTB.jtag_reg[0][4] ), .A3(_04034_ ), .ZN(_04038_ ) );
OAI21_X1 _11203_ ( .A(_04038_ ), .B1(_03895_ ), .B2(_03959_ ), .ZN(_00085_ ) );
NAND3_X1 _11204_ ( .A1(_03958_ ), .A2(\BTB.jtag_reg[0][3] ), .A3(_04034_ ), .ZN(_04039_ ) );
OAI21_X1 _11205_ ( .A(_04039_ ), .B1(_03750_ ), .B2(_03959_ ), .ZN(_00086_ ) );
NAND3_X1 _11206_ ( .A1(_04011_ ), .A2(\BTB.jtag_reg[1][12] ), .A3(_04034_ ), .ZN(_04040_ ) );
OAI21_X1 _11207_ ( .A(_04040_ ), .B1(_03856_ ), .B2(_04010_ ), .ZN(_00087_ ) );
NAND3_X1 _11208_ ( .A1(_04011_ ), .A2(\BTB.jtag_reg[1][11] ), .A3(_04034_ ), .ZN(_04041_ ) );
OAI21_X1 _11209_ ( .A(_04041_ ), .B1(_03858_ ), .B2(_04010_ ), .ZN(_00088_ ) );
NAND3_X1 _11210_ ( .A1(_04011_ ), .A2(\BTB.jtag_reg[1][2] ), .A3(_04034_ ), .ZN(_04042_ ) );
OAI21_X1 _11211_ ( .A(_04042_ ), .B1(_03860_ ), .B2(_04010_ ), .ZN(_00089_ ) );
NAND3_X1 _11212_ ( .A1(_04011_ ), .A2(\BTB.jtag_reg[1][1] ), .A3(_04034_ ), .ZN(_04043_ ) );
OAI21_X1 _11213_ ( .A(_04043_ ), .B1(_03862_ ), .B2(_04010_ ), .ZN(_00090_ ) );
NAND3_X1 _11214_ ( .A1(_04011_ ), .A2(\BTB.jtag_reg[1][0] ), .A3(_04034_ ), .ZN(_04044_ ) );
OAI21_X1 _11215_ ( .A(_04044_ ), .B1(_03864_ ), .B2(_04004_ ), .ZN(_00091_ ) );
BUF_X4 _11216_ ( .A(_03808_ ), .Z(_04045_ ) );
NAND3_X1 _11217_ ( .A1(_04003_ ), .A2(\BTB.jtag_reg[1][10] ), .A3(_04045_ ), .ZN(_04046_ ) );
OAI21_X1 _11218_ ( .A(_04046_ ), .B1(_03867_ ), .B2(_04004_ ), .ZN(_00092_ ) );
NAND3_X1 _11219_ ( .A1(_04003_ ), .A2(\BTB.jtag_reg[1][9] ), .A3(_04045_ ), .ZN(_04047_ ) );
OAI21_X1 _11220_ ( .A(_04047_ ), .B1(_03869_ ), .B2(_04004_ ), .ZN(_00093_ ) );
NAND3_X1 _11221_ ( .A1(_04003_ ), .A2(\BTB.jtag_reg[1][8] ), .A3(_04045_ ), .ZN(_04048_ ) );
OAI21_X1 _11222_ ( .A(_04048_ ), .B1(_03871_ ), .B2(_04004_ ), .ZN(_00094_ ) );
NAND3_X1 _11223_ ( .A1(_04003_ ), .A2(\BTB.jtag_reg[1][7] ), .A3(_04045_ ), .ZN(_04049_ ) );
OAI21_X1 _11224_ ( .A(_04049_ ), .B1(_03873_ ), .B2(_04004_ ), .ZN(_00095_ ) );
NAND3_X1 _11225_ ( .A1(_04003_ ), .A2(\BTB.jtag_reg[1][6] ), .A3(_04045_ ), .ZN(_04050_ ) );
OAI21_X1 _11226_ ( .A(_04050_ ), .B1(_03875_ ), .B2(_04004_ ), .ZN(_00096_ ) );
NAND3_X1 _11227_ ( .A1(_04003_ ), .A2(\BTB.jtag_reg[1][5] ), .A3(_04045_ ), .ZN(_04051_ ) );
OAI21_X1 _11228_ ( .A(_04051_ ), .B1(_03877_ ), .B2(_04004_ ), .ZN(_00097_ ) );
NAND3_X1 _11229_ ( .A1(_04003_ ), .A2(\BTB.jtag_reg[1][4] ), .A3(_04045_ ), .ZN(_04052_ ) );
OAI21_X1 _11230_ ( .A(_04052_ ), .B1(_03895_ ), .B2(_04004_ ), .ZN(_00098_ ) );
NAND3_X1 _11231_ ( .A1(_04003_ ), .A2(\BTB.jtag_reg[1][3] ), .A3(_04045_ ), .ZN(_04053_ ) );
OAI21_X1 _11232_ ( .A(_04053_ ), .B1(_03750_ ), .B2(_04004_ ), .ZN(_00099_ ) );
OAI21_X1 _11233_ ( .A(\Xbar.state [0] ), .B1(\LSU.ls_axi_arvalid ), .B2(\LSU.ls_axi_awvalid ), .ZN(_04054_ ) );
INV_X1 _11234_ ( .A(_04054_ ), .ZN(_04055_ ) );
NOR2_X1 _11235_ ( .A1(_04055_ ), .A2(\Xbar.state [2] ), .ZN(_04056_ ) );
BUF_X4 _11236_ ( .A(_04056_ ), .Z(_04057_ ) );
BUF_X4 _11237_ ( .A(_04057_ ), .Z(_04058_ ) );
MUX2_X1 _11238_ ( .A(\LSU.ls_axi_araddr [9] ), .B(\ICACHE.s_axi_araddr [9] ), .S(_04058_ ), .Z(\io_master_araddr [9] ) );
BUF_X4 _11239_ ( .A(_04056_ ), .Z(_04059_ ) );
BUF_X4 _11240_ ( .A(_04059_ ), .Z(_04060_ ) );
MUX2_X1 _11241_ ( .A(\LSU.ls_axi_araddr [8] ), .B(\ICACHE.s_axi_araddr [8] ), .S(_04060_ ), .Z(\io_master_araddr [8] ) );
MUX2_X1 _11242_ ( .A(\LSU.ls_axi_araddr [11] ), .B(\ICACHE.s_axi_araddr [11] ), .S(_04060_ ), .Z(\io_master_araddr [11] ) );
MUX2_X1 _11243_ ( .A(\LSU.ls_axi_araddr [10] ), .B(\ICACHE.s_axi_araddr [10] ), .S(_04057_ ), .Z(\io_master_araddr [10] ) );
NOR4_X1 _11244_ ( .A1(\io_master_araddr [9] ), .A2(\io_master_araddr [8] ), .A3(\io_master_araddr [11] ), .A4(\io_master_araddr [10] ), .ZN(_04061_ ) );
MUX2_X1 _11245_ ( .A(\LSU.ls_axi_araddr [13] ), .B(\ICACHE.s_axi_araddr [13] ), .S(_04060_ ), .Z(\io_master_araddr [13] ) );
MUX2_X1 _11246_ ( .A(\LSU.ls_axi_araddr [12] ), .B(\ICACHE.s_axi_araddr [12] ), .S(_04060_ ), .Z(\io_master_araddr [12] ) );
MUX2_X1 _11247_ ( .A(\LSU.ls_axi_araddr [15] ), .B(\ICACHE.s_axi_araddr [15] ), .S(_04057_ ), .Z(\io_master_araddr [15] ) );
MUX2_X1 _11248_ ( .A(\LSU.ls_axi_araddr [14] ), .B(\ICACHE.s_axi_araddr [14] ), .S(_04057_ ), .Z(\io_master_araddr [14] ) );
NOR4_X1 _11249_ ( .A1(\io_master_araddr [13] ), .A2(\io_master_araddr [12] ), .A3(\io_master_araddr [15] ), .A4(\io_master_araddr [14] ), .ZN(_04062_ ) );
NAND2_X1 _11250_ ( .A1(_04061_ ), .A2(_04062_ ), .ZN(_04063_ ) );
MUX2_X1 _11251_ ( .A(\LSU.ls_axi_araddr [1] ), .B(\ICACHE.s_axi_araddr [1] ), .S(_04058_ ), .Z(\io_master_araddr [1] ) );
MUX2_X1 _11252_ ( .A(\LSU.ls_axi_araddr [0] ), .B(\ICACHE.s_axi_araddr [0] ), .S(_04060_ ), .Z(\io_master_araddr [0] ) );
NOR2_X1 _11253_ ( .A1(\io_master_araddr [1] ), .A2(\io_master_araddr [0] ), .ZN(_04064_ ) );
MUX2_X1 _11254_ ( .A(\LSU.ls_axi_araddr [7] ), .B(\ICACHE.s_axi_araddr [7] ), .S(_04060_ ), .Z(\io_master_araddr [7] ) );
MUX2_X1 _11255_ ( .A(\LSU.ls_axi_araddr [6] ), .B(\ICACHE.s_axi_araddr [6] ), .S(_04060_ ), .Z(\io_master_araddr [6] ) );
NOR2_X1 _11256_ ( .A1(\io_master_araddr [7] ), .A2(\io_master_araddr [6] ), .ZN(_04065_ ) );
MUX2_X1 _11257_ ( .A(\LSU.ls_axi_araddr [5] ), .B(\ICACHE.s_axi_araddr [5] ), .S(_04060_ ), .Z(\io_master_araddr [5] ) );
MUX2_X1 _11258_ ( .A(\LSU.ls_axi_araddr [4] ), .B(\ICACHE.s_axi_araddr [4] ), .S(_04060_ ), .Z(\io_master_araddr [4] ) );
NOR2_X1 _11259_ ( .A1(\io_master_araddr [5] ), .A2(\io_master_araddr [4] ), .ZN(_04066_ ) );
MUX2_X1 _11260_ ( .A(\LSU.ls_axi_araddr [3] ), .B(\ICACHE.s_axi_araddr [3] ), .S(_04060_ ), .Z(\io_master_araddr [3] ) );
NAND2_X1 _11261_ ( .A1(_04058_ ), .A2(\ICACHE.s_axi_araddr [2] ), .ZN(_04067_ ) );
OAI21_X1 _11262_ ( .A(\LSU.ls_axi_araddr [2] ), .B1(_04055_ ), .B2(\Xbar.state [2] ), .ZN(_04068_ ) );
NAND2_X1 _11263_ ( .A1(_04067_ ), .A2(_04068_ ), .ZN(_04069_ ) );
INV_X1 _11264_ ( .A(_04069_ ), .ZN(_04070_ ) );
NOR2_X1 _11265_ ( .A1(\io_master_araddr [3] ), .A2(_04070_ ), .ZN(_04071_ ) );
NAND4_X1 _11266_ ( .A1(_04064_ ), .A2(_04065_ ), .A3(_04066_ ), .A4(_04071_ ), .ZN(_04072_ ) );
NOR2_X1 _11267_ ( .A1(_04063_ ), .A2(_04072_ ), .ZN(_04073_ ) );
BUF_X4 _11268_ ( .A(_04073_ ), .Z(_04074_ ) );
BUF_X4 _11269_ ( .A(_04074_ ), .Z(_04075_ ) );
BUF_X4 _11270_ ( .A(_04075_ ), .Z(_04076_ ) );
BUF_X4 _11271_ ( .A(_04076_ ), .Z(_04077_ ) );
MUX2_X1 _11272_ ( .A(\LSU.ls_axi_araddr [29] ), .B(\ICACHE.s_axi_araddr [29] ), .S(_04057_ ), .Z(\io_master_araddr [29] ) );
MUX2_X1 _11273_ ( .A(\LSU.ls_axi_araddr [28] ), .B(\ICACHE.s_axi_araddr [28] ), .S(_04059_ ), .Z(\io_master_araddr [28] ) );
MUX2_X1 _11274_ ( .A(\LSU.ls_axi_araddr [31] ), .B(\ICACHE.s_axi_araddr [31] ), .S(_04059_ ), .Z(\io_master_araddr [31] ) );
MUX2_X1 _11275_ ( .A(\LSU.ls_axi_araddr [30] ), .B(\ICACHE.s_axi_araddr [30] ), .S(_04059_ ), .Z(\io_master_araddr [30] ) );
OR4_X1 _11276_ ( .A1(\io_master_araddr [29] ), .A2(\io_master_araddr [28] ), .A3(\io_master_araddr [31] ), .A4(\io_master_araddr [30] ), .ZN(_04078_ ) );
MUX2_X1 _11277_ ( .A(\LSU.ls_axi_araddr [26] ), .B(\ICACHE.s_axi_araddr [26] ), .S(_04059_ ), .Z(\io_master_araddr [26] ) );
MUX2_X1 _11278_ ( .A(\LSU.ls_axi_araddr [27] ), .B(\ICACHE.s_axi_araddr [27] ), .S(_04059_ ), .Z(\io_master_araddr [27] ) );
MUX2_X1 _11279_ ( .A(\LSU.ls_axi_araddr [24] ), .B(\ICACHE.s_axi_araddr [24] ), .S(_04056_ ), .Z(\io_master_araddr [24] ) );
NAND2_X1 _11280_ ( .A1(_04059_ ), .A2(\ICACHE.s_axi_araddr [25] ), .ZN(_04079_ ) );
OAI21_X1 _11281_ ( .A(\LSU.ls_axi_araddr [25] ), .B1(_04055_ ), .B2(\Xbar.state [2] ), .ZN(_04080_ ) );
NAND2_X1 _11282_ ( .A1(_04079_ ), .A2(_04080_ ), .ZN(_04081_ ) );
INV_X1 _11283_ ( .A(_04081_ ), .ZN(_04082_ ) );
OR4_X1 _11284_ ( .A1(\io_master_araddr [26] ), .A2(\io_master_araddr [27] ), .A3(\io_master_araddr [24] ), .A4(_04082_ ), .ZN(_04083_ ) );
MUX2_X1 _11285_ ( .A(\LSU.ls_axi_araddr [19] ), .B(\ICACHE.s_axi_araddr [19] ), .S(_04057_ ), .Z(\io_master_araddr [19] ) );
MUX2_X1 _11286_ ( .A(\LSU.ls_axi_araddr [18] ), .B(\ICACHE.s_axi_araddr [18] ), .S(_04057_ ), .Z(\io_master_araddr [18] ) );
NOR2_X1 _11287_ ( .A1(\io_master_araddr [19] ), .A2(\io_master_araddr [18] ), .ZN(_04084_ ) );
MUX2_X1 _11288_ ( .A(\LSU.ls_axi_araddr [21] ), .B(\ICACHE.s_axi_araddr [21] ), .S(_04057_ ), .Z(\io_master_araddr [21] ) );
MUX2_X1 _11289_ ( .A(\LSU.ls_axi_araddr [20] ), .B(\ICACHE.s_axi_araddr [20] ), .S(_04059_ ), .Z(\io_master_araddr [20] ) );
NOR2_X1 _11290_ ( .A1(\io_master_araddr [21] ), .A2(\io_master_araddr [20] ), .ZN(_04085_ ) );
MUX2_X1 _11291_ ( .A(\LSU.ls_axi_araddr [17] ), .B(\ICACHE.s_axi_araddr [17] ), .S(_04057_ ), .Z(\io_master_araddr [17] ) );
MUX2_X1 _11292_ ( .A(\LSU.ls_axi_araddr [16] ), .B(\ICACHE.s_axi_araddr [16] ), .S(_04059_ ), .Z(\io_master_araddr [16] ) );
NOR2_X1 _11293_ ( .A1(\io_master_araddr [17] ), .A2(\io_master_araddr [16] ), .ZN(_04086_ ) );
MUX2_X1 _11294_ ( .A(\LSU.ls_axi_araddr [23] ), .B(\ICACHE.s_axi_araddr [23] ), .S(_04057_ ), .Z(\io_master_araddr [23] ) );
MUX2_X1 _11295_ ( .A(\LSU.ls_axi_araddr [22] ), .B(\ICACHE.s_axi_araddr [22] ), .S(_04059_ ), .Z(\io_master_araddr [22] ) );
NOR2_X1 _11296_ ( .A1(\io_master_araddr [23] ), .A2(\io_master_araddr [22] ), .ZN(_04087_ ) );
NAND4_X1 _11297_ ( .A1(_04084_ ), .A2(_04085_ ), .A3(_04086_ ), .A4(_04087_ ), .ZN(_04088_ ) );
NOR3_X2 _11298_ ( .A1(_04078_ ), .A2(_04083_ ), .A3(_04088_ ), .ZN(_04089_ ) );
BUF_X4 _11299_ ( .A(_04089_ ), .Z(_04090_ ) );
BUF_X4 _11300_ ( .A(_04090_ ), .Z(_04091_ ) );
BUF_X4 _11301_ ( .A(_04091_ ), .Z(_04092_ ) );
BUF_X4 _11302_ ( .A(_04092_ ), .Z(_04093_ ) );
NAND3_X1 _11303_ ( .A1(_04077_ ), .A2(_04093_ ), .A3(\CLINT.mtime [63] ), .ZN(_04094_ ) );
NOR2_X1 _11304_ ( .A1(\io_master_araddr [3] ), .A2(_04069_ ), .ZN(_04095_ ) );
NAND4_X1 _11305_ ( .A1(_04064_ ), .A2(_04065_ ), .A3(_04066_ ), .A4(_04095_ ), .ZN(_04096_ ) );
NOR2_X1 _11306_ ( .A1(_04063_ ), .A2(_04096_ ), .ZN(_04097_ ) );
BUF_X4 _11307_ ( .A(_04097_ ), .Z(_04098_ ) );
BUF_X4 _11308_ ( .A(_04098_ ), .Z(_04099_ ) );
BUF_X4 _11309_ ( .A(_04099_ ), .Z(_04100_ ) );
BUF_X4 _11310_ ( .A(_04100_ ), .Z(_04101_ ) );
BUF_X4 _11311_ ( .A(_04092_ ), .Z(_04102_ ) );
NAND3_X1 _11312_ ( .A1(_04101_ ), .A2(_04102_ ), .A3(\CLINT.mtime [31] ), .ZN(_04103_ ) );
NAND2_X1 _11313_ ( .A1(_04094_ ), .A2(_04103_ ), .ZN(_04104_ ) );
BUF_X4 _11314_ ( .A(_04058_ ), .Z(_04105_ ) );
NOR2_X1 _11315_ ( .A1(_04105_ ), .A2(io_master_arvalid_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_04106_ ) );
NOR3_X1 _11316_ ( .A1(_04055_ ), .A2(\Xbar.state [2] ), .A3(io_master_arvalid_$_ANDNOT__Y_B_$_MUX__Y_A ), .ZN(_04107_ ) );
OAI21_X1 _11317_ ( .A(\CLINT.c_axi_arready ), .B1(_04106_ ), .B2(_04107_ ), .ZN(_04108_ ) );
AND2_X1 _11318_ ( .A1(_04073_ ), .A2(_04089_ ), .ZN(_04109_ ) );
BUF_X2 _11319_ ( .A(_04109_ ), .Z(_04110_ ) );
INV_X1 _11320_ ( .A(_04110_ ), .ZN(_04111_ ) );
AND2_X1 _11321_ ( .A1(_04097_ ), .A2(_04089_ ), .ZN(_04112_ ) );
BUF_X2 _11322_ ( .A(_04112_ ), .Z(_04113_ ) );
INV_X1 _11323_ ( .A(_04113_ ), .ZN(_04114_ ) );
AOI21_X1 _11324_ ( .A(_04108_ ), .B1(_04111_ ), .B2(_04114_ ), .ZN(_04115_ ) );
AND2_X2 _11325_ ( .A1(_04115_ ), .A2(_03805_ ), .ZN(_04116_ ) );
BUF_X4 _11326_ ( .A(_04116_ ), .Z(_04117_ ) );
MUX2_X1 _11327_ ( .A(\CLINT.c_axi_rdata [31] ), .B(_04104_ ), .S(_04117_ ), .Z(_00100_ ) );
NAND3_X1 _11328_ ( .A1(_04077_ ), .A2(_04093_ ), .A3(\CLINT.mtime [62] ), .ZN(_04118_ ) );
NAND3_X1 _11329_ ( .A1(_04101_ ), .A2(_04102_ ), .A3(\CLINT.mtime [30] ), .ZN(_04119_ ) );
NAND2_X1 _11330_ ( .A1(_04118_ ), .A2(_04119_ ), .ZN(_04120_ ) );
MUX2_X1 _11331_ ( .A(\CLINT.c_axi_rdata [30] ), .B(_04120_ ), .S(_04117_ ), .Z(_00101_ ) );
NAND3_X1 _11332_ ( .A1(_04077_ ), .A2(_04093_ ), .A3(\CLINT.mtime [53] ), .ZN(_04121_ ) );
NAND3_X1 _11333_ ( .A1(_04101_ ), .A2(_04102_ ), .A3(\CLINT.mtime [21] ), .ZN(_04122_ ) );
NAND2_X1 _11334_ ( .A1(_04121_ ), .A2(_04122_ ), .ZN(_04123_ ) );
MUX2_X1 _11335_ ( .A(\CLINT.c_axi_rdata [21] ), .B(_04123_ ), .S(_04117_ ), .Z(_00102_ ) );
NAND3_X1 _11336_ ( .A1(_04077_ ), .A2(_04093_ ), .A3(\CLINT.mtime [52] ), .ZN(_04124_ ) );
NAND3_X1 _11337_ ( .A1(_04101_ ), .A2(_04102_ ), .A3(\CLINT.mtime [20] ), .ZN(_04125_ ) );
NAND2_X1 _11338_ ( .A1(_04124_ ), .A2(_04125_ ), .ZN(_04126_ ) );
MUX2_X1 _11339_ ( .A(\CLINT.c_axi_rdata [20] ), .B(_04126_ ), .S(_04117_ ), .Z(_00103_ ) );
NAND3_X1 _11340_ ( .A1(_04077_ ), .A2(_04093_ ), .A3(\CLINT.mtime [51] ), .ZN(_04127_ ) );
NAND3_X1 _11341_ ( .A1(_04101_ ), .A2(_04102_ ), .A3(\CLINT.mtime [19] ), .ZN(_04128_ ) );
NAND2_X1 _11342_ ( .A1(_04127_ ), .A2(_04128_ ), .ZN(_04129_ ) );
MUX2_X1 _11343_ ( .A(\CLINT.c_axi_rdata [19] ), .B(_04129_ ), .S(_04117_ ), .Z(_00104_ ) );
NAND3_X1 _11344_ ( .A1(_04077_ ), .A2(_04093_ ), .A3(\CLINT.mtime [50] ), .ZN(_04130_ ) );
NAND3_X1 _11345_ ( .A1(_04101_ ), .A2(_04102_ ), .A3(\CLINT.mtime [18] ), .ZN(_04131_ ) );
NAND2_X1 _11346_ ( .A1(_04130_ ), .A2(_04131_ ), .ZN(_04132_ ) );
MUX2_X1 _11347_ ( .A(\CLINT.c_axi_rdata [18] ), .B(_04132_ ), .S(_04117_ ), .Z(_00105_ ) );
NAND3_X1 _11348_ ( .A1(_04077_ ), .A2(_04093_ ), .A3(\CLINT.mtime [49] ), .ZN(_04133_ ) );
BUF_X4 _11349_ ( .A(_04092_ ), .Z(_04134_ ) );
NAND3_X1 _11350_ ( .A1(_04101_ ), .A2(_04134_ ), .A3(\CLINT.mtime [17] ), .ZN(_04135_ ) );
NAND2_X1 _11351_ ( .A1(_04133_ ), .A2(_04135_ ), .ZN(_04136_ ) );
MUX2_X1 _11352_ ( .A(\CLINT.c_axi_rdata [17] ), .B(_04136_ ), .S(_04117_ ), .Z(_00106_ ) );
NAND3_X1 _11353_ ( .A1(_04077_ ), .A2(_04093_ ), .A3(\CLINT.mtime [48] ), .ZN(_04137_ ) );
NAND3_X1 _11354_ ( .A1(_04101_ ), .A2(_04134_ ), .A3(\CLINT.mtime [16] ), .ZN(_04138_ ) );
NAND2_X1 _11355_ ( .A1(_04137_ ), .A2(_04138_ ), .ZN(_04139_ ) );
MUX2_X1 _11356_ ( .A(\CLINT.c_axi_rdata [16] ), .B(_04139_ ), .S(_04117_ ), .Z(_00107_ ) );
BUF_X4 _11357_ ( .A(_04076_ ), .Z(_04140_ ) );
BUF_X4 _11358_ ( .A(_04092_ ), .Z(_04141_ ) );
NAND3_X1 _11359_ ( .A1(_04140_ ), .A2(_04141_ ), .A3(\CLINT.mtime [47] ), .ZN(_04142_ ) );
BUF_X4 _11360_ ( .A(_04100_ ), .Z(_04143_ ) );
NAND3_X1 _11361_ ( .A1(_04143_ ), .A2(_04134_ ), .A3(\CLINT.mtime [15] ), .ZN(_04144_ ) );
NAND2_X1 _11362_ ( .A1(_04142_ ), .A2(_04144_ ), .ZN(_04145_ ) );
BUF_X4 _11363_ ( .A(_04116_ ), .Z(_04146_ ) );
MUX2_X1 _11364_ ( .A(\CLINT.c_axi_rdata [15] ), .B(_04145_ ), .S(_04146_ ), .Z(_00108_ ) );
NAND3_X1 _11365_ ( .A1(_04140_ ), .A2(_04141_ ), .A3(\CLINT.mtime [46] ), .ZN(_04147_ ) );
NAND3_X1 _11366_ ( .A1(_04143_ ), .A2(_04134_ ), .A3(\CLINT.mtime [14] ), .ZN(_04148_ ) );
NAND2_X1 _11367_ ( .A1(_04147_ ), .A2(_04148_ ), .ZN(_04149_ ) );
MUX2_X1 _11368_ ( .A(\CLINT.c_axi_rdata [14] ), .B(_04149_ ), .S(_04146_ ), .Z(_00109_ ) );
NAND3_X1 _11369_ ( .A1(_04140_ ), .A2(_04141_ ), .A3(\CLINT.mtime [45] ), .ZN(_04150_ ) );
NAND3_X1 _11370_ ( .A1(_04143_ ), .A2(_04134_ ), .A3(\CLINT.mtime [13] ), .ZN(_04151_ ) );
NAND2_X1 _11371_ ( .A1(_04150_ ), .A2(_04151_ ), .ZN(_04152_ ) );
MUX2_X1 _11372_ ( .A(\CLINT.c_axi_rdata [13] ), .B(_04152_ ), .S(_04146_ ), .Z(_00110_ ) );
NAND3_X1 _11373_ ( .A1(_04140_ ), .A2(_04141_ ), .A3(\CLINT.mtime [44] ), .ZN(_04153_ ) );
NAND3_X1 _11374_ ( .A1(_04143_ ), .A2(_04134_ ), .A3(\CLINT.mtime [12] ), .ZN(_04154_ ) );
NAND2_X1 _11375_ ( .A1(_04153_ ), .A2(_04154_ ), .ZN(_04155_ ) );
MUX2_X1 _11376_ ( .A(\CLINT.c_axi_rdata [12] ), .B(_04155_ ), .S(_04146_ ), .Z(_00111_ ) );
NAND3_X1 _11377_ ( .A1(_04140_ ), .A2(_04141_ ), .A3(\CLINT.mtime [61] ), .ZN(_04156_ ) );
NAND3_X1 _11378_ ( .A1(_04143_ ), .A2(_04134_ ), .A3(\CLINT.mtime [29] ), .ZN(_04157_ ) );
NAND2_X1 _11379_ ( .A1(_04156_ ), .A2(_04157_ ), .ZN(_04158_ ) );
MUX2_X1 _11380_ ( .A(\CLINT.c_axi_rdata [29] ), .B(_04158_ ), .S(_04146_ ), .Z(_00112_ ) );
NAND3_X1 _11381_ ( .A1(_04140_ ), .A2(_04141_ ), .A3(\CLINT.mtime [43] ), .ZN(_04159_ ) );
NAND3_X1 _11382_ ( .A1(_04143_ ), .A2(_04134_ ), .A3(\CLINT.mtime [11] ), .ZN(_04160_ ) );
NAND2_X1 _11383_ ( .A1(_04159_ ), .A2(_04160_ ), .ZN(_04161_ ) );
MUX2_X1 _11384_ ( .A(\CLINT.c_axi_rdata [11] ), .B(_04161_ ), .S(_04146_ ), .Z(_00113_ ) );
NAND3_X1 _11385_ ( .A1(_04140_ ), .A2(_04141_ ), .A3(\CLINT.mtime [42] ), .ZN(_04162_ ) );
NAND3_X1 _11386_ ( .A1(_04143_ ), .A2(_04134_ ), .A3(\CLINT.mtime [10] ), .ZN(_04163_ ) );
NAND2_X1 _11387_ ( .A1(_04162_ ), .A2(_04163_ ), .ZN(_04164_ ) );
MUX2_X1 _11388_ ( .A(\CLINT.c_axi_rdata [10] ), .B(_04164_ ), .S(_04146_ ), .Z(_00114_ ) );
NAND3_X1 _11389_ ( .A1(_04140_ ), .A2(_04141_ ), .A3(\CLINT.mtime [41] ), .ZN(_04165_ ) );
NAND3_X1 _11390_ ( .A1(_04143_ ), .A2(_04134_ ), .A3(\CLINT.mtime [9] ), .ZN(_04166_ ) );
NAND2_X1 _11391_ ( .A1(_04165_ ), .A2(_04166_ ), .ZN(_04167_ ) );
MUX2_X1 _11392_ ( .A(\CLINT.c_axi_rdata [9] ), .B(_04167_ ), .S(_04146_ ), .Z(_00115_ ) );
NAND3_X1 _11393_ ( .A1(_04140_ ), .A2(_04141_ ), .A3(\CLINT.mtime [40] ), .ZN(_04168_ ) );
BUF_X4 _11394_ ( .A(_04092_ ), .Z(_04169_ ) );
NAND3_X1 _11395_ ( .A1(_04143_ ), .A2(_04169_ ), .A3(\CLINT.mtime [8] ), .ZN(_04170_ ) );
NAND2_X1 _11396_ ( .A1(_04168_ ), .A2(_04170_ ), .ZN(_04171_ ) );
MUX2_X1 _11397_ ( .A(\CLINT.c_axi_rdata [8] ), .B(_04171_ ), .S(_04146_ ), .Z(_00116_ ) );
NAND3_X1 _11398_ ( .A1(_04140_ ), .A2(_04141_ ), .A3(\CLINT.mtime [39] ), .ZN(_04172_ ) );
NAND3_X1 _11399_ ( .A1(_04143_ ), .A2(_04169_ ), .A3(\CLINT.mtime [7] ), .ZN(_04173_ ) );
NAND2_X1 _11400_ ( .A1(_04172_ ), .A2(_04173_ ), .ZN(_04174_ ) );
MUX2_X1 _11401_ ( .A(\CLINT.c_axi_rdata [7] ), .B(_04174_ ), .S(_04146_ ), .Z(_00117_ ) );
BUF_X4 _11402_ ( .A(_04076_ ), .Z(_04175_ ) );
BUF_X4 _11403_ ( .A(_04092_ ), .Z(_04176_ ) );
NAND3_X1 _11404_ ( .A1(_04175_ ), .A2(_04176_ ), .A3(\CLINT.mtime [38] ), .ZN(_04177_ ) );
BUF_X4 _11405_ ( .A(_04100_ ), .Z(_04178_ ) );
NAND3_X1 _11406_ ( .A1(_04178_ ), .A2(_04169_ ), .A3(\CLINT.mtime [6] ), .ZN(_04179_ ) );
NAND2_X1 _11407_ ( .A1(_04177_ ), .A2(_04179_ ), .ZN(_04180_ ) );
BUF_X4 _11408_ ( .A(_04116_ ), .Z(_04181_ ) );
MUX2_X1 _11409_ ( .A(\CLINT.c_axi_rdata [6] ), .B(_04180_ ), .S(_04181_ ), .Z(_00118_ ) );
NAND3_X1 _11410_ ( .A1(_04175_ ), .A2(_04176_ ), .A3(\CLINT.mtime [37] ), .ZN(_04182_ ) );
NAND3_X1 _11411_ ( .A1(_04178_ ), .A2(_04169_ ), .A3(\CLINT.mtime [5] ), .ZN(_04183_ ) );
NAND2_X1 _11412_ ( .A1(_04182_ ), .A2(_04183_ ), .ZN(_04184_ ) );
MUX2_X1 _11413_ ( .A(\CLINT.c_axi_rdata [5] ), .B(_04184_ ), .S(_04181_ ), .Z(_00119_ ) );
NAND3_X1 _11414_ ( .A1(_04175_ ), .A2(_04176_ ), .A3(\CLINT.mtime [36] ), .ZN(_04185_ ) );
NAND3_X1 _11415_ ( .A1(_04178_ ), .A2(_04169_ ), .A3(\CLINT.mtime [4] ), .ZN(_04186_ ) );
NAND2_X1 _11416_ ( .A1(_04185_ ), .A2(_04186_ ), .ZN(_04187_ ) );
MUX2_X1 _11417_ ( .A(\CLINT.c_axi_rdata [4] ), .B(_04187_ ), .S(_04181_ ), .Z(_00120_ ) );
NAND3_X1 _11418_ ( .A1(_04175_ ), .A2(_04176_ ), .A3(\CLINT.mtime [35] ), .ZN(_04188_ ) );
NAND3_X1 _11419_ ( .A1(_04178_ ), .A2(_04169_ ), .A3(\CLINT.mtime [3] ), .ZN(_04189_ ) );
NAND2_X1 _11420_ ( .A1(_04188_ ), .A2(_04189_ ), .ZN(_04190_ ) );
MUX2_X1 _11421_ ( .A(\CLINT.c_axi_rdata [3] ), .B(_04190_ ), .S(_04181_ ), .Z(_00121_ ) );
NAND3_X1 _11422_ ( .A1(_04175_ ), .A2(_04176_ ), .A3(\CLINT.mtime [34] ), .ZN(_04191_ ) );
NAND3_X1 _11423_ ( .A1(_04178_ ), .A2(_04169_ ), .A3(\CLINT.mtime [2] ), .ZN(_04192_ ) );
NAND2_X1 _11424_ ( .A1(_04191_ ), .A2(_04192_ ), .ZN(_04193_ ) );
MUX2_X1 _11425_ ( .A(\CLINT.c_axi_rdata [2] ), .B(_04193_ ), .S(_04181_ ), .Z(_00122_ ) );
NAND3_X1 _11426_ ( .A1(_04175_ ), .A2(_04176_ ), .A3(\CLINT.mtime [60] ), .ZN(_04194_ ) );
NAND3_X1 _11427_ ( .A1(_04178_ ), .A2(_04169_ ), .A3(\CLINT.mtime [28] ), .ZN(_04195_ ) );
NAND2_X1 _11428_ ( .A1(_04194_ ), .A2(_04195_ ), .ZN(_04196_ ) );
MUX2_X1 _11429_ ( .A(\CLINT.c_axi_rdata [28] ), .B(_04196_ ), .S(_04181_ ), .Z(_00123_ ) );
NAND3_X1 _11430_ ( .A1(_04077_ ), .A2(_04093_ ), .A3(\CLINT.mtime [33] ), .ZN(_04197_ ) );
NAND3_X1 _11431_ ( .A1(_04101_ ), .A2(_04102_ ), .A3(\CLINT.mtime [1] ), .ZN(_04198_ ) );
NAND2_X1 _11432_ ( .A1(_04197_ ), .A2(_04198_ ), .ZN(_04199_ ) );
NAND3_X1 _11433_ ( .A1(_04115_ ), .A2(_03809_ ), .A3(_04199_ ), .ZN(_04200_ ) );
INV_X1 _11434_ ( .A(\CLINT.c_axi_rdata [1] ), .ZN(_04201_ ) );
OAI21_X1 _11435_ ( .A(_04200_ ), .B1(_04117_ ), .B2(_04201_ ), .ZN(_00124_ ) );
NAND3_X1 _11436_ ( .A1(_04077_ ), .A2(_04093_ ), .A3(\CLINT.mtime [32] ), .ZN(_04202_ ) );
NAND3_X1 _11437_ ( .A1(_04101_ ), .A2(_04102_ ), .A3(\CLINT.mtime [0] ), .ZN(_04203_ ) );
NAND2_X1 _11438_ ( .A1(_04202_ ), .A2(_04203_ ), .ZN(_04204_ ) );
NAND3_X1 _11439_ ( .A1(_04115_ ), .A2(_03809_ ), .A3(_04204_ ), .ZN(_04205_ ) );
INV_X1 _11440_ ( .A(\CLINT.c_axi_rdata [0] ), .ZN(_04206_ ) );
OAI21_X1 _11441_ ( .A(_04205_ ), .B1(_04117_ ), .B2(_04206_ ), .ZN(_00125_ ) );
NAND3_X1 _11442_ ( .A1(_04175_ ), .A2(_04176_ ), .A3(\CLINT.mtime [59] ), .ZN(_04207_ ) );
NAND3_X1 _11443_ ( .A1(_04178_ ), .A2(_04169_ ), .A3(\CLINT.mtime [27] ), .ZN(_04208_ ) );
NAND2_X1 _11444_ ( .A1(_04207_ ), .A2(_04208_ ), .ZN(_04209_ ) );
MUX2_X1 _11445_ ( .A(\CLINT.c_axi_rdata [27] ), .B(_04209_ ), .S(_04181_ ), .Z(_00126_ ) );
NAND3_X1 _11446_ ( .A1(_04175_ ), .A2(_04176_ ), .A3(\CLINT.mtime [58] ), .ZN(_04210_ ) );
NAND3_X1 _11447_ ( .A1(_04178_ ), .A2(_04169_ ), .A3(\CLINT.mtime [26] ), .ZN(_04211_ ) );
NAND2_X1 _11448_ ( .A1(_04210_ ), .A2(_04211_ ), .ZN(_04212_ ) );
MUX2_X1 _11449_ ( .A(\CLINT.c_axi_rdata [26] ), .B(_04212_ ), .S(_04181_ ), .Z(_00127_ ) );
NAND3_X1 _11450_ ( .A1(_04175_ ), .A2(_04176_ ), .A3(\CLINT.mtime [57] ), .ZN(_04213_ ) );
NAND3_X1 _11451_ ( .A1(_04178_ ), .A2(_04092_ ), .A3(\CLINT.mtime [25] ), .ZN(_04214_ ) );
NAND2_X1 _11452_ ( .A1(_04213_ ), .A2(_04214_ ), .ZN(_04215_ ) );
MUX2_X1 _11453_ ( .A(\CLINT.c_axi_rdata [25] ), .B(_04215_ ), .S(_04181_ ), .Z(_00128_ ) );
NAND3_X1 _11454_ ( .A1(_04175_ ), .A2(_04176_ ), .A3(\CLINT.mtime [56] ), .ZN(_04216_ ) );
NAND3_X1 _11455_ ( .A1(_04178_ ), .A2(_04092_ ), .A3(\CLINT.mtime [24] ), .ZN(_04217_ ) );
NAND2_X1 _11456_ ( .A1(_04216_ ), .A2(_04217_ ), .ZN(_04218_ ) );
MUX2_X1 _11457_ ( .A(\CLINT.c_axi_rdata [24] ), .B(_04218_ ), .S(_04181_ ), .Z(_00129_ ) );
NAND3_X1 _11458_ ( .A1(_04076_ ), .A2(_04102_ ), .A3(\CLINT.mtime [55] ), .ZN(_04219_ ) );
NAND3_X1 _11459_ ( .A1(_04100_ ), .A2(_04092_ ), .A3(\CLINT.mtime [23] ), .ZN(_04220_ ) );
NAND2_X1 _11460_ ( .A1(_04219_ ), .A2(_04220_ ), .ZN(_04221_ ) );
MUX2_X1 _11461_ ( .A(\CLINT.c_axi_rdata [23] ), .B(_04221_ ), .S(_04116_ ), .Z(_00130_ ) );
NAND3_X1 _11462_ ( .A1(_04076_ ), .A2(_04102_ ), .A3(\CLINT.mtime [54] ), .ZN(_04222_ ) );
NAND3_X1 _11463_ ( .A1(_04100_ ), .A2(_04092_ ), .A3(\CLINT.mtime [22] ), .ZN(_04223_ ) );
NAND2_X1 _11464_ ( .A1(_04222_ ), .A2(_04223_ ), .ZN(_04224_ ) );
MUX2_X1 _11465_ ( .A(\CLINT.c_axi_rdata [22] ), .B(_04224_ ), .S(_04116_ ), .Z(_00131_ ) );
NOR4_X1 _11466_ ( .A1(\EXU.dnpc_o [11] ), .A2(\EXU.dnpc_o [10] ), .A3(\EXU.dnpc_o [9] ), .A4(\EXU.dnpc_o [8] ), .ZN(_04225_ ) );
INV_X1 _11467_ ( .A(\EXU.dnpc_o [13] ), .ZN(_04226_ ) );
INV_X1 _11468_ ( .A(\EXU.dnpc_o [12] ), .ZN(_04227_ ) );
NOR2_X1 _11469_ ( .A1(\EXU.dnpc_o [15] ), .A2(\EXU.dnpc_o [14] ), .ZN(_04228_ ) );
NAND4_X1 _11470_ ( .A1(_04225_ ), .A2(_04226_ ), .A3(_04227_ ), .A4(_04228_ ), .ZN(_04229_ ) );
INV_X1 _11471_ ( .A(\EXU.dnpc_o [3] ), .ZN(_04230_ ) );
INV_X1 _11472_ ( .A(\EXU.dnpc_o [2] ), .ZN(_04231_ ) );
INV_X1 _11473_ ( .A(\EXU.dnpc_o [1] ), .ZN(_04232_ ) );
INV_X1 _11474_ ( .A(\EXU.dnpc_o [0] ), .ZN(_04233_ ) );
NAND4_X1 _11475_ ( .A1(_04230_ ), .A2(_04231_ ), .A3(_04232_ ), .A4(_04233_ ), .ZN(_04234_ ) );
INV_X1 _11476_ ( .A(\EXU.dnpc_o [7] ), .ZN(_04235_ ) );
INV_X1 _11477_ ( .A(\EXU.dnpc_o [6] ), .ZN(_04236_ ) );
INV_X1 _11478_ ( .A(\EXU.dnpc_o [5] ), .ZN(_04237_ ) );
INV_X1 _11479_ ( .A(\EXU.dnpc_o [4] ), .ZN(_04238_ ) );
NAND4_X1 _11480_ ( .A1(_04235_ ), .A2(_04236_ ), .A3(_04237_ ), .A4(_04238_ ), .ZN(_04239_ ) );
NOR3_X1 _11481_ ( .A1(_04229_ ), .A2(_04234_ ), .A3(_04239_ ), .ZN(_04240_ ) );
NOR2_X1 _11482_ ( .A1(\EXU.dnpc_o [19] ), .A2(\EXU.dnpc_o [18] ), .ZN(_04241_ ) );
INV_X1 _11483_ ( .A(\EXU.dnpc_o [17] ), .ZN(_04242_ ) );
INV_X1 _11484_ ( .A(\EXU.dnpc_o [16] ), .ZN(_04243_ ) );
NAND3_X1 _11485_ ( .A1(_04241_ ), .A2(_04242_ ), .A3(_04243_ ), .ZN(_04244_ ) );
OR4_X4 _11486_ ( .A1(\EXU.dnpc_o [31] ), .A2(\EXU.dnpc_o [30] ), .A3(\EXU.dnpc_o [29] ), .A4(\EXU.dnpc_o [28] ), .ZN(_04245_ ) );
INV_X1 _11487_ ( .A(\EXU.dnpc_o [27] ), .ZN(_04246_ ) );
INV_X1 _11488_ ( .A(\EXU.dnpc_o [26] ), .ZN(_04247_ ) );
INV_X1 _11489_ ( .A(\EXU.dnpc_o [25] ), .ZN(_04248_ ) );
INV_X1 _11490_ ( .A(\EXU.dnpc_o [24] ), .ZN(_04249_ ) );
NAND4_X1 _11491_ ( .A1(_04246_ ), .A2(_04247_ ), .A3(_04248_ ), .A4(_04249_ ), .ZN(_04250_ ) );
INV_X1 _11492_ ( .A(\EXU.dnpc_o [21] ), .ZN(_04251_ ) );
INV_X1 _11493_ ( .A(\EXU.dnpc_o [20] ), .ZN(_04252_ ) );
INV_X1 _11494_ ( .A(\EXU.dnpc_o [23] ), .ZN(_04253_ ) );
INV_X1 _11495_ ( .A(\EXU.dnpc_o [22] ), .ZN(_04254_ ) );
NAND4_X1 _11496_ ( .A1(_04251_ ), .A2(_04252_ ), .A3(_04253_ ), .A4(_04254_ ), .ZN(_04255_ ) );
NOR4_X1 _11497_ ( .A1(_04244_ ), .A2(_04245_ ), .A3(_04250_ ), .A4(_04255_ ), .ZN(_04256_ ) );
NAND2_X1 _11498_ ( .A1(_04240_ ), .A2(_04256_ ), .ZN(_04257_ ) );
NOR2_X1 _11499_ ( .A1(\EXU.pc_i [23] ), .A2(\EXU.pc_i [22] ), .ZN(_04258_ ) );
NOR2_X1 _11500_ ( .A1(\EXU.pc_i [21] ), .A2(\EXU.pc_i [20] ), .ZN(_04259_ ) );
AND2_X1 _11501_ ( .A1(_04258_ ), .A2(_04259_ ), .ZN(_04260_ ) );
INV_X1 _11502_ ( .A(\EXU.pc_i [19] ), .ZN(_04261_ ) );
INV_X1 _11503_ ( .A(\EXU.pc_i [18] ), .ZN(_04262_ ) );
NOR2_X1 _11504_ ( .A1(\EXU.pc_i [17] ), .A2(\EXU.pc_i [16] ), .ZN(_04263_ ) );
NAND4_X1 _11505_ ( .A1(_04260_ ), .A2(_04261_ ), .A3(_04262_ ), .A4(_04263_ ), .ZN(_04264_ ) );
NOR4_X1 _11506_ ( .A1(\EXU.pc_i [31] ), .A2(\EXU.pc_i [30] ), .A3(\EXU.pc_i [29] ), .A4(\EXU.pc_i [28] ), .ZN(_04265_ ) );
NOR4_X1 _11507_ ( .A1(\EXU.pc_i [27] ), .A2(\EXU.pc_i [26] ), .A3(\EXU.pc_i [25] ), .A4(\EXU.pc_i [24] ), .ZN(_04266_ ) );
NAND2_X1 _11508_ ( .A1(_04265_ ), .A2(_04266_ ), .ZN(_04267_ ) );
NOR2_X1 _11509_ ( .A1(_04264_ ), .A2(_04267_ ), .ZN(_04268_ ) );
OR4_X1 _11510_ ( .A1(\EXU.pc_i [3] ), .A2(\EXU.pc_i [2] ), .A3(\EXU.add_pc_4 [1] ), .A4(\EXU.add_pc_4 [0] ), .ZN(_04269_ ) );
INV_X1 _11511_ ( .A(\EXU.pc_i [7] ), .ZN(_04270_ ) );
INV_X1 _11512_ ( .A(\EXU.pc_i [6] ), .ZN(_04271_ ) );
INV_X1 _11513_ ( .A(\EXU.pc_i [5] ), .ZN(_04272_ ) );
INV_X1 _11514_ ( .A(\EXU.pc_i [4] ), .ZN(_04273_ ) );
NAND4_X1 _11515_ ( .A1(_04270_ ), .A2(_04271_ ), .A3(_04272_ ), .A4(_04273_ ), .ZN(_04274_ ) );
INV_X1 _11516_ ( .A(\EXU.pc_i [15] ), .ZN(_04275_ ) );
INV_X1 _11517_ ( .A(\EXU.pc_i [14] ), .ZN(_04276_ ) );
INV_X1 _11518_ ( .A(\EXU.pc_i [13] ), .ZN(_04277_ ) );
INV_X1 _11519_ ( .A(\EXU.pc_i [12] ), .ZN(_04278_ ) );
NAND4_X1 _11520_ ( .A1(_04275_ ), .A2(_04276_ ), .A3(_04277_ ), .A4(_04278_ ), .ZN(_04279_ ) );
INV_X1 _11521_ ( .A(\EXU.pc_i [11] ), .ZN(_04280_ ) );
INV_X1 _11522_ ( .A(\EXU.pc_i [10] ), .ZN(_04281_ ) );
INV_X1 _11523_ ( .A(\EXU.pc_i [9] ), .ZN(_04282_ ) );
INV_X1 _11524_ ( .A(\EXU.pc_i [8] ), .ZN(_04283_ ) );
NAND4_X1 _11525_ ( .A1(_04280_ ), .A2(_04281_ ), .A3(_04282_ ), .A4(_04283_ ), .ZN(_04284_ ) );
NOR4_X1 _11526_ ( .A1(_04269_ ), .A2(_04274_ ), .A3(_04279_ ), .A4(_04284_ ), .ZN(_04285_ ) );
NAND2_X1 _11527_ ( .A1(_04268_ ), .A2(_04285_ ), .ZN(_04286_ ) );
AND3_X2 _11528_ ( .A1(_04257_ ), .A2(CHazarden ), .A3(_04286_ ), .ZN(_04287_ ) );
XNOR2_X1 _11529_ ( .A(\EXU.dnpc_o [2] ), .B(\EXU.pc_i [2] ), .ZN(_04288_ ) );
XNOR2_X1 _11530_ ( .A(\EXU.dnpc_o [1] ), .B(\EXU.add_pc_4 [1] ), .ZN(_04289_ ) );
XNOR2_X1 _11531_ ( .A(\EXU.dnpc_o [10] ), .B(\EXU.pc_i [10] ), .ZN(_04290_ ) );
XNOR2_X1 _11532_ ( .A(\EXU.dnpc_o [5] ), .B(\EXU.pc_i [5] ), .ZN(_04291_ ) );
AND4_X1 _11533_ ( .A1(_04288_ ), .A2(_04289_ ), .A3(_04290_ ), .A4(_04291_ ), .ZN(_04292_ ) );
XNOR2_X1 _11534_ ( .A(\EXU.dnpc_o [19] ), .B(\EXU.pc_i [19] ), .ZN(_04293_ ) );
XNOR2_X1 _11535_ ( .A(\EXU.dnpc_o [18] ), .B(\EXU.pc_i [18] ), .ZN(_04294_ ) );
XNOR2_X1 _11536_ ( .A(\EXU.dnpc_o [28] ), .B(\EXU.pc_i [28] ), .ZN(_04295_ ) );
XNOR2_X1 _11537_ ( .A(\EXU.dnpc_o [24] ), .B(\EXU.pc_i [24] ), .ZN(_04296_ ) );
AND4_X1 _11538_ ( .A1(_04293_ ), .A2(_04294_ ), .A3(_04295_ ), .A4(_04296_ ), .ZN(_04297_ ) );
XNOR2_X1 _11539_ ( .A(\EXU.dnpc_o [9] ), .B(\EXU.pc_i [9] ), .ZN(_04298_ ) );
XNOR2_X1 _11540_ ( .A(\EXU.dnpc_o [6] ), .B(\EXU.pc_i [6] ), .ZN(_04299_ ) );
XNOR2_X1 _11541_ ( .A(\EXU.dnpc_o [20] ), .B(\EXU.pc_i [20] ), .ZN(_04300_ ) );
XNOR2_X1 _11542_ ( .A(\EXU.dnpc_o [16] ), .B(\EXU.pc_i [16] ), .ZN(_04301_ ) );
AND4_X1 _11543_ ( .A1(_04298_ ), .A2(_04299_ ), .A3(_04300_ ), .A4(_04301_ ), .ZN(_04302_ ) );
XNOR2_X1 _11544_ ( .A(\EXU.dnpc_o [30] ), .B(\EXU.pc_i [30] ), .ZN(_04303_ ) );
XNOR2_X1 _11545_ ( .A(\EXU.dnpc_o [27] ), .B(\EXU.pc_i [27] ), .ZN(_04304_ ) );
XNOR2_X1 _11546_ ( .A(\EXU.dnpc_o [7] ), .B(\EXU.pc_i [7] ), .ZN(_04305_ ) );
XNOR2_X1 _11547_ ( .A(\EXU.dnpc_o [26] ), .B(\EXU.pc_i [26] ), .ZN(_04306_ ) );
AND4_X1 _11548_ ( .A1(_04303_ ), .A2(_04304_ ), .A3(_04305_ ), .A4(_04306_ ), .ZN(_04307_ ) );
AND4_X1 _11549_ ( .A1(_04292_ ), .A2(_04297_ ), .A3(_04302_ ), .A4(_04307_ ), .ZN(_04308_ ) );
XNOR2_X1 _11550_ ( .A(\EXU.dnpc_o [14] ), .B(\EXU.pc_i [14] ), .ZN(_04309_ ) );
XNOR2_X1 _11551_ ( .A(\EXU.dnpc_o [8] ), .B(\EXU.pc_i [8] ), .ZN(_04310_ ) );
XNOR2_X1 _11552_ ( .A(\EXU.dnpc_o [3] ), .B(\EXU.pc_i [3] ), .ZN(_04311_ ) );
XNOR2_X1 _11553_ ( .A(\EXU.dnpc_o [4] ), .B(\EXU.pc_i [4] ), .ZN(_04312_ ) );
AND4_X1 _11554_ ( .A1(_04309_ ), .A2(_04310_ ), .A3(_04311_ ), .A4(_04312_ ), .ZN(_04313_ ) );
XNOR2_X1 _11555_ ( .A(\EXU.dnpc_o [23] ), .B(\EXU.pc_i [23] ), .ZN(_04314_ ) );
XNOR2_X1 _11556_ ( .A(\EXU.dnpc_o [22] ), .B(\EXU.pc_i [22] ), .ZN(_04315_ ) );
XNOR2_X1 _11557_ ( .A(\EXU.dnpc_o [21] ), .B(\EXU.pc_i [21] ), .ZN(_04316_ ) );
XNOR2_X1 _11558_ ( .A(\EXU.dnpc_o [17] ), .B(\EXU.pc_i [17] ), .ZN(_04317_ ) );
AND4_X1 _11559_ ( .A1(_04314_ ), .A2(_04315_ ), .A3(_04316_ ), .A4(_04317_ ), .ZN(_04318_ ) );
XNOR2_X1 _11560_ ( .A(\EXU.dnpc_o [12] ), .B(\EXU.pc_i [12] ), .ZN(_04319_ ) );
XNOR2_X1 _11561_ ( .A(\EXU.dnpc_o [15] ), .B(\EXU.pc_i [15] ), .ZN(_04320_ ) );
XNOR2_X1 _11562_ ( .A(\EXU.dnpc_o [13] ), .B(\EXU.pc_i [13] ), .ZN(_04321_ ) );
XNOR2_X1 _11563_ ( .A(\EXU.dnpc_o [0] ), .B(\EXU.add_pc_4 [0] ), .ZN(_04322_ ) );
AND4_X1 _11564_ ( .A1(_04319_ ), .A2(_04320_ ), .A3(_04321_ ), .A4(_04322_ ), .ZN(_04323_ ) );
XNOR2_X1 _11565_ ( .A(\EXU.dnpc_o [11] ), .B(\EXU.pc_i [11] ), .ZN(_04324_ ) );
XNOR2_X1 _11566_ ( .A(\EXU.dnpc_o [29] ), .B(\EXU.pc_i [29] ), .ZN(_04325_ ) );
XNOR2_X1 _11567_ ( .A(\EXU.dnpc_o [31] ), .B(\EXU.pc_i [31] ), .ZN(_04326_ ) );
XNOR2_X1 _11568_ ( .A(\EXU.dnpc_o [25] ), .B(\EXU.pc_i [25] ), .ZN(_04327_ ) );
AND4_X1 _11569_ ( .A1(_04324_ ), .A2(_04325_ ), .A3(_04326_ ), .A4(_04327_ ), .ZN(_04328_ ) );
AND4_X1 _11570_ ( .A1(_04313_ ), .A2(_04318_ ), .A3(_04323_ ), .A4(_04328_ ), .ZN(_04329_ ) );
NAND2_X1 _11571_ ( .A1(_04308_ ), .A2(_04329_ ), .ZN(_04330_ ) );
AND2_X1 _11572_ ( .A1(_04287_ ), .A2(_04330_ ), .ZN(_04331_ ) );
NOR2_X2 _11573_ ( .A1(_04331_ ), .A2(\LSU.ls_read_done_$_OR__B_Y_$_ORNOT__A_Y_$_ANDNOT__A_Y_$_OR__A_1_B ), .ZN(_04332_ ) );
INV_X16 _11574_ ( .A(\EXU.imm_i [0] ), .ZN(_04333_ ) );
AND2_X2 _11575_ ( .A1(_04333_ ), .A2(\EXU.imm_i [1] ), .ZN(_04334_ ) );
AND3_X1 _11576_ ( .A1(\EXU.imm_i [9] ), .A2(\EXU.imm_i [6] ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_04335_ ) );
AND2_X4 _11577_ ( .A1(_04334_ ), .A2(_04335_ ), .ZN(_04336_ ) );
AND2_X4 _11578_ ( .A1(\EXU.op_i [3] ), .A2(\EXU.op_i [2] ), .ZN(_04337_ ) );
NOR2_X4 _11579_ ( .A1(\EXU.op_i [1] ), .A2(\EXU.op_i [0] ), .ZN(_04338_ ) );
AND2_X4 _11580_ ( .A1(_04337_ ), .A2(_04338_ ), .ZN(_04339_ ) );
BUF_X8 _11581_ ( .A(_04339_ ), .Z(_04340_ ) );
AND3_X1 _11582_ ( .A1(_04336_ ), .A2(fanout_net_7 ), .A3(_04340_ ), .ZN(_04341_ ) );
INV_X1 _11583_ ( .A(_04341_ ), .ZN(_04342_ ) );
AND2_X4 _11584_ ( .A1(_04340_ ), .A2(fanout_net_7 ), .ZN(_04343_ ) );
INV_X1 _11585_ ( .A(\EXU.imm_i [11] ), .ZN(_04344_ ) );
NOR2_X2 _11586_ ( .A1(\EXU.imm_i [1] ), .A2(\EXU.imm_i [0] ), .ZN(_04345_ ) );
INV_X1 _11587_ ( .A(\EXU.imm_i [9] ), .ZN(_04346_ ) );
INV_X16 _11588_ ( .A(\EXU.imm_i [6] ), .ZN(_04347_ ) );
AND4_X2 _11589_ ( .A1(_04344_ ), .A2(_04345_ ), .A3(_04346_ ), .A4(_04347_ ), .ZN(_04348_ ) );
NOR2_X4 _11590_ ( .A1(_04333_ ), .A2(\EXU.imm_i [1] ), .ZN(_04349_ ) );
AND2_X2 _11591_ ( .A1(_04335_ ), .A2(_04349_ ), .ZN(_04350_ ) );
OAI21_X2 _11592_ ( .A(_04343_ ), .B1(_04348_ ), .B2(_04350_ ), .ZN(_04351_ ) );
AND3_X2 _11593_ ( .A1(_04347_ ), .A2(\EXU.imm_i [9] ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_04352_ ) );
AND2_X2 _11594_ ( .A1(_04352_ ), .A2(_04349_ ), .ZN(_04353_ ) );
NAND3_X1 _11595_ ( .A1(_04353_ ), .A2(fanout_net_7 ), .A3(_04340_ ), .ZN(_04354_ ) );
AND2_X2 _11596_ ( .A1(_04352_ ), .A2(_04345_ ), .ZN(_04355_ ) );
NAND2_X2 _11597_ ( .A1(_04343_ ), .A2(_04355_ ), .ZN(_04356_ ) );
NAND4_X2 _11598_ ( .A1(_04342_ ), .A2(_04351_ ), .A3(_04354_ ), .A4(_04356_ ), .ZN(_04357_ ) );
AND2_X4 _11599_ ( .A1(_04343_ ), .A2(_04348_ ), .ZN(_04358_ ) );
BUF_X8 _11600_ ( .A(_04358_ ), .Z(_04359_ ) );
INV_X4 _11601_ ( .A(_04359_ ), .ZN(_04360_ ) );
AND2_X4 _11602_ ( .A1(_04357_ ), .A2(_04360_ ), .ZN(_04361_ ) );
INV_X1 _11603_ ( .A(_04361_ ), .ZN(_04362_ ) );
INV_X1 _11604_ ( .A(\EXU.counter [1] ), .ZN(_04363_ ) );
XNOR2_X2 _11605_ ( .A(_04359_ ), .B(_04363_ ), .ZN(_04364_ ) );
INV_X1 _11606_ ( .A(_04364_ ), .ZN(_04365_ ) );
NAND3_X1 _11607_ ( .A1(_04362_ ), .A2(\EXU.counter [0] ), .A3(_04365_ ), .ZN(_04366_ ) );
INV_X1 _11608_ ( .A(\EXU.counter [0] ), .ZN(_04367_ ) );
OAI21_X2 _11609_ ( .A(_04364_ ), .B1(_04361_ ), .B2(_04367_ ), .ZN(_04368_ ) );
AND2_X2 _11610_ ( .A1(_04366_ ), .A2(_04368_ ), .ZN(_04369_ ) );
BUF_X8 _11611_ ( .A(_04369_ ), .Z(_04370_ ) );
BUF_X4 _11612_ ( .A(_04370_ ), .Z(_04371_ ) );
XOR2_X2 _11613_ ( .A(_04361_ ), .B(\EXU.counter_$_SDFFE_PP0N__Q_1_D [0] ), .Z(_04372_ ) );
INV_X4 _11614_ ( .A(_04372_ ), .ZN(_04373_ ) );
BUF_X2 _11615_ ( .A(_04373_ ), .Z(_04374_ ) );
AND3_X1 _11616_ ( .A1(_04371_ ), .A2(_04341_ ), .A3(_04374_ ), .ZN(_04375_ ) );
NOR2_X2 _11617_ ( .A1(_04373_ ), .A2(_04370_ ), .ZN(_04376_ ) );
BUF_X4 _11618_ ( .A(_04376_ ), .Z(_04377_ ) );
OAI21_X1 _11619_ ( .A(_04332_ ), .B1(_04375_ ), .B2(_04377_ ), .ZN(_04378_ ) );
INV_X1 _11620_ ( .A(\LSU.ls_axi_bready ), .ZN(_04379_ ) );
NOR2_X1 _11621_ ( .A1(_04056_ ), .A2(_04379_ ), .ZN(io_master_bready ) );
AND2_X1 _11622_ ( .A1(io_master_bready ), .A2(io_master_bvalid ), .ZN(_04380_ ) );
INV_X32 _11623_ ( .A(\EXU.op_i [2] ), .ZN(_04381_ ) );
AND3_X4 _11624_ ( .A1(_04338_ ), .A2(\EXU.op_i [3] ), .A3(_04381_ ), .ZN(_04382_ ) );
INV_X32 _11625_ ( .A(fanout_net_7 ), .ZN(_04383_ ) );
AND2_X4 _11626_ ( .A1(_04382_ ), .A2(_04383_ ), .ZN(_04384_ ) );
INV_X32 _11627_ ( .A(fanout_net_8 ), .ZN(_04385_ ) );
NOR3_X4 _11628_ ( .A1(_04385_ ), .A2(\EXU.op_i [1] ), .A3(\EXU.op_i [0] ), .ZN(_04386_ ) );
BUF_X8 _11629_ ( .A(_04386_ ), .Z(_04387_ ) );
NOR2_X4 _11630_ ( .A1(\EXU.op_i [3] ), .A2(\EXU.op_i [2] ), .ZN(_04388_ ) );
AND2_X4 _11631_ ( .A1(_04387_ ), .A2(_04388_ ), .ZN(_04389_ ) );
NOR2_X1 _11632_ ( .A1(_04384_ ), .A2(_04389_ ), .ZN(_04390_ ) );
NOR3_X1 _11633_ ( .A1(_04380_ ), .A2(_04390_ ), .A3(\LSU.ls_read_done ), .ZN(_04391_ ) );
NOR2_X4 _11634_ ( .A1(_04373_ ), .A2(_04391_ ), .ZN(_04392_ ) );
AND2_X2 _11635_ ( .A1(_04392_ ), .A2(_04370_ ), .ZN(_04393_ ) );
AND2_X2 _11636_ ( .A1(_04373_ ), .A2(_04370_ ), .ZN(_04394_ ) );
INV_X2 _11637_ ( .A(_04332_ ), .ZN(_04395_ ) );
NOR4_X1 _11638_ ( .A1(_04393_ ), .A2(_04394_ ), .A3(_04376_ ), .A4(_04395_ ), .ZN(_04396_ ) );
INV_X1 _11639_ ( .A(\LSU.ls_read_done_$_OR__B_Y_$_ORNOT__A_Y_$_ANDNOT__A_Y_$_OR__A_1_B ), .ZN(_04397_ ) );
AOI21_X1 _11640_ ( .A(_04397_ ), .B1(_04287_ ), .B2(_04330_ ), .ZN(_04398_ ) );
NOR2_X2 _11641_ ( .A1(_04396_ ), .A2(_04398_ ), .ZN(_04399_ ) );
BUF_X4 _11642_ ( .A(_04399_ ), .Z(_04400_ ) );
INV_X1 _11643_ ( .A(fanout_net_3 ), .ZN(_04401_ ) );
BUF_X4 _11644_ ( .A(_04401_ ), .Z(_04402_ ) );
OAI21_X1 _11645_ ( .A(_04378_ ), .B1(_04400_ ), .B2(_04402_ ), .ZN(_00199_ ) );
NAND3_X1 _11646_ ( .A1(_04374_ ), .A2(_04371_ ), .A3(_04332_ ), .ZN(_04403_ ) );
OR2_X1 _11647_ ( .A1(_04403_ ), .A2(_04354_ ), .ZN(_04404_ ) );
INV_X1 _11648_ ( .A(fanout_net_4 ), .ZN(_04405_ ) );
BUF_X4 _11649_ ( .A(_04405_ ), .Z(_04406_ ) );
OAI21_X1 _11650_ ( .A(_04404_ ), .B1(_04400_ ), .B2(_04406_ ), .ZN(_00200_ ) );
OR2_X1 _11651_ ( .A1(_04403_ ), .A2(_04356_ ), .ZN(_04407_ ) );
INV_X1 _11652_ ( .A(fanout_net_2 ), .ZN(_04408_ ) );
BUF_X4 _11653_ ( .A(_04408_ ), .Z(_04409_ ) );
OAI21_X1 _11654_ ( .A(_04407_ ), .B1(_04400_ ), .B2(_04409_ ), .ZN(_00201_ ) );
OR2_X1 _11655_ ( .A1(_04403_ ), .A2(_04351_ ), .ZN(_04410_ ) );
INV_X1 _11656_ ( .A(fanout_net_1 ), .ZN(_04411_ ) );
BUF_X4 _11657_ ( .A(_04411_ ), .Z(_04412_ ) );
OAI21_X1 _11658_ ( .A(_04410_ ), .B1(_04400_ ), .B2(_04412_ ), .ZN(_00202_ ) );
INV_X1 _11659_ ( .A(_04384_ ), .ZN(_04413_ ) );
INV_X2 _11660_ ( .A(_04389_ ), .ZN(_04414_ ) );
AND3_X4 _11661_ ( .A1(_04381_ ), .A2(fanout_net_7 ), .A3(\EXU.op_i [3] ), .ZN(_04415_ ) );
INV_X1 _11662_ ( .A(\EXU.op_i [0] ), .ZN(_04416_ ) );
NOR2_X2 _11663_ ( .A1(_04416_ ), .A2(\EXU.op_i [1] ), .ZN(_04417_ ) );
AND2_X1 _11664_ ( .A1(_04415_ ), .A2(_04417_ ), .ZN(_04418_ ) );
INV_X1 _11665_ ( .A(_04418_ ), .ZN(_04419_ ) );
NAND3_X4 _11666_ ( .A1(_04413_ ), .A2(_04414_ ), .A3(_04419_ ), .ZN(_04420_ ) );
AND2_X4 _11667_ ( .A1(_04339_ ), .A2(_04383_ ), .ZN(_04421_ ) );
BUF_X8 _11668_ ( .A(_04421_ ), .Z(_04422_ ) );
NOR2_X4 _11669_ ( .A1(_04381_ ), .A2(\EXU.op_i [3] ), .ZN(_04423_ ) );
AND2_X4 _11670_ ( .A1(_04386_ ), .A2(_04423_ ), .ZN(_04424_ ) );
NOR2_X4 _11671_ ( .A1(_04422_ ), .A2(_04424_ ), .ZN(_04425_ ) );
INV_X4 _11672_ ( .A(_04425_ ), .ZN(_04426_ ) );
BUF_X2 _11673_ ( .A(_04426_ ), .Z(_04427_ ) );
OAI21_X1 _11674_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_A ), .B1(_04420_ ), .B2(_04427_ ), .ZN(_04428_ ) );
NAND4_X1 _11675_ ( .A1(_04390_ ), .A2(_04425_ ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_B ), .A4(_04419_ ), .ZN(_04429_ ) );
AND2_X1 _11676_ ( .A1(_04428_ ), .A2(_04429_ ), .ZN(_04430_ ) );
BUF_X4 _11677_ ( .A(_04338_ ), .Z(_04431_ ) );
BUF_X2 _11678_ ( .A(_04431_ ), .Z(_04432_ ) );
NAND4_X1 _11679_ ( .A1(_04337_ ), .A2(_04432_ ), .A3(_04383_ ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04433_ ) );
BUF_X4 _11680_ ( .A(_04422_ ), .Z(_04434_ ) );
BUF_X4 _11681_ ( .A(_04434_ ), .Z(_04435_ ) );
BUF_X4 _11682_ ( .A(_04435_ ), .Z(_04436_ ) );
INV_X1 _11683_ ( .A(_04436_ ), .ZN(_04437_ ) );
NAND2_X1 _11684_ ( .A1(_04437_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_04438_ ) );
NAND3_X1 _11685_ ( .A1(_04430_ ), .A2(_04433_ ), .A3(_04438_ ), .ZN(_04439_ ) );
NOR2_X4 _11686_ ( .A1(_04420_ ), .A2(_04426_ ), .ZN(_04440_ ) );
BUF_X8 _11687_ ( .A(_04440_ ), .Z(_04441_ ) );
MUX2_X1 _11688_ ( .A(\EXU.r1_i [6] ), .B(\EXU.pc_i [6] ), .S(_04441_ ), .Z(_04442_ ) );
MUX2_X1 _11689_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_18_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_wdata_i_$_MUX__Y_17_A_$_ANDNOT__Y_B ), .S(_04434_ ), .Z(_04443_ ) );
XNOR2_X1 _11690_ ( .A(_04442_ ), .B(_04443_ ), .ZN(_04444_ ) );
MUX2_X1 _11691_ ( .A(\EXU.r1_i [4] ), .B(\EXU.pc_i [4] ), .S(_04441_ ), .Z(_04445_ ) );
INV_X1 _11692_ ( .A(_04445_ ), .ZN(_04446_ ) );
MUX2_X1 _11693_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_20_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_wdata_i_$_MUX__Y_19_A_$_ANDNOT__Y_B ), .S(_04422_ ), .Z(_04447_ ) );
OR2_X1 _11694_ ( .A1(_04446_ ), .A2(_04447_ ), .ZN(_04448_ ) );
MUX2_X1 _11695_ ( .A(\EXU.r1_i [1] ), .B(\EXU.add_pc_4 [1] ), .S(_04440_ ), .Z(_04449_ ) );
MUX2_X1 _11696_ ( .A(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_wdata_i_$_MUX__Y_22_A_$_ANDNOT__Y_B ), .S(_04422_ ), .Z(_04450_ ) );
INV_X2 _11697_ ( .A(_04450_ ), .ZN(_04451_ ) );
NAND2_X1 _11698_ ( .A1(_04449_ ), .A2(_04451_ ), .ZN(_04452_ ) );
XNOR2_X2 _11699_ ( .A(_04449_ ), .B(_04451_ ), .ZN(_04453_ ) );
MUX2_X1 _11700_ ( .A(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_A ), .B(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_B ), .S(_04440_ ), .Z(_04454_ ) );
MUX2_X1 _11701_ ( .A(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_wdata_i_$_MUX__Y_23_A_$_ANDNOT__Y_B ), .S(_04422_ ), .Z(_04455_ ) );
OR2_X4 _11702_ ( .A1(_04454_ ), .A2(_04455_ ), .ZN(_04456_ ) );
OAI21_X4 _11703_ ( .A(_04452_ ), .B1(_04453_ ), .B2(_04456_ ), .ZN(_04457_ ) );
INV_X1 _11704_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_B_$_MUX__Y_A ), .ZN(_04458_ ) );
NOR2_X2 _11705_ ( .A1(_04441_ ), .A2(_04458_ ), .ZN(_04459_ ) );
MUX2_X1 _11706_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_wdata_i_$_MUX__Y_21_A_$_ANDNOT__Y_B ), .S(_04422_ ), .Z(_04460_ ) );
AND4_X1 _11707_ ( .A1(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_B_$_MUX__Y_B ), .A2(_04390_ ), .A3(_04425_ ), .A4(_04419_ ), .ZN(_04461_ ) );
OR3_X4 _11708_ ( .A1(_04459_ ), .A2(_04460_ ), .A3(_04461_ ), .ZN(_04462_ ) );
OAI21_X1 _11709_ ( .A(_04460_ ), .B1(_04459_ ), .B2(_04461_ ), .ZN(_04463_ ) );
AND2_X4 _11710_ ( .A1(_04462_ ), .A2(_04463_ ), .ZN(_04464_ ) );
NAND2_X2 _11711_ ( .A1(_04457_ ), .A2(_04464_ ), .ZN(_04465_ ) );
AND2_X2 _11712_ ( .A1(_04465_ ), .A2(_04462_ ), .ZN(_04466_ ) );
INV_X2 _11713_ ( .A(_04466_ ), .ZN(_04467_ ) );
MUX2_X1 _11714_ ( .A(\EXU.r1_i [3] ), .B(\EXU.pc_i [3] ), .S(_04441_ ), .Z(_04468_ ) );
MUX2_X1 _11715_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_21_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_wdata_i_$_MUX__Y_20_A_$_ANDNOT__Y_B ), .S(_04422_ ), .Z(_04469_ ) );
XNOR2_X2 _11716_ ( .A(_04468_ ), .B(_04469_ ), .ZN(_04470_ ) );
NAND2_X2 _11717_ ( .A1(_04467_ ), .A2(_04470_ ), .ZN(_04471_ ) );
INV_X1 _11718_ ( .A(_04469_ ), .ZN(_04472_ ) );
NAND2_X1 _11719_ ( .A1(_04468_ ), .A2(_04472_ ), .ZN(_04473_ ) );
AND2_X4 _11720_ ( .A1(_04471_ ), .A2(_04473_ ), .ZN(_04474_ ) );
AND2_X1 _11721_ ( .A1(_04446_ ), .A2(_04447_ ), .ZN(_04475_ ) );
OAI21_X4 _11722_ ( .A(_04448_ ), .B1(_04474_ ), .B2(_04475_ ), .ZN(_04476_ ) );
MUX2_X1 _11723_ ( .A(\EXU.r1_i [5] ), .B(\EXU.pc_i [5] ), .S(_04441_ ), .Z(_04477_ ) );
MUX2_X1 _11724_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_19_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_wdata_i_$_MUX__Y_18_A_$_ANDNOT__Y_B ), .S(_04434_ ), .Z(_04478_ ) );
XNOR2_X1 _11725_ ( .A(_04477_ ), .B(_04478_ ), .ZN(_04479_ ) );
AND2_X4 _11726_ ( .A1(_04476_ ), .A2(_04479_ ), .ZN(_04480_ ) );
INV_X1 _11727_ ( .A(_04478_ ), .ZN(_04481_ ) );
AND2_X1 _11728_ ( .A1(_04477_ ), .A2(_04481_ ), .ZN(_04482_ ) );
OAI21_X4 _11729_ ( .A(_04444_ ), .B1(_04480_ ), .B2(_04482_ ), .ZN(_04483_ ) );
INV_X1 _11730_ ( .A(_04442_ ), .ZN(_04484_ ) );
OAI21_X4 _11731_ ( .A(_04483_ ), .B1(_04443_ ), .B2(_04484_ ), .ZN(_04485_ ) );
BUF_X8 _11732_ ( .A(_04441_ ), .Z(_04486_ ) );
MUX2_X1 _11733_ ( .A(\EXU.r1_i [7] ), .B(\EXU.pc_i [7] ), .S(_04486_ ), .Z(_04487_ ) );
MUX2_X1 _11734_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_17_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_wdata_i_$_MUX__Y_16_A_$_ANDNOT__Y_B ), .S(_04435_ ), .Z(_04488_ ) );
XNOR2_X1 _11735_ ( .A(_04487_ ), .B(_04488_ ), .ZN(_04489_ ) );
NAND2_X4 _11736_ ( .A1(_04485_ ), .A2(_04489_ ), .ZN(_04490_ ) );
INV_X1 _11737_ ( .A(_04488_ ), .ZN(_04491_ ) );
NAND2_X1 _11738_ ( .A1(_04487_ ), .A2(_04491_ ), .ZN(_04492_ ) );
NAND2_X4 _11739_ ( .A1(_04490_ ), .A2(_04492_ ), .ZN(_04493_ ) );
MUX2_X1 _11740_ ( .A(\EXU.r1_i [14] ), .B(\EXU.pc_i [14] ), .S(_04441_ ), .Z(_04494_ ) );
INV_X1 _11741_ ( .A(_04494_ ), .ZN(_04495_ ) );
MUX2_X1 _11742_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_11_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_11_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04434_ ), .Z(_04496_ ) );
NOR2_X1 _11743_ ( .A1(_04495_ ), .A2(_04496_ ), .ZN(_04497_ ) );
INV_X1 _11744_ ( .A(_04497_ ), .ZN(_04498_ ) );
MUX2_X1 _11745_ ( .A(\EXU.r1_i [15] ), .B(\EXU.pc_i [15] ), .S(_04441_ ), .Z(_04499_ ) );
MUX2_X1 _11746_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_10_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_10_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04434_ ), .Z(_04500_ ) );
XNOR2_X2 _11747_ ( .A(_04499_ ), .B(_04500_ ), .ZN(_04501_ ) );
NAND2_X1 _11748_ ( .A1(_04495_ ), .A2(_04496_ ), .ZN(_04502_ ) );
AND3_X1 _11749_ ( .A1(_04498_ ), .A2(_04501_ ), .A3(_04502_ ), .ZN(_04503_ ) );
MUX2_X1 _11750_ ( .A(\EXU.r1_i [13] ), .B(\EXU.pc_i [13] ), .S(_04441_ ), .Z(_04504_ ) );
MUX2_X1 _11751_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04434_ ), .Z(_04505_ ) );
XNOR2_X1 _11752_ ( .A(_04504_ ), .B(_04505_ ), .ZN(_04506_ ) );
MUX2_X1 _11753_ ( .A(\EXU.r1_i [12] ), .B(\EXU.pc_i [12] ), .S(_04441_ ), .Z(_04507_ ) );
MUX2_X1 _11754_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ), .S(_04434_ ), .Z(_04508_ ) );
XNOR2_X1 _11755_ ( .A(_04507_ ), .B(_04508_ ), .ZN(_04509_ ) );
AND2_X1 _11756_ ( .A1(_04506_ ), .A2(_04509_ ), .ZN(_04510_ ) );
MUX2_X1 _11757_ ( .A(\EXU.r1_i [11] ), .B(\EXU.pc_i [11] ), .S(_04486_ ), .Z(_04511_ ) );
MUX2_X1 _11758_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04434_ ), .Z(_04512_ ) );
XNOR2_X1 _11759_ ( .A(_04511_ ), .B(_04512_ ), .ZN(_04513_ ) );
INV_X1 _11760_ ( .A(_04513_ ), .ZN(_04514_ ) );
MUX2_X1 _11761_ ( .A(\EXU.r1_i [10] ), .B(\EXU.pc_i [10] ), .S(_04486_ ), .Z(_04515_ ) );
MUX2_X1 _11762_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_14_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_14_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04435_ ), .Z(_04516_ ) );
XOR2_X1 _11763_ ( .A(_04515_ ), .B(_04516_ ), .Z(_04517_ ) );
NOR2_X1 _11764_ ( .A1(_04514_ ), .A2(_04517_ ), .ZN(_04518_ ) );
MUX2_X1 _11765_ ( .A(\EXU.r1_i [9] ), .B(\EXU.pc_i [9] ), .S(_04486_ ), .Z(_04519_ ) );
MUX2_X1 _11766_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_15_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_15_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04434_ ), .Z(_04520_ ) );
XNOR2_X2 _11767_ ( .A(_04519_ ), .B(_04520_ ), .ZN(_04521_ ) );
MUX2_X1 _11768_ ( .A(\EXU.r1_i [8] ), .B(\EXU.pc_i [8] ), .S(_04486_ ), .Z(_04522_ ) );
MUX2_X1 _11769_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_16_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_16_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04435_ ), .Z(_04523_ ) );
XNOR2_X1 _11770_ ( .A(_04522_ ), .B(_04523_ ), .ZN(_04524_ ) );
AND2_X1 _11771_ ( .A1(_04521_ ), .A2(_04524_ ), .ZN(_04525_ ) );
AND2_X1 _11772_ ( .A1(_04518_ ), .A2(_04525_ ), .ZN(_04526_ ) );
NAND4_X4 _11773_ ( .A1(_04493_ ), .A2(_04503_ ), .A3(_04510_ ), .A4(_04526_ ), .ZN(_04527_ ) );
NAND2_X1 _11774_ ( .A1(_04503_ ), .A2(_04510_ ), .ZN(_04528_ ) );
INV_X1 _11775_ ( .A(_04523_ ), .ZN(_04529_ ) );
NAND3_X1 _11776_ ( .A1(_04521_ ), .A2(_04529_ ), .A3(_04522_ ), .ZN(_04530_ ) );
INV_X1 _11777_ ( .A(_04519_ ), .ZN(_04531_ ) );
OAI21_X1 _11778_ ( .A(_04530_ ), .B1(_04520_ ), .B2(_04531_ ), .ZN(_04532_ ) );
NAND2_X1 _11779_ ( .A1(_04532_ ), .A2(_04518_ ), .ZN(_04533_ ) );
INV_X1 _11780_ ( .A(_04515_ ), .ZN(_04534_ ) );
NOR2_X1 _11781_ ( .A1(_04534_ ), .A2(_04516_ ), .ZN(_04535_ ) );
AND2_X2 _11782_ ( .A1(_04513_ ), .A2(_04535_ ), .ZN(_04536_ ) );
INV_X1 _11783_ ( .A(_04512_ ), .ZN(_04537_ ) );
AOI21_X1 _11784_ ( .A(_04536_ ), .B1(_04537_ ), .B2(_04511_ ), .ZN(_04538_ ) );
AOI21_X1 _11785_ ( .A(_04528_ ), .B1(_04533_ ), .B2(_04538_ ), .ZN(_04539_ ) );
INV_X1 _11786_ ( .A(_04500_ ), .ZN(_04540_ ) );
AND2_X1 _11787_ ( .A1(_04499_ ), .A2(_04540_ ), .ZN(_04541_ ) );
INV_X1 _11788_ ( .A(_04508_ ), .ZN(_04542_ ) );
NAND3_X1 _11789_ ( .A1(_04506_ ), .A2(_04542_ ), .A3(_04507_ ), .ZN(_04543_ ) );
INV_X1 _11790_ ( .A(_04504_ ), .ZN(_04544_ ) );
OAI21_X1 _11791_ ( .A(_04543_ ), .B1(_04505_ ), .B2(_04544_ ), .ZN(_04545_ ) );
AND2_X1 _11792_ ( .A1(_04545_ ), .A2(_04503_ ), .ZN(_04546_ ) );
AND2_X1 _11793_ ( .A1(_04501_ ), .A2(_04497_ ), .ZN(_04547_ ) );
NOR4_X4 _11794_ ( .A1(_04539_ ), .A2(_04541_ ), .A3(_04546_ ), .A4(_04547_ ), .ZN(_04548_ ) );
AND2_X4 _11795_ ( .A1(_04527_ ), .A2(_04548_ ), .ZN(_04549_ ) );
INV_X4 _11796_ ( .A(_04549_ ), .ZN(_04550_ ) );
MUX2_X1 _11797_ ( .A(\EXU.r1_i [22] ), .B(\EXU.pc_i [22] ), .S(_04486_ ), .Z(_04551_ ) );
MUX2_X1 _11798_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_5_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_5_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04435_ ), .Z(_04552_ ) );
XOR2_X1 _11799_ ( .A(_04551_ ), .B(_04552_ ), .Z(_04553_ ) );
BUF_X4 _11800_ ( .A(_04486_ ), .Z(_04554_ ) );
MUX2_X1 _11801_ ( .A(\EXU.r1_i [23] ), .B(\EXU.pc_i [23] ), .S(_04554_ ), .Z(_04555_ ) );
MUX2_X1 _11802_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_4_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_4_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04435_ ), .Z(_04556_ ) );
INV_X1 _11803_ ( .A(_04556_ ), .ZN(_04557_ ) );
AND2_X1 _11804_ ( .A1(_04555_ ), .A2(_04557_ ), .ZN(_04558_ ) );
NOR2_X1 _11805_ ( .A1(_04555_ ), .A2(_04557_ ), .ZN(_04559_ ) );
NOR3_X1 _11806_ ( .A1(_04553_ ), .A2(_04558_ ), .A3(_04559_ ), .ZN(_04560_ ) );
MUX2_X1 _11807_ ( .A(\EXU.r1_i [21] ), .B(\EXU.pc_i [21] ), .S(_04486_ ), .Z(_04561_ ) );
MUX2_X1 _11808_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04435_ ), .Z(_04562_ ) );
XNOR2_X1 _11809_ ( .A(_04561_ ), .B(_04562_ ), .ZN(_04563_ ) );
MUX2_X1 _11810_ ( .A(\EXU.r1_i [20] ), .B(\EXU.pc_i [20] ), .S(_04486_ ), .Z(_04564_ ) );
MUX2_X1 _11811_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ), .S(_04435_ ), .Z(_04565_ ) );
XNOR2_X1 _11812_ ( .A(_04564_ ), .B(_04565_ ), .ZN(_04566_ ) );
AND2_X1 _11813_ ( .A1(_04563_ ), .A2(_04566_ ), .ZN(_04567_ ) );
MUX2_X1 _11814_ ( .A(\EXU.r1_i [19] ), .B(\EXU.pc_i [19] ), .S(_04486_ ), .Z(_04568_ ) );
MUX2_X1 _11815_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_7_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_7_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04435_ ), .Z(_04569_ ) );
XNOR2_X1 _11816_ ( .A(_04568_ ), .B(_04569_ ), .ZN(_04570_ ) );
INV_X1 _11817_ ( .A(_04570_ ), .ZN(_04571_ ) );
MUX2_X1 _11818_ ( .A(\EXU.r1_i [18] ), .B(\EXU.pc_i [18] ), .S(_04554_ ), .Z(_04572_ ) );
MUX2_X1 _11819_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_8_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_8_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04436_ ), .Z(_04573_ ) );
XOR2_X1 _11820_ ( .A(_04572_ ), .B(_04573_ ), .Z(_04574_ ) );
NOR2_X1 _11821_ ( .A1(_04571_ ), .A2(_04574_ ), .ZN(_04575_ ) );
MUX2_X1 _11822_ ( .A(\EXU.r1_i [17] ), .B(\EXU.pc_i [17] ), .S(_04554_ ), .Z(_04576_ ) );
MUX2_X1 _11823_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04435_ ), .Z(_04577_ ) );
XNOR2_X1 _11824_ ( .A(_04576_ ), .B(_04577_ ), .ZN(_04578_ ) );
MUX2_X1 _11825_ ( .A(\EXU.r1_i [16] ), .B(\EXU.pc_i [16] ), .S(_04554_ ), .Z(_04579_ ) );
MUX2_X1 _11826_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ), .S(_04436_ ), .Z(_04580_ ) );
XNOR2_X1 _11827_ ( .A(_04579_ ), .B(_04580_ ), .ZN(_04581_ ) );
AND2_X1 _11828_ ( .A1(_04578_ ), .A2(_04581_ ), .ZN(_04582_ ) );
AND2_X1 _11829_ ( .A1(_04575_ ), .A2(_04582_ ), .ZN(_04583_ ) );
NAND4_X4 _11830_ ( .A1(_04550_ ), .A2(_04560_ ), .A3(_04567_ ), .A4(_04583_ ), .ZN(_04584_ ) );
NAND2_X1 _11831_ ( .A1(_04560_ ), .A2(_04567_ ), .ZN(_04585_ ) );
INV_X1 _11832_ ( .A(_04580_ ), .ZN(_04586_ ) );
NAND3_X1 _11833_ ( .A1(_04578_ ), .A2(_04586_ ), .A3(_04579_ ), .ZN(_04587_ ) );
INV_X1 _11834_ ( .A(_04576_ ), .ZN(_04588_ ) );
OAI21_X1 _11835_ ( .A(_04587_ ), .B1(_04577_ ), .B2(_04588_ ), .ZN(_04589_ ) );
NAND2_X1 _11836_ ( .A1(_04589_ ), .A2(_04575_ ), .ZN(_04590_ ) );
INV_X1 _11837_ ( .A(_04572_ ), .ZN(_04591_ ) );
NOR2_X1 _11838_ ( .A1(_04591_ ), .A2(_04573_ ), .ZN(_04592_ ) );
AND2_X1 _11839_ ( .A1(_04570_ ), .A2(_04592_ ), .ZN(_04593_ ) );
INV_X1 _11840_ ( .A(_04569_ ), .ZN(_04594_ ) );
AOI21_X1 _11841_ ( .A(_04593_ ), .B1(_04594_ ), .B2(_04568_ ), .ZN(_04595_ ) );
AOI21_X1 _11842_ ( .A(_04585_ ), .B1(_04590_ ), .B2(_04595_ ), .ZN(_04596_ ) );
INV_X1 _11843_ ( .A(_04565_ ), .ZN(_04597_ ) );
NAND3_X1 _11844_ ( .A1(_04563_ ), .A2(_04597_ ), .A3(_04564_ ), .ZN(_04598_ ) );
INV_X1 _11845_ ( .A(_04561_ ), .ZN(_04599_ ) );
OAI21_X1 _11846_ ( .A(_04598_ ), .B1(_04562_ ), .B2(_04599_ ), .ZN(_04600_ ) );
AND2_X1 _11847_ ( .A1(_04600_ ), .A2(_04560_ ), .ZN(_04601_ ) );
INV_X1 _11848_ ( .A(_04551_ ), .ZN(_04602_ ) );
NOR4_X1 _11849_ ( .A1(_04558_ ), .A2(_04559_ ), .A3(_04552_ ), .A4(_04602_ ), .ZN(_04603_ ) );
NOR4_X1 _11850_ ( .A1(_04596_ ), .A2(_04558_ ), .A3(_04601_ ), .A4(_04603_ ), .ZN(_04604_ ) );
AND2_X4 _11851_ ( .A1(_04584_ ), .A2(_04604_ ), .ZN(_04605_ ) );
INV_X4 _11852_ ( .A(_04605_ ), .ZN(_04606_ ) );
MUX2_X1 _11853_ ( .A(\EXU.r1_i [26] ), .B(\EXU.pc_i [26] ), .S(_04554_ ), .Z(_04607_ ) );
MUX2_X1 _11854_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .S(_04436_ ), .Z(_04608_ ) );
INV_X1 _11855_ ( .A(_04608_ ), .ZN(_04609_ ) );
XNOR2_X1 _11856_ ( .A(_04607_ ), .B(_04609_ ), .ZN(_04610_ ) );
MUX2_X1 _11857_ ( .A(\EXU.r1_i [27] ), .B(\EXU.pc_i [27] ), .S(_04554_ ), .Z(_04611_ ) );
AND4_X1 _11858_ ( .A1(_04383_ ), .A2(_04337_ ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_2_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .A4(_04432_ ), .ZN(_04612_ ) );
AOI21_X1 _11859_ ( .A(_04612_ ), .B1(_04437_ ), .B2(\LSU.ls_addr_i_$_ANDNOT__Y_2_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_04613_ ) );
XNOR2_X1 _11860_ ( .A(_04611_ ), .B(_04613_ ), .ZN(_04614_ ) );
NOR2_X1 _11861_ ( .A1(_04610_ ), .A2(_04614_ ), .ZN(_04615_ ) );
MUX2_X1 _11862_ ( .A(\EXU.r1_i [25] ), .B(\EXU.pc_i [25] ), .S(_04554_ ), .Z(_04616_ ) );
MUX2_X1 _11863_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A ), .S(_04436_ ), .Z(_04617_ ) );
XNOR2_X1 _11864_ ( .A(_04616_ ), .B(_04617_ ), .ZN(_04618_ ) );
MUX2_X1 _11865_ ( .A(\EXU.r1_i [24] ), .B(\EXU.pc_i [24] ), .S(_04554_ ), .Z(_04619_ ) );
MUX2_X1 _11866_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_A ), .S(_04436_ ), .Z(_04620_ ) );
XNOR2_X1 _11867_ ( .A(_04619_ ), .B(_04620_ ), .ZN(_04621_ ) );
AND2_X1 _11868_ ( .A1(_04618_ ), .A2(_04621_ ), .ZN(_04622_ ) );
NAND3_X4 _11869_ ( .A1(_04606_ ), .A2(_04615_ ), .A3(_04622_ ), .ZN(_04623_ ) );
NAND2_X1 _11870_ ( .A1(_04607_ ), .A2(_04609_ ), .ZN(_04624_ ) );
NOR2_X1 _11871_ ( .A1(_04614_ ), .A2(_04624_ ), .ZN(_04625_ ) );
INV_X1 _11872_ ( .A(_04620_ ), .ZN(_04626_ ) );
NAND3_X1 _11873_ ( .A1(_04618_ ), .A2(_04626_ ), .A3(_04619_ ), .ZN(_04627_ ) );
INV_X1 _11874_ ( .A(_04616_ ), .ZN(_04628_ ) );
OAI21_X1 _11875_ ( .A(_04627_ ), .B1(_04617_ ), .B2(_04628_ ), .ZN(_04629_ ) );
AOI221_X4 _11876_ ( .A(_04625_ ), .B1(_04613_ ), .B2(_04611_ ), .C1(_04629_ ), .C2(_04615_ ), .ZN(_04630_ ) );
AND2_X4 _11877_ ( .A1(_04623_ ), .A2(_04630_ ), .ZN(_04631_ ) );
INV_X4 _11878_ ( .A(_04631_ ), .ZN(_04632_ ) );
MUX2_X1 _11879_ ( .A(\EXU.r1_i [29] ), .B(\EXU.pc_i [29] ), .S(_04554_ ), .Z(_04633_ ) );
MUX2_X1 _11880_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ), .S(_04436_ ), .Z(_04634_ ) );
XNOR2_X1 _11881_ ( .A(_04633_ ), .B(_04634_ ), .ZN(_04635_ ) );
OAI21_X1 _11882_ ( .A(\EXU.r1_i [28] ), .B1(_04420_ ), .B2(_04427_ ), .ZN(_04636_ ) );
MUX2_X1 _11883_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_A ), .S(_04436_ ), .Z(_04637_ ) );
NAND4_X1 _11884_ ( .A1(_04390_ ), .A2(_04425_ ), .A3(\EXU.pc_i [28] ), .A4(_04419_ ), .ZN(_04638_ ) );
AND3_X1 _11885_ ( .A1(_04636_ ), .A2(_04637_ ), .A3(_04638_ ), .ZN(_04639_ ) );
AOI21_X1 _11886_ ( .A(_04637_ ), .B1(_04636_ ), .B2(_04638_ ), .ZN(_04640_ ) );
NOR2_X1 _11887_ ( .A1(_04639_ ), .A2(_04640_ ), .ZN(_04641_ ) );
AND3_X4 _11888_ ( .A1(_04632_ ), .A2(_04635_ ), .A3(_04641_ ), .ZN(_04642_ ) );
INV_X1 _11889_ ( .A(_04634_ ), .ZN(_04643_ ) );
AND2_X1 _11890_ ( .A1(_04633_ ), .A2(_04643_ ), .ZN(_04644_ ) );
AND2_X1 _11891_ ( .A1(_04635_ ), .A2(_04640_ ), .ZN(_04645_ ) );
NOR3_X4 _11892_ ( .A1(_04642_ ), .A2(_04644_ ), .A3(_04645_ ), .ZN(_04646_ ) );
NAND2_X1 _11893_ ( .A1(_04438_ ), .A2(_04433_ ), .ZN(_04647_ ) );
XOR2_X1 _11894_ ( .A(_04430_ ), .B(_04647_ ), .Z(_04648_ ) );
OAI21_X2 _11895_ ( .A(_04439_ ), .B1(_04646_ ), .B2(_04648_ ), .ZN(_04649_ ) );
MUX2_X1 _11896_ ( .A(\EXU.r1_i [31] ), .B(\EXU.pc_i [31] ), .S(_04554_ ), .Z(_04650_ ) );
MUX2_X1 _11897_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A ), .S(_04436_ ), .Z(_04651_ ) );
XNOR2_X1 _11898_ ( .A(_04650_ ), .B(_04651_ ), .ZN(_04652_ ) );
XOR2_X2 _11899_ ( .A(_04649_ ), .B(_04652_ ), .Z(_04653_ ) );
XNOR2_X1 _11900_ ( .A(\EXU.r1_i [1] ), .B(\EXU.r2_i [1] ), .ZN(_04654_ ) );
INV_X1 _11901_ ( .A(_04654_ ), .ZN(_04655_ ) );
XNOR2_X1 _11902_ ( .A(\EXU.r1_i [30] ), .B(\EXU.r2_i [30] ), .ZN(_04656_ ) );
INV_X1 _11903_ ( .A(_04656_ ), .ZN(_04657_ ) );
XOR2_X1 _11904_ ( .A(\EXU.r1_i [0] ), .B(\EXU.r2_i [0] ), .Z(_04658_ ) );
XOR2_X1 _11905_ ( .A(\EXU.r1_i [31] ), .B(\EXU.r2_i [31] ), .Z(_04659_ ) );
NOR4_X1 _11906_ ( .A1(_04655_ ), .A2(_04657_ ), .A3(_04658_ ), .A4(_04659_ ), .ZN(_04660_ ) );
XNOR2_X1 _11907_ ( .A(\EXU.r1_i [3] ), .B(\EXU.r2_i [3] ), .ZN(_04661_ ) );
XNOR2_X1 _11908_ ( .A(\EXU.r1_i [2] ), .B(\EXU.r2_i [2] ), .ZN(_04662_ ) );
XNOR2_X1 _11909_ ( .A(\EXU.r1_i [29] ), .B(\EXU.r2_i [29] ), .ZN(_04663_ ) );
XNOR2_X1 _11910_ ( .A(\EXU.r1_i [28] ), .B(\EXU.r2_i [28] ), .ZN(_04664_ ) );
AND4_X1 _11911_ ( .A1(_04661_ ), .A2(_04662_ ), .A3(_04663_ ), .A4(_04664_ ), .ZN(_04665_ ) );
AND2_X1 _11912_ ( .A1(_04660_ ), .A2(_04665_ ), .ZN(_04666_ ) );
XNOR2_X1 _11913_ ( .A(\EXU.r1_i [7] ), .B(\EXU.r2_i [7] ), .ZN(_04667_ ) );
XNOR2_X1 _11914_ ( .A(\EXU.r1_i [6] ), .B(\EXU.r2_i [6] ), .ZN(_04668_ ) );
AND2_X1 _11915_ ( .A1(_04667_ ), .A2(_04668_ ), .ZN(_04669_ ) );
XNOR2_X1 _11916_ ( .A(\EXU.r1_i [5] ), .B(\EXU.r2_i [5] ), .ZN(_04670_ ) );
XNOR2_X1 _11917_ ( .A(\EXU.r1_i [4] ), .B(\EXU.r2_i [4] ), .ZN(_04671_ ) );
AND2_X1 _11918_ ( .A1(_04670_ ), .A2(_04671_ ), .ZN(_04672_ ) );
XNOR2_X1 _11919_ ( .A(\EXU.r1_i [25] ), .B(\EXU.r2_i [25] ), .ZN(_04673_ ) );
XNOR2_X1 _11920_ ( .A(\EXU.r1_i [24] ), .B(\EXU.r2_i [24] ), .ZN(_04674_ ) );
AND2_X1 _11921_ ( .A1(_04673_ ), .A2(_04674_ ), .ZN(_04675_ ) );
XNOR2_X1 _11922_ ( .A(\EXU.r1_i [27] ), .B(\EXU.r2_i [27] ), .ZN(_04676_ ) );
XNOR2_X1 _11923_ ( .A(\EXU.r1_i [26] ), .B(\EXU.r2_i [26] ), .ZN(_04677_ ) );
AND3_X1 _11924_ ( .A1(_04675_ ), .A2(_04676_ ), .A3(_04677_ ), .ZN(_04678_ ) );
AND4_X1 _11925_ ( .A1(_04666_ ), .A2(_04669_ ), .A3(_04672_ ), .A4(_04678_ ), .ZN(_04679_ ) );
XNOR2_X1 _11926_ ( .A(\EXU.r1_i [15] ), .B(\EXU.r2_i [15] ), .ZN(_04680_ ) );
XNOR2_X1 _11927_ ( .A(\EXU.r1_i [14] ), .B(\EXU.r2_i [14] ), .ZN(_04681_ ) );
NAND2_X1 _11928_ ( .A1(_04680_ ), .A2(_04681_ ), .ZN(_04682_ ) );
XNOR2_X1 _11929_ ( .A(\EXU.r1_i [13] ), .B(\EXU.r2_i [13] ), .ZN(_04683_ ) );
INV_X1 _11930_ ( .A(_04683_ ), .ZN(_04684_ ) );
XNOR2_X1 _11931_ ( .A(\EXU.r1_i [12] ), .B(\EXU.r2_i [12] ), .ZN(_04685_ ) );
INV_X1 _11932_ ( .A(_04685_ ), .ZN(_04686_ ) );
NOR3_X1 _11933_ ( .A1(_04682_ ), .A2(_04684_ ), .A3(_04686_ ), .ZN(_04687_ ) );
XNOR2_X1 _11934_ ( .A(\EXU.r1_i [21] ), .B(\EXU.r2_i [21] ), .ZN(_04688_ ) );
XNOR2_X1 _11935_ ( .A(\EXU.r1_i [20] ), .B(\EXU.r2_i [20] ), .ZN(_04689_ ) );
AND2_X1 _11936_ ( .A1(_04688_ ), .A2(_04689_ ), .ZN(_04690_ ) );
XNOR2_X1 _11937_ ( .A(\EXU.r1_i [23] ), .B(\EXU.r2_i [23] ), .ZN(_04691_ ) );
XNOR2_X1 _11938_ ( .A(\EXU.r1_i [22] ), .B(\EXU.r2_i [22] ), .ZN(_04692_ ) );
AND3_X1 _11939_ ( .A1(_04690_ ), .A2(_04691_ ), .A3(_04692_ ), .ZN(_04693_ ) );
XNOR2_X1 _11940_ ( .A(\EXU.r1_i [11] ), .B(\EXU.r2_i [11] ), .ZN(_04694_ ) );
XNOR2_X1 _11941_ ( .A(\EXU.r1_i [10] ), .B(\EXU.r2_i [10] ), .ZN(_04695_ ) );
AND2_X1 _11942_ ( .A1(_04694_ ), .A2(_04695_ ), .ZN(_04696_ ) );
XNOR2_X1 _11943_ ( .A(\EXU.r1_i [9] ), .B(\EXU.r2_i [9] ), .ZN(_04697_ ) );
XNOR2_X1 _11944_ ( .A(\EXU.r1_i [8] ), .B(\EXU.r2_i [8] ), .ZN(_04698_ ) );
AND2_X1 _11945_ ( .A1(_04697_ ), .A2(_04698_ ), .ZN(_04699_ ) );
AND2_X1 _11946_ ( .A1(_04696_ ), .A2(_04699_ ), .ZN(_04700_ ) );
XNOR2_X1 _11947_ ( .A(\EXU.r1_i [19] ), .B(\EXU.r2_i [19] ), .ZN(_04701_ ) );
XNOR2_X1 _11948_ ( .A(\EXU.r1_i [18] ), .B(\EXU.r2_i [18] ), .ZN(_04702_ ) );
AND2_X1 _11949_ ( .A1(_04701_ ), .A2(_04702_ ), .ZN(_04703_ ) );
XNOR2_X1 _11950_ ( .A(\EXU.r1_i [17] ), .B(\EXU.r2_i [17] ), .ZN(_04704_ ) );
XNOR2_X1 _11951_ ( .A(\EXU.r1_i [16] ), .B(\EXU.r2_i [16] ), .ZN(_04705_ ) );
AND2_X1 _11952_ ( .A1(_04704_ ), .A2(_04705_ ), .ZN(_04706_ ) );
AND2_X1 _11953_ ( .A1(_04703_ ), .A2(_04706_ ), .ZN(_04707_ ) );
AND4_X1 _11954_ ( .A1(_04687_ ), .A2(_04693_ ), .A3(_04700_ ), .A4(_04707_ ), .ZN(_04708_ ) );
NOR2_X1 _11955_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .ZN(_04709_ ) );
INV_X1 _11956_ ( .A(\EXU.funct3_i [2] ), .ZN(_04710_ ) );
AND2_X2 _11957_ ( .A1(_04709_ ), .A2(_04710_ ), .ZN(_04711_ ) );
AND3_X1 _11958_ ( .A1(_04679_ ), .A2(_04708_ ), .A3(_04711_ ), .ZN(_04712_ ) );
NAND2_X1 _11959_ ( .A1(_04679_ ), .A2(_04708_ ), .ZN(_04713_ ) );
INV_X32 _11960_ ( .A(fanout_net_5 ), .ZN(_04714_ ) );
NOR2_X1 _11961_ ( .A1(_04714_ ), .A2(fanout_net_6 ), .ZN(_04715_ ) );
AND2_X2 _11962_ ( .A1(_04715_ ), .A2(_04710_ ), .ZN(_04716_ ) );
INV_X2 _11963_ ( .A(_04424_ ), .ZN(_04717_ ) );
BUF_X4 _11964_ ( .A(_04717_ ), .Z(_04718_ ) );
BUF_X4 _11965_ ( .A(_04718_ ), .Z(_04719_ ) );
NAND2_X1 _11966_ ( .A1(_04719_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04720_ ) );
BUF_X4 _11967_ ( .A(_04423_ ), .Z(_04721_ ) );
BUF_X4 _11968_ ( .A(_04431_ ), .Z(_04722_ ) );
NAND4_X1 _11969_ ( .A1(_04721_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04722_ ), .ZN(_04723_ ) );
NAND2_X1 _11970_ ( .A1(_04720_ ), .A2(_04723_ ), .ZN(_04724_ ) );
INV_X1 _11971_ ( .A(\EXU.r1_i [31] ), .ZN(_04725_ ) );
AND2_X1 _11972_ ( .A1(_04724_ ), .A2(_04725_ ), .ZN(_04726_ ) );
NOR2_X1 _11973_ ( .A1(_04724_ ), .A2(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ), .ZN(_04727_ ) );
NOR2_X1 _11974_ ( .A1(_04726_ ), .A2(_04727_ ), .ZN(_04728_ ) );
INV_X1 _11975_ ( .A(_04728_ ), .ZN(_04729_ ) );
BUF_X4 _11976_ ( .A(_04719_ ), .Z(_04730_ ) );
NAND2_X1 _11977_ ( .A1(_04730_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04731_ ) );
BUF_X4 _11978_ ( .A(_04721_ ), .Z(_04732_ ) );
NAND4_X1 _11979_ ( .A1(_04732_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04432_ ), .ZN(_04733_ ) );
NAND2_X1 _11980_ ( .A1(_04731_ ), .A2(_04733_ ), .ZN(_04734_ ) );
NOR2_X1 _11981_ ( .A1(_04734_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_A ), .ZN(_04735_ ) );
INV_X1 _11982_ ( .A(\EXU.r1_i [30] ), .ZN(_04736_ ) );
AND2_X1 _11983_ ( .A1(_04734_ ), .A2(_04736_ ), .ZN(_04737_ ) );
OAI21_X1 _11984_ ( .A(_04729_ ), .B1(_04735_ ), .B2(_04737_ ), .ZN(_04738_ ) );
NAND2_X1 _11985_ ( .A1(_04718_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_8_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04739_ ) );
NAND4_X1 _11986_ ( .A1(_04423_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_8_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04338_ ), .ZN(_04740_ ) );
NAND2_X1 _11987_ ( .A1(_04739_ ), .A2(_04740_ ), .ZN(_04741_ ) );
INV_X1 _11988_ ( .A(\EXU.r1_i [18] ), .ZN(_04742_ ) );
AND2_X1 _11989_ ( .A1(_04741_ ), .A2(_04742_ ), .ZN(_04743_ ) );
NOR2_X1 _11990_ ( .A1(_04741_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_13_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04744_ ) );
OR2_X1 _11991_ ( .A1(_04743_ ), .A2(_04744_ ), .ZN(_04745_ ) );
NAND2_X1 _11992_ ( .A1(_04718_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_7_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04746_ ) );
BUF_X4 _11993_ ( .A(_04423_ ), .Z(_04747_ ) );
NAND4_X1 _11994_ ( .A1(_04747_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_7_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04431_ ), .ZN(_04748_ ) );
NAND2_X1 _11995_ ( .A1(_04746_ ), .A2(_04748_ ), .ZN(_04749_ ) );
INV_X1 _11996_ ( .A(\EXU.r1_i [19] ), .ZN(_04750_ ) );
AND2_X1 _11997_ ( .A1(_04749_ ), .A2(_04750_ ), .ZN(_04751_ ) );
INV_X1 _11998_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_12_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04752_ ) );
AND3_X1 _11999_ ( .A1(_04746_ ), .A2(_04752_ ), .A3(_04748_ ), .ZN(_04753_ ) );
OAI21_X1 _12000_ ( .A(_04745_ ), .B1(_04751_ ), .B2(_04753_ ), .ZN(_04754_ ) );
INV_X1 _12001_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04755_ ) );
INV_X1 _12002_ ( .A(\EXU.r1_i [17] ), .ZN(_04756_ ) );
NAND2_X1 _12003_ ( .A1(_04718_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04757_ ) );
NAND4_X1 _12004_ ( .A1(_04423_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04338_ ), .ZN(_04758_ ) );
NAND2_X1 _12005_ ( .A1(_04757_ ), .A2(_04758_ ), .ZN(_04759_ ) );
MUX2_X1 _12006_ ( .A(_04755_ ), .B(_04756_ ), .S(_04759_ ), .Z(_04760_ ) );
NAND2_X1 _12007_ ( .A1(_04718_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ), .ZN(_04761_ ) );
NAND4_X1 _12008_ ( .A1(_04747_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A4(_04431_ ), .ZN(_04762_ ) );
NAND2_X1 _12009_ ( .A1(_04761_ ), .A2(_04762_ ), .ZN(_04763_ ) );
INV_X1 _12010_ ( .A(\EXU.r1_i [16] ), .ZN(_04764_ ) );
AND2_X1 _12011_ ( .A1(_04763_ ), .A2(_04764_ ), .ZN(_04765_ ) );
NOR2_X1 _12012_ ( .A1(_04763_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04766_ ) );
OAI21_X1 _12013_ ( .A(_04760_ ), .B1(_04765_ ), .B2(_04766_ ), .ZN(_04767_ ) );
NAND2_X1 _12014_ ( .A1(_04719_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ), .ZN(_04768_ ) );
NAND4_X1 _12015_ ( .A1(_04721_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A4(_04722_ ), .ZN(_04769_ ) );
NAND2_X1 _12016_ ( .A1(_04768_ ), .A2(_04769_ ), .ZN(_04770_ ) );
INV_X1 _12017_ ( .A(\EXU.r1_i [29] ), .ZN(_04771_ ) );
NAND2_X1 _12018_ ( .A1(_04770_ ), .A2(_04771_ ), .ZN(_04772_ ) );
OAI21_X1 _12019_ ( .A(_04772_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_2_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B2(_04770_ ), .ZN(_04773_ ) );
NAND2_X1 _12020_ ( .A1(_04730_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04774_ ) );
NAND4_X1 _12021_ ( .A1(_04732_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04432_ ), .ZN(_04775_ ) );
NAND2_X1 _12022_ ( .A1(_04774_ ), .A2(_04775_ ), .ZN(_04776_ ) );
NOR2_X1 _12023_ ( .A1(_04776_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_3_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04777_ ) );
INV_X1 _12024_ ( .A(\EXU.r1_i [28] ), .ZN(_04778_ ) );
AND2_X1 _12025_ ( .A1(_04776_ ), .A2(_04778_ ), .ZN(_04779_ ) );
OAI21_X1 _12026_ ( .A(_04773_ ), .B1(_04777_ ), .B2(_04779_ ), .ZN(_04780_ ) );
NOR4_X1 _12027_ ( .A1(_04738_ ), .A2(_04754_ ), .A3(_04767_ ), .A4(_04780_ ), .ZN(_04781_ ) );
NAND2_X1 _12028_ ( .A1(_04718_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_5_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04782_ ) );
NAND4_X1 _12029_ ( .A1(_04423_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_5_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04338_ ), .ZN(_04783_ ) );
NAND2_X1 _12030_ ( .A1(_04782_ ), .A2(_04783_ ), .ZN(_04784_ ) );
INV_X1 _12031_ ( .A(\EXU.r1_i [22] ), .ZN(_04785_ ) );
AND2_X1 _12032_ ( .A1(_04784_ ), .A2(_04785_ ), .ZN(_04786_ ) );
NOR2_X1 _12033_ ( .A1(_04784_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ), .ZN(_04787_ ) );
OR2_X1 _12034_ ( .A1(_04786_ ), .A2(_04787_ ), .ZN(_04788_ ) );
NAND2_X1 _12035_ ( .A1(_04718_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_4_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04789_ ) );
NAND4_X1 _12036_ ( .A1(_04747_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_4_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04431_ ), .ZN(_04790_ ) );
NAND2_X1 _12037_ ( .A1(_04789_ ), .A2(_04790_ ), .ZN(_04791_ ) );
INV_X1 _12038_ ( .A(\EXU.r1_i [23] ), .ZN(_04792_ ) );
AND2_X1 _12039_ ( .A1(_04791_ ), .A2(_04792_ ), .ZN(_04793_ ) );
INV_X1 _12040_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_8_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04794_ ) );
AND3_X1 _12041_ ( .A1(_04789_ ), .A2(_04794_ ), .A3(_04790_ ), .ZN(_04795_ ) );
OAI21_X1 _12042_ ( .A(_04788_ ), .B1(_04793_ ), .B2(_04795_ ), .ZN(_04796_ ) );
INV_X1 _12043_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_2_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04797_ ) );
OR2_X1 _12044_ ( .A1(_04424_ ), .A2(_04797_ ), .ZN(_04798_ ) );
NAND4_X1 _12045_ ( .A1(_04721_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_2_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04722_ ), .ZN(_04799_ ) );
NAND2_X1 _12046_ ( .A1(_04798_ ), .A2(_04799_ ), .ZN(_04800_ ) );
INV_X1 _12047_ ( .A(\EXU.r1_i [27] ), .ZN(_04801_ ) );
NAND2_X1 _12048_ ( .A1(_04800_ ), .A2(_04801_ ), .ZN(_04802_ ) );
OAI21_X1 _12049_ ( .A(_04802_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_4_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B2(_04800_ ), .ZN(_04803_ ) );
NAND2_X1 _12050_ ( .A1(_04719_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04804_ ) );
NAND4_X1 _12051_ ( .A1(_04721_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04722_ ), .ZN(_04805_ ) );
NAND2_X1 _12052_ ( .A1(_04804_ ), .A2(_04805_ ), .ZN(_04806_ ) );
NOR2_X1 _12053_ ( .A1(_04806_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_5_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04807_ ) );
INV_X1 _12054_ ( .A(\EXU.r1_i [26] ), .ZN(_04808_ ) );
AND2_X1 _12055_ ( .A1(_04806_ ), .A2(_04808_ ), .ZN(_04809_ ) );
OAI21_X1 _12056_ ( .A(_04803_ ), .B1(_04807_ ), .B2(_04809_ ), .ZN(_04810_ ) );
NAND2_X1 _12057_ ( .A1(_04719_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A ), .ZN(_04811_ ) );
NAND4_X1 _12058_ ( .A1(_04747_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A4(_04431_ ), .ZN(_04812_ ) );
NAND2_X1 _12059_ ( .A1(_04811_ ), .A2(_04812_ ), .ZN(_04813_ ) );
INV_X1 _12060_ ( .A(\EXU.r1_i [25] ), .ZN(_04814_ ) );
NAND2_X1 _12061_ ( .A1(_04813_ ), .A2(_04814_ ), .ZN(_04815_ ) );
OAI21_X1 _12062_ ( .A(_04815_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_6_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B2(_04813_ ), .ZN(_04816_ ) );
NAND2_X1 _12063_ ( .A1(_04730_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04817_ ) );
NAND4_X1 _12064_ ( .A1(_04732_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04722_ ), .ZN(_04818_ ) );
NAND2_X1 _12065_ ( .A1(_04817_ ), .A2(_04818_ ), .ZN(_04819_ ) );
NOR2_X1 _12066_ ( .A1(_04819_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ), .ZN(_04820_ ) );
INV_X1 _12067_ ( .A(\EXU.r1_i [24] ), .ZN(_04821_ ) );
AND2_X1 _12068_ ( .A1(_04819_ ), .A2(_04821_ ), .ZN(_04822_ ) );
OAI21_X1 _12069_ ( .A(_04816_ ), .B1(_04820_ ), .B2(_04822_ ), .ZN(_04823_ ) );
NAND2_X1 _12070_ ( .A1(_04718_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04824_ ) );
INV_X1 _12071_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04825_ ) );
NAND4_X1 _12072_ ( .A1(_04747_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04431_ ), .ZN(_04826_ ) );
NAND3_X1 _12073_ ( .A1(_04824_ ), .A2(_04825_ ), .A3(_04826_ ), .ZN(_04827_ ) );
NAND2_X1 _12074_ ( .A1(_04824_ ), .A2(_04826_ ), .ZN(_04828_ ) );
INV_X1 _12075_ ( .A(_04828_ ), .ZN(_04829_ ) );
OAI21_X1 _12076_ ( .A(_04827_ ), .B1(_04829_ ), .B2(\EXU.r1_i [21] ), .ZN(_04830_ ) );
NAND2_X1 _12077_ ( .A1(_04719_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ), .ZN(_04831_ ) );
NAND4_X1 _12078_ ( .A1(_04721_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A4(_04722_ ), .ZN(_04832_ ) );
NAND2_X1 _12079_ ( .A1(_04831_ ), .A2(_04832_ ), .ZN(_04833_ ) );
NOR2_X1 _12080_ ( .A1(_04833_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_11_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04834_ ) );
INV_X1 _12081_ ( .A(\EXU.r1_i [20] ), .ZN(_04835_ ) );
AND2_X1 _12082_ ( .A1(_04833_ ), .A2(_04835_ ), .ZN(_04836_ ) );
OAI21_X1 _12083_ ( .A(_04830_ ), .B1(_04834_ ), .B2(_04836_ ), .ZN(_04837_ ) );
NOR4_X1 _12084_ ( .A1(_04796_ ), .A2(_04810_ ), .A3(_04823_ ), .A4(_04837_ ), .ZN(_04838_ ) );
AND2_X1 _12085_ ( .A1(_04781_ ), .A2(_04838_ ), .ZN(_04839_ ) );
INV_X1 _12086_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_20_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04840_ ) );
INV_X1 _12087_ ( .A(\EXU.r1_i [11] ), .ZN(_04841_ ) );
NAND2_X1 _12088_ ( .A1(_04719_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04842_ ) );
NAND4_X1 _12089_ ( .A1(_04721_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04722_ ), .ZN(_04843_ ) );
NAND2_X1 _12090_ ( .A1(_04842_ ), .A2(_04843_ ), .ZN(_04844_ ) );
MUX2_X1 _12091_ ( .A(_04840_ ), .B(_04841_ ), .S(_04844_ ), .Z(_04845_ ) );
NAND2_X1 _12092_ ( .A1(_04730_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_14_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04846_ ) );
NAND4_X1 _12093_ ( .A1(_04732_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_14_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(fanout_net_8 ), .A4(_04432_ ), .ZN(_04847_ ) );
NAND2_X1 _12094_ ( .A1(_04846_ ), .A2(_04847_ ), .ZN(_04848_ ) );
INV_X1 _12095_ ( .A(\EXU.r1_i [10] ), .ZN(_04849_ ) );
NAND2_X1 _12096_ ( .A1(_04848_ ), .A2(_04849_ ), .ZN(_04850_ ) );
OAI21_X1 _12097_ ( .A(_04850_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_21_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B2(_04848_ ), .ZN(_04851_ ) );
AND2_X1 _12098_ ( .A1(_04845_ ), .A2(_04851_ ), .ZN(_04852_ ) );
NAND2_X1 _12099_ ( .A1(_04730_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_10_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04853_ ) );
INV_X1 _12100_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_16_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04854_ ) );
NAND4_X1 _12101_ ( .A1(_04732_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_10_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04432_ ), .ZN(_04855_ ) );
NAND3_X1 _12102_ ( .A1(_04853_ ), .A2(_04854_ ), .A3(_04855_ ), .ZN(_04856_ ) );
NAND2_X1 _12103_ ( .A1(_04853_ ), .A2(_04855_ ), .ZN(_04857_ ) );
INV_X1 _12104_ ( .A(_04857_ ), .ZN(_04858_ ) );
OAI21_X1 _12105_ ( .A(_04856_ ), .B1(_04858_ ), .B2(\EXU.r1_i [15] ), .ZN(_04859_ ) );
NAND2_X1 _12106_ ( .A1(_04730_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_11_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04860_ ) );
NAND4_X1 _12107_ ( .A1(_04732_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_11_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04432_ ), .ZN(_04861_ ) );
NAND2_X1 _12108_ ( .A1(_04860_ ), .A2(_04861_ ), .ZN(_04862_ ) );
NOR2_X1 _12109_ ( .A1(_04862_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04863_ ) );
INV_X1 _12110_ ( .A(\EXU.r1_i [14] ), .ZN(_04864_ ) );
AND2_X1 _12111_ ( .A1(_04862_ ), .A2(_04864_ ), .ZN(_04865_ ) );
OAI21_X1 _12112_ ( .A(_04859_ ), .B1(_04863_ ), .B2(_04865_ ), .ZN(_04866_ ) );
NAND2_X1 _12113_ ( .A1(_04719_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04867_ ) );
NAND4_X1 _12114_ ( .A1(_04721_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04722_ ), .ZN(_04868_ ) );
NAND2_X1 _12115_ ( .A1(_04867_ ), .A2(_04868_ ), .ZN(_04869_ ) );
OR2_X1 _12116_ ( .A1(_04869_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04870_ ) );
INV_X1 _12117_ ( .A(_04869_ ), .ZN(_04871_ ) );
OAI21_X1 _12118_ ( .A(_04870_ ), .B1(_04871_ ), .B2(\EXU.r1_i [13] ), .ZN(_04872_ ) );
NAND2_X1 _12119_ ( .A1(_04730_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ), .ZN(_04873_ ) );
NAND4_X1 _12120_ ( .A1(_04732_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A4(_04432_ ), .ZN(_04874_ ) );
NAND2_X1 _12121_ ( .A1(_04873_ ), .A2(_04874_ ), .ZN(_04875_ ) );
NOR2_X1 _12122_ ( .A1(_04875_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_19_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04876_ ) );
INV_X1 _12123_ ( .A(\EXU.r1_i [12] ), .ZN(_04877_ ) );
AND2_X1 _12124_ ( .A1(_04875_ ), .A2(_04877_ ), .ZN(_04878_ ) );
OAI21_X1 _12125_ ( .A(_04872_ ), .B1(_04876_ ), .B2(_04878_ ), .ZN(_04879_ ) );
INV_X1 _12126_ ( .A(\LSU.ls_wdata_i_$_MUX__Y_20_A_$_ANDNOT__Y_B ), .ZN(_04880_ ) );
OR2_X1 _12127_ ( .A1(_04424_ ), .A2(_04880_ ), .ZN(_04881_ ) );
INV_X1 _12128_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04882_ ) );
NAND4_X1 _12129_ ( .A1(_04423_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_21_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04338_ ), .ZN(_04883_ ) );
NAND3_X1 _12130_ ( .A1(_04881_ ), .A2(_04882_ ), .A3(_04883_ ), .ZN(_04884_ ) );
NAND2_X2 _12131_ ( .A1(_04881_ ), .A2(_04883_ ), .ZN(_04885_ ) );
INV_X1 _12132_ ( .A(_04885_ ), .ZN(_04886_ ) );
OAI21_X1 _12133_ ( .A(_04884_ ), .B1(_04886_ ), .B2(\EXU.r1_i [3] ), .ZN(_04887_ ) );
INV_X1 _12134_ ( .A(\LSU.ls_wdata_i_$_MUX__Y_21_A_$_ANDNOT__Y_B ), .ZN(_04888_ ) );
OR2_X1 _12135_ ( .A1(_04424_ ), .A2(_04888_ ), .ZN(_04889_ ) );
NAND4_X1 _12136_ ( .A1(_04747_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .A4(_04431_ ), .ZN(_04890_ ) );
AND3_X1 _12137_ ( .A1(_04889_ ), .A2(_04458_ ), .A3(_04890_ ), .ZN(_04891_ ) );
NAND2_X1 _12138_ ( .A1(_04889_ ), .A2(_04890_ ), .ZN(_04892_ ) );
INV_X1 _12139_ ( .A(\EXU.r1_i [2] ), .ZN(_04893_ ) );
AND2_X1 _12140_ ( .A1(_04892_ ), .A2(_04893_ ), .ZN(_04894_ ) );
OAI21_X1 _12141_ ( .A(_04887_ ), .B1(_04891_ ), .B2(_04894_ ), .ZN(_04895_ ) );
INV_X1 _12142_ ( .A(\LSU.ls_wdata_i_$_MUX__Y_22_A_$_ANDNOT__Y_B ), .ZN(_04896_ ) );
OR2_X1 _12143_ ( .A1(_04424_ ), .A2(_04896_ ), .ZN(_04897_ ) );
INV_X1 _12144_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04898_ ) );
NAND4_X1 _12145_ ( .A1(_04747_ ), .A2(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(fanout_net_8 ), .A4(_04431_ ), .ZN(_04899_ ) );
NAND3_X1 _12146_ ( .A1(_04897_ ), .A2(_04898_ ), .A3(_04899_ ), .ZN(_04900_ ) );
NAND2_X2 _12147_ ( .A1(_04897_ ), .A2(_04899_ ), .ZN(_04901_ ) );
INV_X1 _12148_ ( .A(_04901_ ), .ZN(_04902_ ) );
OAI21_X1 _12149_ ( .A(_04900_ ), .B1(_04902_ ), .B2(\EXU.r1_i [1] ), .ZN(_04903_ ) );
INV_X1 _12150_ ( .A(\EXU.r2_i [0] ), .ZN(_04904_ ) );
OR2_X1 _12151_ ( .A1(_04424_ ), .A2(_04904_ ), .ZN(_04905_ ) );
BUF_X2 _12152_ ( .A(_04905_ ), .Z(_04906_ ) );
NAND4_X2 _12153_ ( .A1(_04747_ ), .A2(\EXU.imm_i [0] ), .A3(fanout_net_8 ), .A4(_04338_ ), .ZN(_04907_ ) );
NAND2_X2 _12154_ ( .A1(_04906_ ), .A2(_04907_ ), .ZN(_04908_ ) );
INV_X1 _12155_ ( .A(_04908_ ), .ZN(_04909_ ) );
AND2_X1 _12156_ ( .A1(_04909_ ), .A2(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_A ), .ZN(_04910_ ) );
INV_X1 _12157_ ( .A(\EXU.r1_i [0] ), .ZN(_04911_ ) );
AOI21_X1 _12158_ ( .A(_04911_ ), .B1(_04906_ ), .B2(_04907_ ), .ZN(_04912_ ) );
OAI21_X1 _12159_ ( .A(_04903_ ), .B1(_04910_ ), .B2(_04912_ ), .ZN(_04913_ ) );
NOR4_X1 _12160_ ( .A1(_04866_ ), .A2(_04879_ ), .A3(_04895_ ), .A4(_04913_ ), .ZN(_04914_ ) );
NAND2_X1 _12161_ ( .A1(_04730_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_15_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04915_ ) );
NAND4_X1 _12162_ ( .A1(_04732_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_15_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04432_ ), .ZN(_04916_ ) );
NAND2_X1 _12163_ ( .A1(_04915_ ), .A2(_04916_ ), .ZN(_04917_ ) );
INV_X1 _12164_ ( .A(\EXU.r1_i [9] ), .ZN(_04918_ ) );
AND2_X1 _12165_ ( .A1(_04917_ ), .A2(_04918_ ), .ZN(_04919_ ) );
NOR2_X1 _12166_ ( .A1(_04917_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_22_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04920_ ) );
NOR2_X1 _12167_ ( .A1(_04919_ ), .A2(_04920_ ), .ZN(_04921_ ) );
NAND2_X1 _12168_ ( .A1(_04730_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_16_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ), .ZN(_04922_ ) );
NAND4_X1 _12169_ ( .A1(_04732_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_16_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04432_ ), .ZN(_04923_ ) );
NAND2_X1 _12170_ ( .A1(_04922_ ), .A2(_04923_ ), .ZN(_04924_ ) );
OR2_X1 _12171_ ( .A1(_04924_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04925_ ) );
INV_X1 _12172_ ( .A(\EXU.r1_i [8] ), .ZN(_04926_ ) );
NAND2_X1 _12173_ ( .A1(_04924_ ), .A2(_04926_ ), .ZN(_04927_ ) );
AOI21_X1 _12174_ ( .A(_04921_ ), .B1(_04925_ ), .B2(_04927_ ), .ZN(_04928_ ) );
INV_X1 _12175_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_24_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04929_ ) );
INV_X1 _12176_ ( .A(\EXU.r1_i [7] ), .ZN(_04930_ ) );
NOR2_X1 _12177_ ( .A1(_04718_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_17_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_04931_ ) );
AOI21_X1 _12178_ ( .A(\LSU.ls_wdata_i_$_MUX__Y_16_A_$_ANDNOT__Y_B ), .B1(_04387_ ), .B2(_04747_ ), .ZN(_04932_ ) );
NOR2_X1 _12179_ ( .A1(_04931_ ), .A2(_04932_ ), .ZN(_04933_ ) );
MUX2_X1 _12180_ ( .A(_04929_ ), .B(_04930_ ), .S(_04933_ ), .Z(_04934_ ) );
NAND2_X1 _12181_ ( .A1(_04719_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_17_A_$_ANDNOT__Y_B ), .ZN(_04935_ ) );
INV_X1 _12182_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04936_ ) );
NAND4_X1 _12183_ ( .A1(_04721_ ), .A2(fanout_net_8 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_18_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04722_ ), .ZN(_04937_ ) );
AND3_X1 _12184_ ( .A1(_04935_ ), .A2(_04936_ ), .A3(_04937_ ), .ZN(_04938_ ) );
NAND2_X1 _12185_ ( .A1(_04935_ ), .A2(_04937_ ), .ZN(_04939_ ) );
INV_X1 _12186_ ( .A(\EXU.r1_i [6] ), .ZN(_04940_ ) );
AND2_X1 _12187_ ( .A1(_04939_ ), .A2(_04940_ ), .ZN(_04941_ ) );
OAI21_X1 _12188_ ( .A(_04934_ ), .B1(_04938_ ), .B2(_04941_ ), .ZN(_04942_ ) );
NAND2_X1 _12189_ ( .A1(_04719_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_18_A_$_ANDNOT__Y_B ), .ZN(_04943_ ) );
INV_X1 _12190_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_26_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04944_ ) );
NAND4_X1 _12191_ ( .A1(_04721_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_19_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04722_ ), .ZN(_04945_ ) );
NAND3_X1 _12192_ ( .A1(_04943_ ), .A2(_04944_ ), .A3(_04945_ ), .ZN(_04946_ ) );
NAND2_X1 _12193_ ( .A1(_04943_ ), .A2(_04945_ ), .ZN(_04947_ ) );
INV_X1 _12194_ ( .A(_04947_ ), .ZN(_04948_ ) );
OAI21_X1 _12195_ ( .A(_04946_ ), .B1(_04948_ ), .B2(\EXU.r1_i [5] ), .ZN(_04949_ ) );
NAND2_X1 _12196_ ( .A1(_04718_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_19_A_$_ANDNOT__Y_B ), .ZN(_04950_ ) );
INV_X1 _12197_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_27_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_04951_ ) );
NAND4_X1 _12198_ ( .A1(_04747_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_20_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04431_ ), .ZN(_04952_ ) );
AND3_X1 _12199_ ( .A1(_04950_ ), .A2(_04951_ ), .A3(_04952_ ), .ZN(_04953_ ) );
NAND2_X2 _12200_ ( .A1(_04950_ ), .A2(_04952_ ), .ZN(_04954_ ) );
INV_X1 _12201_ ( .A(\EXU.r1_i [4] ), .ZN(_04955_ ) );
AND2_X1 _12202_ ( .A1(_04954_ ), .A2(_04955_ ), .ZN(_04956_ ) );
OAI21_X1 _12203_ ( .A(_04949_ ), .B1(_04953_ ), .B2(_04956_ ), .ZN(_04957_ ) );
NOR2_X1 _12204_ ( .A1(_04942_ ), .A2(_04957_ ), .ZN(_04958_ ) );
AND4_X1 _12205_ ( .A1(_04852_ ), .A2(_04914_ ), .A3(_04928_ ), .A4(_04958_ ), .ZN(_04959_ ) );
AND2_X1 _12206_ ( .A1(_04839_ ), .A2(_04959_ ), .ZN(_04960_ ) );
NAND2_X1 _12207_ ( .A1(_04382_ ), .A2(_04385_ ), .ZN(_04961_ ) );
NOR2_X1 _12208_ ( .A1(_04823_ ), .A2(_04810_ ), .ZN(_04962_ ) );
AND3_X1 _12209_ ( .A1(_04761_ ), .A2(_04764_ ), .A3(_04762_ ), .ZN(_04963_ ) );
AND2_X1 _12210_ ( .A1(_04760_ ), .A2(_04963_ ), .ZN(_04964_ ) );
AND3_X1 _12211_ ( .A1(_04757_ ), .A2(_04756_ ), .A3(_04758_ ), .ZN(_04965_ ) );
OAI221_X1 _12212_ ( .A(_04745_ ), .B1(_04751_ ), .B2(_04753_ ), .C1(_04964_ ), .C2(_04965_ ), .ZN(_04966_ ) );
AOI21_X1 _12213_ ( .A(_04753_ ), .B1(_04750_ ), .B2(_04749_ ), .ZN(_04967_ ) );
NAND3_X1 _12214_ ( .A1(_04739_ ), .A2(_04742_ ), .A3(_04740_ ), .ZN(_04968_ ) );
OAI221_X1 _12215_ ( .A(_04966_ ), .B1(\EXU.r1_i [19] ), .B2(_04749_ ), .C1(_04967_ ), .C2(_04968_ ), .ZN(_04969_ ) );
NOR2_X1 _12216_ ( .A1(_04796_ ), .A2(_04837_ ), .ZN(_04970_ ) );
AND2_X1 _12217_ ( .A1(_04969_ ), .A2(_04970_ ), .ZN(_04971_ ) );
AND3_X1 _12218_ ( .A1(_04831_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_11_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A3(_04832_ ), .ZN(_04972_ ) );
INV_X1 _12219_ ( .A(\EXU.r1_i [21] ), .ZN(_04973_ ) );
AOI22_X1 _12220_ ( .A1(_04830_ ), .A2(_04972_ ), .B1(_04973_ ), .B2(_04829_ ), .ZN(_04974_ ) );
OR2_X1 _12221_ ( .A1(_04796_ ), .A2(_04974_ ), .ZN(_04975_ ) );
AOI21_X1 _12222_ ( .A(_04795_ ), .B1(_04792_ ), .B2(_04791_ ), .ZN(_04976_ ) );
NAND3_X1 _12223_ ( .A1(_04782_ ), .A2(_04785_ ), .A3(_04783_ ), .ZN(_04977_ ) );
OAI221_X1 _12224_ ( .A(_04975_ ), .B1(\EXU.r1_i [23] ), .B2(_04791_ ), .C1(_04976_ ), .C2(_04977_ ), .ZN(_04978_ ) );
OAI21_X1 _12225_ ( .A(_04962_ ), .B1(_04971_ ), .B2(_04978_ ), .ZN(_04979_ ) );
AND3_X1 _12226_ ( .A1(_04817_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ), .A3(_04818_ ), .ZN(_04980_ ) );
AND2_X1 _12227_ ( .A1(_04816_ ), .A2(_04980_ ), .ZN(_04981_ ) );
AND3_X1 _12228_ ( .A1(_04811_ ), .A2(_04814_ ), .A3(_04812_ ), .ZN(_04982_ ) );
OAI221_X1 _12229_ ( .A(_04803_ ), .B1(_04807_ ), .B2(_04809_ ), .C1(_04981_ ), .C2(_04982_ ), .ZN(_04983_ ) );
BUF_X4 _12230_ ( .A(_04424_ ), .Z(_04984_ ) );
OAI211_X1 _12231_ ( .A(_04801_ ), .B(_04799_ ), .C1(_04984_ ), .C2(_04797_ ), .ZN(_04985_ ) );
NAND4_X1 _12232_ ( .A1(_04803_ ), .A2(_04808_ ), .A3(_04804_ ), .A4(_04805_ ), .ZN(_04986_ ) );
AND3_X1 _12233_ ( .A1(_04983_ ), .A2(_04985_ ), .A3(_04986_ ), .ZN(_04987_ ) );
AOI211_X1 _12234_ ( .A(_04738_ ), .B(_04780_ ), .C1(_04979_ ), .C2(_04987_ ), .ZN(_04988_ ) );
NAND3_X1 _12235_ ( .A1(_04768_ ), .A2(_04771_ ), .A3(_04769_ ), .ZN(_04989_ ) );
AND3_X1 _12236_ ( .A1(_04774_ ), .A2(_04778_ ), .A3(_04775_ ), .ZN(_04990_ ) );
NAND2_X1 _12237_ ( .A1(_04773_ ), .A2(_04990_ ), .ZN(_04991_ ) );
AOI21_X1 _12238_ ( .A(_04738_ ), .B1(_04989_ ), .B2(_04991_ ), .ZN(_04992_ ) );
AND3_X1 _12239_ ( .A1(_04720_ ), .A2(_04725_ ), .A3(_04723_ ), .ZN(_04993_ ) );
NOR3_X1 _12240_ ( .A1(_04728_ ), .A2(\EXU.r1_i [30] ), .A3(_04734_ ), .ZN(_04994_ ) );
NOR4_X1 _12241_ ( .A1(_04988_ ), .A2(_04992_ ), .A3(_04993_ ), .A4(_04994_ ), .ZN(_04995_ ) );
INV_X1 _12242_ ( .A(_04892_ ), .ZN(_04996_ ) );
NAND3_X1 _12243_ ( .A1(_04887_ ), .A2(_04893_ ), .A3(_04996_ ), .ZN(_04997_ ) );
NOR2_X1 _12244_ ( .A1(_04908_ ), .A2(_04911_ ), .ZN(_04998_ ) );
INV_X1 _12245_ ( .A(_04998_ ), .ZN(_04999_ ) );
INV_X1 _12246_ ( .A(\EXU.r1_i [1] ), .ZN(_05000_ ) );
AOI22_X1 _12247_ ( .A1(_04903_ ), .A2(_04999_ ), .B1(_05000_ ), .B2(_04902_ ), .ZN(_05001_ ) );
OAI221_X1 _12248_ ( .A(_04997_ ), .B1(\EXU.r1_i [3] ), .B2(_04885_ ), .C1(_05001_ ), .C2(_04895_ ), .ZN(_05002_ ) );
AND2_X1 _12249_ ( .A1(_04958_ ), .A2(_05002_ ), .ZN(_05003_ ) );
NAND4_X1 _12250_ ( .A1(_04934_ ), .A2(_04940_ ), .A3(_04935_ ), .A4(_04937_ ), .ZN(_05004_ ) );
AND3_X1 _12251_ ( .A1(_04950_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_27_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A3(_04952_ ), .ZN(_05005_ ) );
INV_X1 _12252_ ( .A(\EXU.r1_i [5] ), .ZN(_05006_ ) );
AOI22_X1 _12253_ ( .A1(_04949_ ), .A2(_05005_ ), .B1(_05006_ ), .B2(_04948_ ), .ZN(_05007_ ) );
OAI221_X1 _12254_ ( .A(_05004_ ), .B1(\EXU.r1_i [7] ), .B2(_04933_ ), .C1(_04942_ ), .C2(_05007_ ), .ZN(_05008_ ) );
OAI211_X1 _12255_ ( .A(_04852_ ), .B(_04928_ ), .C1(_05003_ ), .C2(_05008_ ), .ZN(_05009_ ) );
NAND4_X1 _12256_ ( .A1(_04845_ ), .A2(_04849_ ), .A3(_04846_ ), .A4(_04847_ ), .ZN(_05010_ ) );
OAI21_X1 _12257_ ( .A(_05010_ ), .B1(\EXU.r1_i [11] ), .B2(_04844_ ), .ZN(_05011_ ) );
NAND3_X1 _12258_ ( .A1(_04922_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_04923_ ), .ZN(_05012_ ) );
OAI22_X1 _12259_ ( .A1(_04921_ ), .A2(_05012_ ), .B1(\EXU.r1_i [9] ), .B2(_04917_ ), .ZN(_05013_ ) );
AOI21_X1 _12260_ ( .A(_05011_ ), .B1(_04852_ ), .B2(_05013_ ), .ZN(_05014_ ) );
AOI211_X1 _12261_ ( .A(_04866_ ), .B(_04879_ ), .C1(_05009_ ), .C2(_05014_ ), .ZN(_05015_ ) );
AND3_X1 _12262_ ( .A1(_04860_ ), .A2(_04864_ ), .A3(_04861_ ), .ZN(_05016_ ) );
INV_X1 _12263_ ( .A(\EXU.r1_i [15] ), .ZN(_05017_ ) );
AOI22_X1 _12264_ ( .A1(_04859_ ), .A2(_05016_ ), .B1(_05017_ ), .B2(_04858_ ), .ZN(_05018_ ) );
AND3_X1 _12265_ ( .A1(_04873_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_19_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A3(_04874_ ), .ZN(_05019_ ) );
INV_X1 _12266_ ( .A(\EXU.r1_i [13] ), .ZN(_05020_ ) );
AOI22_X1 _12267_ ( .A1(_04872_ ), .A2(_05019_ ), .B1(_05020_ ), .B2(_04871_ ), .ZN(_05021_ ) );
OAI21_X1 _12268_ ( .A(_05018_ ), .B1(_05021_ ), .B2(_04866_ ), .ZN(_05022_ ) );
OAI21_X1 _12269_ ( .A(_04839_ ), .B1(_05015_ ), .B2(_05022_ ), .ZN(_05023_ ) );
NAND2_X1 _12270_ ( .A1(_04995_ ), .A2(_05023_ ), .ZN(_05024_ ) );
NAND3_X1 _12271_ ( .A1(_04710_ ), .A2(_04714_ ), .A3(fanout_net_6 ), .ZN(_05025_ ) );
INV_X1 _12272_ ( .A(fanout_net_10 ), .ZN(_05026_ ) );
AOI22_X1 _12273_ ( .A1(_04715_ ), .A2(_05026_ ), .B1(_04709_ ), .B2(\EXU.funct3_i [2] ), .ZN(_05027_ ) );
AOI21_X1 _12274_ ( .A(_04729_ ), .B1(_05025_ ), .B2(_05027_ ), .ZN(_05028_ ) );
AOI221_X4 _12275_ ( .A(_04960_ ), .B1(_04425_ ), .B2(_04961_ ), .C1(_05024_ ), .C2(_05028_ ), .ZN(_05029_ ) );
OR2_X1 _12276_ ( .A1(_05024_ ), .A2(_05028_ ), .ZN(_05030_ ) );
AND2_X1 _12277_ ( .A1(_05029_ ), .A2(_05030_ ), .ZN(_05031_ ) );
XNOR2_X1 _12278_ ( .A(_05031_ ), .B(_04714_ ), .ZN(_05032_ ) );
AOI221_X4 _12279_ ( .A(_04712_ ), .B1(_04713_ ), .B2(_04716_ ), .C1(_05032_ ), .C2(_05026_ ), .ZN(_05033_ ) );
NOR2_X1 _12280_ ( .A1(_05033_ ), .A2(_04961_ ), .ZN(_05034_ ) );
AND2_X1 _12281_ ( .A1(\EXU.op_i [1] ), .A2(\EXU.op_i [0] ), .ZN(_05035_ ) );
AND2_X1 _12282_ ( .A1(_04415_ ), .A2(_05035_ ), .ZN(_05036_ ) );
NOR2_X1 _12283_ ( .A1(_04418_ ), .A2(_05036_ ), .ZN(_05037_ ) );
INV_X1 _12284_ ( .A(_05037_ ), .ZN(_05038_ ) );
BUF_X2 _12285_ ( .A(_05038_ ), .Z(_05039_ ) );
NOR2_X1 _12286_ ( .A1(_05034_ ), .A2(_05039_ ), .ZN(_05040_ ) );
BUF_X4 _12287_ ( .A(_05040_ ), .Z(_05041_ ) );
BUF_X4 _12288_ ( .A(_05041_ ), .Z(_05042_ ) );
NOR2_X1 _12289_ ( .A1(_04653_ ), .A2(_05042_ ), .ZN(_05043_ ) );
BUF_X4 _12290_ ( .A(_04343_ ), .Z(_05044_ ) );
BUF_X2 _12291_ ( .A(_05044_ ), .Z(_05045_ ) );
BUF_X2 _12292_ ( .A(_04348_ ), .Z(_05046_ ) );
CLKBUF_X3 _12293_ ( .A(_05046_ ), .Z(_05047_ ) );
AND3_X1 _12294_ ( .A1(_05045_ ), .A2(\EXU.mtvec_i [31] ), .A3(_05047_ ), .ZN(_05048_ ) );
INV_X1 _12295_ ( .A(_05040_ ), .ZN(_05049_ ) );
BUF_X4 _12296_ ( .A(_04360_ ), .Z(_05050_ ) );
BUF_X2 _12297_ ( .A(_05050_ ), .Z(_05051_ ) );
NOR2_X1 _12298_ ( .A1(_04346_ ), .A2(\EXU.imm_i [6] ), .ZN(_05052_ ) );
AND3_X2 _12299_ ( .A1(_04334_ ), .A2(_04344_ ), .A3(_05052_ ), .ZN(_05053_ ) );
BUF_X2 _12300_ ( .A(_05053_ ), .Z(_05054_ ) );
BUF_X4 _12301_ ( .A(_04340_ ), .Z(_05055_ ) );
NAND4_X1 _12302_ ( .A1(_05054_ ), .A2(fanout_net_7 ), .A3(\EXU.mepc_i [31] ), .A4(_05055_ ), .ZN(_05056_ ) );
AND2_X1 _12303_ ( .A1(\EXU.pc_i [3] ), .A2(\EXU.pc_i [2] ), .ZN(_05057_ ) );
AND2_X1 _12304_ ( .A1(_05057_ ), .A2(\EXU.pc_i [4] ), .ZN(_05058_ ) );
AND2_X1 _12305_ ( .A1(_05058_ ), .A2(\EXU.pc_i [5] ), .ZN(_05059_ ) );
AND2_X1 _12306_ ( .A1(_05059_ ), .A2(\EXU.pc_i [6] ), .ZN(_05060_ ) );
AND2_X1 _12307_ ( .A1(_05060_ ), .A2(\EXU.pc_i [7] ), .ZN(_05061_ ) );
AND3_X1 _12308_ ( .A1(_05061_ ), .A2(\EXU.pc_i [9] ), .A3(\EXU.pc_i [8] ), .ZN(_05062_ ) );
AND3_X1 _12309_ ( .A1(_05062_ ), .A2(\EXU.pc_i [11] ), .A3(\EXU.pc_i [10] ), .ZN(_05063_ ) );
AND3_X1 _12310_ ( .A1(_05063_ ), .A2(\EXU.pc_i [13] ), .A3(\EXU.pc_i [12] ), .ZN(_05064_ ) );
AND3_X1 _12311_ ( .A1(_05064_ ), .A2(\EXU.pc_i [15] ), .A3(\EXU.pc_i [14] ), .ZN(_05065_ ) );
AND3_X1 _12312_ ( .A1(_05065_ ), .A2(\EXU.pc_i [17] ), .A3(\EXU.pc_i [16] ), .ZN(_05066_ ) );
AND3_X1 _12313_ ( .A1(_05066_ ), .A2(\EXU.pc_i [19] ), .A3(\EXU.pc_i [18] ), .ZN(_05067_ ) );
AND3_X1 _12314_ ( .A1(_05067_ ), .A2(\EXU.pc_i [21] ), .A3(\EXU.pc_i [20] ), .ZN(_05068_ ) );
AND3_X1 _12315_ ( .A1(_05068_ ), .A2(\EXU.pc_i [23] ), .A3(\EXU.pc_i [22] ), .ZN(_05069_ ) );
AND3_X1 _12316_ ( .A1(_05069_ ), .A2(\EXU.pc_i [25] ), .A3(\EXU.pc_i [24] ), .ZN(_05070_ ) );
AND3_X1 _12317_ ( .A1(_05070_ ), .A2(\EXU.pc_i [27] ), .A3(\EXU.pc_i [26] ), .ZN(_05071_ ) );
AND2_X1 _12318_ ( .A1(_05071_ ), .A2(\EXU.pc_i [28] ), .ZN(_05072_ ) );
NAND2_X1 _12319_ ( .A1(_05072_ ), .A2(\EXU.pc_i [29] ), .ZN(_05073_ ) );
NOR2_X1 _12320_ ( .A1(_05073_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_B ), .ZN(_05074_ ) );
XNOR2_X1 _12321_ ( .A(_05074_ ), .B(\EXU.pc_i [31] ), .ZN(_05075_ ) );
AND2_X1 _12322_ ( .A1(_04343_ ), .A2(_05053_ ), .ZN(_05076_ ) );
BUF_X4 _12323_ ( .A(_05076_ ), .Z(_05077_ ) );
OAI21_X1 _12324_ ( .A(_05056_ ), .B1(_05075_ ), .B2(_05077_ ), .ZN(_05078_ ) );
AOI211_X1 _12325_ ( .A(_05048_ ), .B(_05049_ ), .C1(_05051_ ), .C2(_05078_ ), .ZN(_05079_ ) );
NOR2_X1 _12326_ ( .A1(_04331_ ), .A2(fanout_net_11 ), .ZN(_05080_ ) );
AND2_X1 _12327_ ( .A1(_05080_ ), .A2(_04397_ ), .ZN(_05081_ ) );
AND2_X2 _12328_ ( .A1(_04393_ ), .A2(_05081_ ), .ZN(_05082_ ) );
INV_X1 _12329_ ( .A(_05082_ ), .ZN(_05083_ ) );
OR2_X1 _12330_ ( .A1(_05079_ ), .A2(_05083_ ), .ZN(_05084_ ) );
INV_X1 _12331_ ( .A(\EXU.dnpc_o [31] ), .ZN(_05085_ ) );
INV_X1 _12332_ ( .A(_05080_ ), .ZN(_05086_ ) );
OR2_X2 _12333_ ( .A1(_05082_ ), .A2(_05086_ ), .ZN(_05087_ ) );
BUF_X4 _12334_ ( .A(_05087_ ), .Z(_05088_ ) );
OAI22_X1 _12335_ ( .A1(_05043_ ), .A2(_05084_ ), .B1(_05085_ ), .B2(_05088_ ), .ZN(_00203_ ) );
XOR2_X1 _12336_ ( .A(_04646_ ), .B(_04648_ ), .Z(_05089_ ) );
AND2_X1 _12337_ ( .A1(_05089_ ), .A2(_05049_ ), .ZN(_05090_ ) );
BUF_X4 _12338_ ( .A(_05041_ ), .Z(_05091_ ) );
BUF_X4 _12339_ ( .A(_05047_ ), .Z(_05092_ ) );
BUF_X4 _12340_ ( .A(_05092_ ), .Z(_05093_ ) );
BUF_X4 _12341_ ( .A(_05055_ ), .Z(_05094_ ) );
NAND4_X1 _12342_ ( .A1(_05093_ ), .A2(fanout_net_7 ), .A3(\EXU.mtvec_i [30] ), .A4(_05094_ ), .ZN(_05095_ ) );
CLKBUF_X2 _12343_ ( .A(_04340_ ), .Z(_05096_ ) );
AND4_X1 _12344_ ( .A1(fanout_net_7 ), .A2(_05054_ ), .A3(\EXU.mepc_i [30] ), .A4(_05096_ ), .ZN(_05097_ ) );
XNOR2_X1 _12345_ ( .A(_05073_ ), .B(\EXU.pc_i [30] ), .ZN(_05098_ ) );
INV_X1 _12346_ ( .A(_05076_ ), .ZN(_05099_ ) );
BUF_X4 _12347_ ( .A(_05099_ ), .Z(_05100_ ) );
BUF_X4 _12348_ ( .A(_05100_ ), .Z(_05101_ ) );
AOI21_X1 _12349_ ( .A(_05097_ ), .B1(_05098_ ), .B2(_05101_ ), .ZN(_05102_ ) );
BUF_X4 _12350_ ( .A(_04359_ ), .Z(_05103_ ) );
BUF_X4 _12351_ ( .A(_05103_ ), .Z(_05104_ ) );
OAI21_X1 _12352_ ( .A(_05095_ ), .B1(_05102_ ), .B2(_05104_ ), .ZN(_05105_ ) );
AOI21_X1 _12353_ ( .A(_05090_ ), .B1(_05091_ ), .B2(_05105_ ), .ZN(_05106_ ) );
INV_X1 _12354_ ( .A(\EXU.dnpc_o [30] ), .ZN(_05107_ ) );
OAI22_X1 _12355_ ( .A1(_05106_ ), .A2(_05083_ ), .B1(_05107_ ), .B2(_05088_ ), .ZN(_00204_ ) );
AND2_X1 _12356_ ( .A1(_04564_ ), .A2(_04597_ ), .ZN(_05108_ ) );
NAND2_X1 _12357_ ( .A1(_04550_ ), .A2(_04583_ ), .ZN(_05109_ ) );
AND2_X1 _12358_ ( .A1(_04590_ ), .A2(_04595_ ), .ZN(_05110_ ) );
AND2_X1 _12359_ ( .A1(_05109_ ), .A2(_05110_ ), .ZN(_05111_ ) );
INV_X1 _12360_ ( .A(_05111_ ), .ZN(_05112_ ) );
AOI21_X1 _12361_ ( .A(_05108_ ), .B1(_05112_ ), .B2(_04566_ ), .ZN(_05113_ ) );
XNOR2_X1 _12362_ ( .A(_05113_ ), .B(_04563_ ), .ZN(_05114_ ) );
NOR2_X1 _12363_ ( .A1(_05114_ ), .A2(_05042_ ), .ZN(_05115_ ) );
BUF_X4 _12364_ ( .A(_05082_ ), .Z(_05116_ ) );
BUF_X4 _12365_ ( .A(_05049_ ), .Z(_05117_ ) );
NAND4_X1 _12366_ ( .A1(_05093_ ), .A2(fanout_net_7 ), .A3(\EXU.mtvec_i [21] ), .A4(_05094_ ), .ZN(_05118_ ) );
CLKBUF_X2 _12367_ ( .A(_04340_ ), .Z(_05119_ ) );
AND4_X1 _12368_ ( .A1(fanout_net_7 ), .A2(_05053_ ), .A3(\EXU.mepc_i [21] ), .A4(_05119_ ), .ZN(_05120_ ) );
AND4_X1 _12369_ ( .A1(\EXU.pc_i [9] ), .A2(\EXU.pc_i [8] ), .A3(\EXU.pc_i [7] ), .A4(\EXU.pc_i [6] ), .ZN(_05121_ ) );
AND2_X2 _12370_ ( .A1(_05059_ ), .A2(_05121_ ), .ZN(_05122_ ) );
AND4_X1 _12371_ ( .A1(\EXU.pc_i [17] ), .A2(\EXU.pc_i [16] ), .A3(\EXU.pc_i [15] ), .A4(\EXU.pc_i [14] ), .ZN(_05123_ ) );
AND2_X1 _12372_ ( .A1(\EXU.pc_i [11] ), .A2(\EXU.pc_i [10] ), .ZN(_05124_ ) );
AND4_X1 _12373_ ( .A1(\EXU.pc_i [13] ), .A2(_05123_ ), .A3(\EXU.pc_i [12] ), .A4(_05124_ ), .ZN(_05125_ ) );
NAND2_X1 _12374_ ( .A1(_05122_ ), .A2(_05125_ ), .ZN(_05126_ ) );
NOR3_X1 _12375_ ( .A1(_05126_ ), .A2(_04261_ ), .A3(_04262_ ), .ZN(_05127_ ) );
NAND2_X1 _12376_ ( .A1(_05127_ ), .A2(\EXU.pc_i [20] ), .ZN(_05128_ ) );
XNOR2_X1 _12377_ ( .A(_05128_ ), .B(\EXU.pc_i [21] ), .ZN(_05129_ ) );
AOI21_X1 _12378_ ( .A(_05120_ ), .B1(_05129_ ), .B2(_05101_ ), .ZN(_05130_ ) );
OAI21_X1 _12379_ ( .A(_05118_ ), .B1(_05130_ ), .B2(_05104_ ), .ZN(_05131_ ) );
OAI21_X1 _12380_ ( .A(_05116_ ), .B1(_05117_ ), .B2(_05131_ ), .ZN(_05132_ ) );
OAI22_X1 _12381_ ( .A1(_05115_ ), .A2(_05132_ ), .B1(_04251_ ), .B2(_05088_ ), .ZN(_00205_ ) );
XNOR2_X1 _12382_ ( .A(_05111_ ), .B(_04566_ ), .ZN(_05133_ ) );
NOR2_X1 _12383_ ( .A1(_05133_ ), .A2(_05042_ ), .ZN(_05134_ ) );
BUF_X4 _12384_ ( .A(_05082_ ), .Z(_05135_ ) );
NAND4_X1 _12385_ ( .A1(_05093_ ), .A2(fanout_net_7 ), .A3(\EXU.mtvec_i [20] ), .A4(_05094_ ), .ZN(_05136_ ) );
AND4_X1 _12386_ ( .A1(fanout_net_7 ), .A2(_05053_ ), .A3(\EXU.mepc_i [20] ), .A4(_05119_ ), .ZN(_05137_ ) );
AND2_X1 _12387_ ( .A1(_05122_ ), .A2(_05125_ ), .ZN(_05138_ ) );
NAND3_X1 _12388_ ( .A1(_05138_ ), .A2(\EXU.pc_i [19] ), .A3(\EXU.pc_i [18] ), .ZN(_05139_ ) );
XNOR2_X1 _12389_ ( .A(_05139_ ), .B(\EXU.pc_i [20] ), .ZN(_05140_ ) );
AOI21_X1 _12390_ ( .A(_05137_ ), .B1(_05140_ ), .B2(_05101_ ), .ZN(_05141_ ) );
OAI21_X1 _12391_ ( .A(_05136_ ), .B1(_05141_ ), .B2(_05104_ ), .ZN(_05142_ ) );
OAI21_X1 _12392_ ( .A(_05135_ ), .B1(_05117_ ), .B2(_05142_ ), .ZN(_05143_ ) );
OAI22_X1 _12393_ ( .A1(_05134_ ), .A2(_05143_ ), .B1(_04252_ ), .B2(_05088_ ), .ZN(_00206_ ) );
AOI21_X1 _12394_ ( .A(_04589_ ), .B1(_04550_ ), .B2(_04582_ ), .ZN(_05144_ ) );
NOR2_X1 _12395_ ( .A1(_05144_ ), .A2(_04574_ ), .ZN(_05145_ ) );
NOR2_X1 _12396_ ( .A1(_05145_ ), .A2(_04592_ ), .ZN(_05146_ ) );
XNOR2_X1 _12397_ ( .A(_05146_ ), .B(_04570_ ), .ZN(_05147_ ) );
NOR2_X1 _12398_ ( .A1(_05147_ ), .A2(_05042_ ), .ZN(_05148_ ) );
NAND4_X1 _12399_ ( .A1(_05093_ ), .A2(fanout_net_7 ), .A3(\EXU.mtvec_i [19] ), .A4(_05094_ ), .ZN(_05149_ ) );
AND4_X1 _12400_ ( .A1(fanout_net_7 ), .A2(_05053_ ), .A3(\EXU.mepc_i [19] ), .A4(_05119_ ), .ZN(_05150_ ) );
NAND3_X1 _12401_ ( .A1(_05122_ ), .A2(\EXU.pc_i [18] ), .A3(_05125_ ), .ZN(_05151_ ) );
XNOR2_X1 _12402_ ( .A(_05151_ ), .B(\EXU.pc_i [19] ), .ZN(_05152_ ) );
AOI21_X1 _12403_ ( .A(_05150_ ), .B1(_05152_ ), .B2(_05101_ ), .ZN(_05153_ ) );
OAI21_X1 _12404_ ( .A(_05149_ ), .B1(_05153_ ), .B2(_05104_ ), .ZN(_05154_ ) );
OAI21_X1 _12405_ ( .A(_05135_ ), .B1(_05117_ ), .B2(_05154_ ), .ZN(_05155_ ) );
INV_X1 _12406_ ( .A(\EXU.dnpc_o [19] ), .ZN(_05156_ ) );
OAI22_X1 _12407_ ( .A1(_05148_ ), .A2(_05155_ ), .B1(_05156_ ), .B2(_05088_ ), .ZN(_00207_ ) );
XOR2_X1 _12408_ ( .A(_05144_ ), .B(_04574_ ), .Z(_05157_ ) );
NOR2_X1 _12409_ ( .A1(_05157_ ), .A2(_05042_ ), .ZN(_05158_ ) );
NAND4_X1 _12410_ ( .A1(_05092_ ), .A2(fanout_net_7 ), .A3(\EXU.mtvec_i [18] ), .A4(_05094_ ), .ZN(_05159_ ) );
AND4_X1 _12411_ ( .A1(fanout_net_7 ), .A2(_05053_ ), .A3(\EXU.mepc_i [18] ), .A4(_05119_ ), .ZN(_05160_ ) );
XNOR2_X1 _12412_ ( .A(_05126_ ), .B(\EXU.pc_i [18] ), .ZN(_05161_ ) );
AOI21_X1 _12413_ ( .A(_05160_ ), .B1(_05161_ ), .B2(_05101_ ), .ZN(_05162_ ) );
OAI21_X1 _12414_ ( .A(_05159_ ), .B1(_05162_ ), .B2(_05104_ ), .ZN(_05163_ ) );
OAI21_X1 _12415_ ( .A(_05135_ ), .B1(_05117_ ), .B2(_05163_ ), .ZN(_05164_ ) );
INV_X1 _12416_ ( .A(\EXU.dnpc_o [18] ), .ZN(_05165_ ) );
OAI22_X1 _12417_ ( .A1(_05158_ ), .A2(_05164_ ), .B1(_05165_ ), .B2(_05088_ ), .ZN(_00208_ ) );
NAND4_X1 _12418_ ( .A1(_05093_ ), .A2(fanout_net_7 ), .A3(\EXU.mtvec_i [17] ), .A4(_05094_ ), .ZN(_05166_ ) );
AND4_X1 _12419_ ( .A1(fanout_net_7 ), .A2(_05054_ ), .A3(\EXU.mepc_i [17] ), .A4(_05096_ ), .ZN(_05167_ ) );
AND3_X1 _12420_ ( .A1(_05124_ ), .A2(\EXU.pc_i [13] ), .A3(\EXU.pc_i [12] ), .ZN(_05168_ ) );
NAND2_X1 _12421_ ( .A1(_05122_ ), .A2(_05168_ ), .ZN(_05169_ ) );
NOR3_X1 _12422_ ( .A1(_05169_ ), .A2(_04275_ ), .A3(_04276_ ), .ZN(_05170_ ) );
NAND2_X1 _12423_ ( .A1(_05170_ ), .A2(\EXU.pc_i [16] ), .ZN(_05171_ ) );
XNOR2_X1 _12424_ ( .A(_05171_ ), .B(\EXU.pc_i [17] ), .ZN(_05172_ ) );
AOI21_X1 _12425_ ( .A(_05167_ ), .B1(_05172_ ), .B2(_05101_ ), .ZN(_05173_ ) );
OAI21_X1 _12426_ ( .A(_05166_ ), .B1(_05173_ ), .B2(_05104_ ), .ZN(_05174_ ) );
OAI21_X1 _12427_ ( .A(_05116_ ), .B1(_05117_ ), .B2(_05174_ ), .ZN(_05175_ ) );
AND2_X1 _12428_ ( .A1(_04579_ ), .A2(_04586_ ), .ZN(_05176_ ) );
AOI21_X1 _12429_ ( .A(_05176_ ), .B1(_04550_ ), .B2(_04581_ ), .ZN(_05177_ ) );
XNOR2_X1 _12430_ ( .A(_05177_ ), .B(_04578_ ), .ZN(_05178_ ) );
NOR2_X1 _12431_ ( .A1(_05178_ ), .A2(_05091_ ), .ZN(_05179_ ) );
OAI22_X1 _12432_ ( .A1(_05175_ ), .A2(_05179_ ), .B1(_04242_ ), .B2(_05088_ ), .ZN(_00209_ ) );
NAND4_X1 _12433_ ( .A1(_05093_ ), .A2(fanout_net_7 ), .A3(\EXU.mtvec_i [16] ), .A4(_05094_ ), .ZN(_05180_ ) );
AND4_X1 _12434_ ( .A1(fanout_net_7 ), .A2(_05054_ ), .A3(\EXU.mepc_i [16] ), .A4(_05119_ ), .ZN(_05181_ ) );
INV_X1 _12435_ ( .A(\EXU.pc_i [16] ), .ZN(_05182_ ) );
XNOR2_X1 _12436_ ( .A(_05170_ ), .B(_05182_ ), .ZN(_05183_ ) );
AOI21_X1 _12437_ ( .A(_05181_ ), .B1(_05183_ ), .B2(_05101_ ), .ZN(_05184_ ) );
OAI21_X1 _12438_ ( .A(_05180_ ), .B1(_05184_ ), .B2(_05104_ ), .ZN(_05185_ ) );
OAI21_X1 _12439_ ( .A(_05116_ ), .B1(_05117_ ), .B2(_05185_ ), .ZN(_05186_ ) );
XNOR2_X1 _12440_ ( .A(_04549_ ), .B(_04581_ ), .ZN(_05187_ ) );
INV_X1 _12441_ ( .A(_05034_ ), .ZN(_05188_ ) );
BUF_X2 _12442_ ( .A(_05037_ ), .Z(_05189_ ) );
AOI21_X1 _12443_ ( .A(_05187_ ), .B1(_05188_ ), .B2(_05189_ ), .ZN(_05190_ ) );
OAI22_X1 _12444_ ( .A1(_05186_ ), .A2(_05190_ ), .B1(_04243_ ), .B2(_05088_ ), .ZN(_00210_ ) );
NAND2_X1 _12445_ ( .A1(_04493_ ), .A2(_04526_ ), .ZN(_05191_ ) );
AND2_X1 _12446_ ( .A1(_04533_ ), .A2(_04538_ ), .ZN(_05192_ ) );
AND2_X1 _12447_ ( .A1(_05191_ ), .A2(_05192_ ), .ZN(_05193_ ) );
INV_X1 _12448_ ( .A(_05193_ ), .ZN(_05194_ ) );
AOI21_X1 _12449_ ( .A(_04545_ ), .B1(_05194_ ), .B2(_04510_ ), .ZN(_05195_ ) );
XOR2_X1 _12450_ ( .A(_04494_ ), .B(_04496_ ), .Z(_05196_ ) );
OAI21_X1 _12451_ ( .A(_04498_ ), .B1(_05195_ ), .B2(_05196_ ), .ZN(_05197_ ) );
XOR2_X1 _12452_ ( .A(_05197_ ), .B(_04501_ ), .Z(_05198_ ) );
NOR2_X1 _12453_ ( .A1(_05198_ ), .A2(_05042_ ), .ZN(_05199_ ) );
NAND4_X1 _12454_ ( .A1(_05092_ ), .A2(fanout_net_7 ), .A3(\EXU.mtvec_i [15] ), .A4(_05055_ ), .ZN(_05200_ ) );
AND4_X1 _12455_ ( .A1(fanout_net_7 ), .A2(_05053_ ), .A3(\EXU.mepc_i [15] ), .A4(_05119_ ), .ZN(_05201_ ) );
NAND3_X1 _12456_ ( .A1(_05122_ ), .A2(\EXU.pc_i [14] ), .A3(_05168_ ), .ZN(_05202_ ) );
XNOR2_X1 _12457_ ( .A(_05202_ ), .B(\EXU.pc_i [15] ), .ZN(_05203_ ) );
AOI21_X1 _12458_ ( .A(_05201_ ), .B1(_05203_ ), .B2(_05101_ ), .ZN(_05204_ ) );
OAI21_X1 _12459_ ( .A(_05200_ ), .B1(_05204_ ), .B2(_05103_ ), .ZN(_05205_ ) );
OAI21_X1 _12460_ ( .A(_05135_ ), .B1(_05117_ ), .B2(_05205_ ), .ZN(_05206_ ) );
INV_X1 _12461_ ( .A(\EXU.dnpc_o [15] ), .ZN(_05207_ ) );
BUF_X4 _12462_ ( .A(_05087_ ), .Z(_05208_ ) );
OAI22_X1 _12463_ ( .A1(_05199_ ), .A2(_05206_ ), .B1(_05207_ ), .B2(_05208_ ), .ZN(_00211_ ) );
XOR2_X1 _12464_ ( .A(_05195_ ), .B(_05196_ ), .Z(_05209_ ) );
NOR2_X1 _12465_ ( .A1(_05209_ ), .A2(_05040_ ), .ZN(_05210_ ) );
BUF_X4 _12466_ ( .A(_05039_ ), .Z(_05211_ ) );
AND4_X1 _12467_ ( .A1(fanout_net_7 ), .A2(_05047_ ), .A3(\EXU.mtvec_i [14] ), .A4(_04340_ ), .ZN(_05212_ ) );
OAI21_X1 _12468_ ( .A(_04360_ ), .B1(_05099_ ), .B2(\EXU.mepc_i [14] ), .ZN(_05213_ ) );
XNOR2_X1 _12469_ ( .A(_05169_ ), .B(_04276_ ), .ZN(_05214_ ) );
AOI21_X1 _12470_ ( .A(_05213_ ), .B1(_05214_ ), .B2(_05100_ ), .ZN(_05215_ ) );
NOR4_X1 _12471_ ( .A1(_05034_ ), .A2(_05211_ ), .A3(_05212_ ), .A4(_05215_ ), .ZN(_05216_ ) );
OR3_X1 _12472_ ( .A1(_05210_ ), .A2(_05083_ ), .A3(_05216_ ), .ZN(_05217_ ) );
INV_X1 _12473_ ( .A(\EXU.dnpc_o [14] ), .ZN(_05218_ ) );
OAI21_X1 _12474_ ( .A(_05217_ ), .B1(_05218_ ), .B2(_05088_ ), .ZN(_00212_ ) );
NAND4_X1 _12475_ ( .A1(_05054_ ), .A2(fanout_net_7 ), .A3(\EXU.mepc_i [13] ), .A4(_05096_ ), .ZN(_05219_ ) );
NAND3_X1 _12476_ ( .A1(_05059_ ), .A2(_05121_ ), .A3(_05124_ ), .ZN(_05220_ ) );
NOR2_X1 _12477_ ( .A1(_05220_ ), .A2(_04278_ ), .ZN(_05221_ ) );
XNOR2_X1 _12478_ ( .A(_05221_ ), .B(\EXU.pc_i [13] ), .ZN(_05222_ ) );
OAI21_X1 _12479_ ( .A(_05219_ ), .B1(_05222_ ), .B2(_05077_ ), .ZN(_05223_ ) );
MUX2_X1 _12480_ ( .A(\EXU.mtvec_i [13] ), .B(_05223_ ), .S(_05050_ ), .Z(_05224_ ) );
OAI21_X1 _12481_ ( .A(_05116_ ), .B1(_05117_ ), .B2(_05224_ ), .ZN(_05225_ ) );
AND2_X1 _12482_ ( .A1(_04507_ ), .A2(_04542_ ), .ZN(_05226_ ) );
AOI21_X1 _12483_ ( .A(_05226_ ), .B1(_05194_ ), .B2(_04509_ ), .ZN(_05227_ ) );
XNOR2_X1 _12484_ ( .A(_05227_ ), .B(_04506_ ), .ZN(_05228_ ) );
NOR2_X1 _12485_ ( .A1(_05228_ ), .A2(_05091_ ), .ZN(_05229_ ) );
OAI22_X1 _12486_ ( .A1(_05225_ ), .A2(_05229_ ), .B1(_04226_ ), .B2(_05208_ ), .ZN(_00213_ ) );
NAND4_X1 _12487_ ( .A1(_05093_ ), .A2(fanout_net_7 ), .A3(\EXU.mtvec_i [12] ), .A4(_05094_ ), .ZN(_05230_ ) );
AND4_X1 _12488_ ( .A1(fanout_net_7 ), .A2(_05054_ ), .A3(\EXU.mepc_i [12] ), .A4(_05119_ ), .ZN(_05231_ ) );
XNOR2_X1 _12489_ ( .A(_05220_ ), .B(\EXU.pc_i [12] ), .ZN(_05232_ ) );
AOI21_X1 _12490_ ( .A(_05231_ ), .B1(_05232_ ), .B2(_05101_ ), .ZN(_05233_ ) );
OAI21_X1 _12491_ ( .A(_05230_ ), .B1(_05233_ ), .B2(_05104_ ), .ZN(_05234_ ) );
OAI21_X1 _12492_ ( .A(_05116_ ), .B1(_05117_ ), .B2(_05234_ ), .ZN(_05235_ ) );
XNOR2_X1 _12493_ ( .A(_05193_ ), .B(_04509_ ), .ZN(_05236_ ) );
AOI21_X1 _12494_ ( .A(_05236_ ), .B1(_05188_ ), .B2(_05189_ ), .ZN(_05237_ ) );
OAI22_X1 _12495_ ( .A1(_05235_ ), .A2(_05237_ ), .B1(_04227_ ), .B2(_05208_ ), .ZN(_00214_ ) );
NAND3_X1 _12496_ ( .A1(_05045_ ), .A2(\EXU.mtvec_i [29] ), .A3(_05093_ ), .ZN(_05238_ ) );
AND4_X1 _12497_ ( .A1(fanout_net_7 ), .A2(_05054_ ), .A3(\EXU.mepc_i [29] ), .A4(_05119_ ), .ZN(_05239_ ) );
NAND4_X1 _12498_ ( .A1(\EXU.pc_i [25] ), .A2(\EXU.pc_i [24] ), .A3(\EXU.pc_i [23] ), .A4(\EXU.pc_i [22] ), .ZN(_05240_ ) );
NAND2_X1 _12499_ ( .A1(\EXU.pc_i [21] ), .A2(\EXU.pc_i [20] ), .ZN(_05241_ ) );
NOR4_X1 _12500_ ( .A1(_05240_ ), .A2(_05241_ ), .A3(_04261_ ), .A4(_04262_ ), .ZN(_05242_ ) );
AND2_X1 _12501_ ( .A1(_05138_ ), .A2(_05242_ ), .ZN(_05243_ ) );
AND3_X1 _12502_ ( .A1(_05243_ ), .A2(\EXU.pc_i [27] ), .A3(\EXU.pc_i [26] ), .ZN(_05244_ ) );
NAND2_X1 _12503_ ( .A1(_05244_ ), .A2(\EXU.pc_i [28] ), .ZN(_05245_ ) );
XNOR2_X1 _12504_ ( .A(_05245_ ), .B(\EXU.pc_i [29] ), .ZN(_05246_ ) );
AOI21_X1 _12505_ ( .A(_05239_ ), .B1(_05246_ ), .B2(_05101_ ), .ZN(_05247_ ) );
OAI211_X1 _12506_ ( .A(_05041_ ), .B(_05238_ ), .C1(_05104_ ), .C2(_05247_ ), .ZN(_05248_ ) );
AOI21_X1 _12507_ ( .A(_04640_ ), .B1(_04632_ ), .B2(_04641_ ), .ZN(_05249_ ) );
XNOR2_X1 _12508_ ( .A(_05249_ ), .B(_04635_ ), .ZN(_05250_ ) );
OAI211_X1 _12509_ ( .A(_05116_ ), .B(_05248_ ), .C1(_05250_ ), .C2(_05091_ ), .ZN(_05251_ ) );
BUF_X2 _12510_ ( .A(_05080_ ), .Z(_05252_ ) );
INV_X1 _12511_ ( .A(_04393_ ), .ZN(_05253_ ) );
OAI211_X1 _12512_ ( .A(\EXU.dnpc_o [29] ), .B(_05252_ ), .C1(_05253_ ), .C2(\LSU.ls_read_done_$_OR__B_Y_$_ORNOT__A_Y_$_ANDNOT__A_Y_$_OR__A_1_B ), .ZN(_05254_ ) );
NAND2_X1 _12513_ ( .A1(_05251_ ), .A2(_05254_ ), .ZN(_00215_ ) );
AOI21_X1 _12514_ ( .A(_04532_ ), .B1(_04493_ ), .B2(_04525_ ), .ZN(_05255_ ) );
NOR2_X1 _12515_ ( .A1(_05255_ ), .A2(_04517_ ), .ZN(_05256_ ) );
OR2_X1 _12516_ ( .A1(_05256_ ), .A2(_04535_ ), .ZN(_05257_ ) );
XNOR2_X1 _12517_ ( .A(_05257_ ), .B(_04514_ ), .ZN(_05258_ ) );
NOR2_X1 _12518_ ( .A1(_05042_ ), .A2(_05258_ ), .ZN(_05259_ ) );
AND4_X1 _12519_ ( .A1(fanout_net_7 ), .A2(_05047_ ), .A3(\EXU.mtvec_i [11] ), .A4(_05096_ ), .ZN(_05260_ ) );
NAND3_X1 _12520_ ( .A1(_05059_ ), .A2(\EXU.pc_i [10] ), .A3(_05121_ ), .ZN(_05261_ ) );
XNOR2_X1 _12521_ ( .A(_05261_ ), .B(\EXU.pc_i [11] ), .ZN(_05262_ ) );
MUX2_X1 _12522_ ( .A(\EXU.mepc_i [11] ), .B(_05262_ ), .S(_05099_ ), .Z(_05263_ ) );
BUF_X4 _12523_ ( .A(_05050_ ), .Z(_05264_ ) );
AOI21_X1 _12524_ ( .A(_05260_ ), .B1(_05263_ ), .B2(_05264_ ), .ZN(_05265_ ) );
OAI211_X1 _12525_ ( .A(_05189_ ), .B(_05265_ ), .C1(_05033_ ), .C2(_04961_ ), .ZN(_05266_ ) );
NAND2_X1 _12526_ ( .A1(_05266_ ), .A2(_05116_ ), .ZN(_05267_ ) );
INV_X1 _12527_ ( .A(\EXU.dnpc_o [11] ), .ZN(_05268_ ) );
OAI22_X1 _12528_ ( .A1(_05259_ ), .A2(_05267_ ), .B1(_05268_ ), .B2(_05208_ ), .ZN(_00216_ ) );
XOR2_X1 _12529_ ( .A(_05255_ ), .B(_04517_ ), .Z(_05269_ ) );
INV_X1 _12530_ ( .A(_05269_ ), .ZN(_05270_ ) );
AND4_X1 _12531_ ( .A1(fanout_net_7 ), .A2(_05047_ ), .A3(\EXU.mtvec_i [10] ), .A4(_05096_ ), .ZN(_05271_ ) );
XNOR2_X1 _12532_ ( .A(_05122_ ), .B(_04281_ ), .ZN(_05272_ ) );
MUX2_X1 _12533_ ( .A(\EXU.mepc_i [10] ), .B(_05272_ ), .S(_05100_ ), .Z(_05273_ ) );
AOI21_X1 _12534_ ( .A(_05271_ ), .B1(_05273_ ), .B2(_05264_ ), .ZN(_05274_ ) );
MUX2_X1 _12535_ ( .A(_05270_ ), .B(_05274_ ), .S(_05041_ ), .Z(_05275_ ) );
INV_X1 _12536_ ( .A(\EXU.dnpc_o [10] ), .ZN(_05276_ ) );
OAI22_X1 _12537_ ( .A1(_05275_ ), .A2(_05083_ ), .B1(_05276_ ), .B2(_05208_ ), .ZN(_00217_ ) );
NAND2_X1 _12538_ ( .A1(_04493_ ), .A2(_04524_ ), .ZN(_05277_ ) );
NAND2_X1 _12539_ ( .A1(_04522_ ), .A2(_04529_ ), .ZN(_05278_ ) );
NAND2_X1 _12540_ ( .A1(_05277_ ), .A2(_05278_ ), .ZN(_05279_ ) );
XOR2_X1 _12541_ ( .A(_05279_ ), .B(_04521_ ), .Z(_05280_ ) );
OAI21_X1 _12542_ ( .A(_05116_ ), .B1(_05091_ ), .B2(_05280_ ), .ZN(_05281_ ) );
AND4_X1 _12543_ ( .A1(fanout_net_7 ), .A2(_05092_ ), .A3(\EXU.mtvec_i [9] ), .A4(_05096_ ), .ZN(_05282_ ) );
AND2_X1 _12544_ ( .A1(_05061_ ), .A2(\EXU.pc_i [8] ), .ZN(_05283_ ) );
XNOR2_X1 _12545_ ( .A(_05283_ ), .B(_04282_ ), .ZN(_05284_ ) );
MUX2_X1 _12546_ ( .A(\EXU.mepc_i [9] ), .B(_05284_ ), .S(_05100_ ), .Z(_05285_ ) );
AOI21_X1 _12547_ ( .A(_05282_ ), .B1(_05285_ ), .B2(_05051_ ), .ZN(_05286_ ) );
AND3_X1 _12548_ ( .A1(_05188_ ), .A2(_05189_ ), .A3(_05286_ ), .ZN(_05287_ ) );
INV_X1 _12549_ ( .A(\EXU.dnpc_o [9] ), .ZN(_05288_ ) );
OAI22_X1 _12550_ ( .A1(_05281_ ), .A2(_05287_ ), .B1(_05288_ ), .B2(_05208_ ), .ZN(_00218_ ) );
NAND4_X1 _12551_ ( .A1(_05093_ ), .A2(\EXU.op_i [4] ), .A3(\EXU.mtvec_i [8] ), .A4(_05094_ ), .ZN(_05289_ ) );
BUF_X4 _12552_ ( .A(_05050_ ), .Z(_05290_ ) );
OR2_X1 _12553_ ( .A1(_05100_ ), .A2(\EXU.mepc_i [8] ), .ZN(_05291_ ) );
XNOR2_X1 _12554_ ( .A(_05061_ ), .B(_04283_ ), .ZN(_05292_ ) );
OAI211_X1 _12555_ ( .A(_05290_ ), .B(_05291_ ), .C1(_05292_ ), .C2(_05077_ ), .ZN(_05293_ ) );
AND4_X1 _12556_ ( .A1(_05189_ ), .A2(_05188_ ), .A3(_05289_ ), .A4(_05293_ ), .ZN(_05294_ ) );
XOR2_X1 _12557_ ( .A(_04493_ ), .B(_04524_ ), .Z(_05295_ ) );
OAI21_X1 _12558_ ( .A(_05135_ ), .B1(_05091_ ), .B2(_05295_ ), .ZN(_05296_ ) );
INV_X1 _12559_ ( .A(\EXU.dnpc_o [8] ), .ZN(_05297_ ) );
OAI22_X1 _12560_ ( .A1(_05294_ ), .A2(_05296_ ), .B1(_05297_ ), .B2(_05208_ ), .ZN(_00219_ ) );
NAND4_X1 _12561_ ( .A1(_05093_ ), .A2(\EXU.op_i [4] ), .A3(\EXU.mtvec_i [7] ), .A4(_05094_ ), .ZN(_05298_ ) );
OR2_X1 _12562_ ( .A1(_05100_ ), .A2(\EXU.mepc_i [7] ), .ZN(_05299_ ) );
XNOR2_X1 _12563_ ( .A(_05060_ ), .B(_04270_ ), .ZN(_05300_ ) );
OAI211_X1 _12564_ ( .A(_05290_ ), .B(_05299_ ), .C1(_05300_ ), .C2(_05077_ ), .ZN(_05301_ ) );
AND4_X1 _12565_ ( .A1(_05189_ ), .A2(_05188_ ), .A3(_05298_ ), .A4(_05301_ ), .ZN(_05302_ ) );
XOR2_X1 _12566_ ( .A(_04485_ ), .B(_04489_ ), .Z(_05303_ ) );
OAI21_X1 _12567_ ( .A(_05135_ ), .B1(_05091_ ), .B2(_05303_ ), .ZN(_05304_ ) );
OAI22_X1 _12568_ ( .A1(_05302_ ), .A2(_05304_ ), .B1(_04235_ ), .B2(_05208_ ), .ZN(_00220_ ) );
AOI21_X1 _12569_ ( .A(_04480_ ), .B1(_04481_ ), .B2(_04477_ ), .ZN(_05305_ ) );
XNOR2_X1 _12570_ ( .A(_05305_ ), .B(_04444_ ), .ZN(_05306_ ) );
OAI21_X1 _12571_ ( .A(_05116_ ), .B1(_05091_ ), .B2(_05306_ ), .ZN(_05307_ ) );
AND4_X1 _12572_ ( .A1(\EXU.op_i [4] ), .A2(_05047_ ), .A3(\EXU.mtvec_i [6] ), .A4(_05096_ ), .ZN(_05308_ ) );
XNOR2_X1 _12573_ ( .A(_05059_ ), .B(_04271_ ), .ZN(_05309_ ) );
MUX2_X1 _12574_ ( .A(_05309_ ), .B(\EXU.mepc_i [6] ), .S(_05077_ ), .Z(_05310_ ) );
AOI21_X1 _12575_ ( .A(_05308_ ), .B1(_05310_ ), .B2(_05051_ ), .ZN(_05311_ ) );
AND3_X1 _12576_ ( .A1(_05188_ ), .A2(_05189_ ), .A3(_05311_ ), .ZN(_05312_ ) );
OAI22_X1 _12577_ ( .A1(_05307_ ), .A2(_05312_ ), .B1(_04236_ ), .B2(_05208_ ), .ZN(_00221_ ) );
XOR2_X1 _12578_ ( .A(_04476_ ), .B(_04479_ ), .Z(_05313_ ) );
OAI21_X1 _12579_ ( .A(_05116_ ), .B1(_05091_ ), .B2(_05313_ ), .ZN(_05314_ ) );
AND4_X1 _12580_ ( .A1(\EXU.op_i [4] ), .A2(_05047_ ), .A3(\EXU.mtvec_i [5] ), .A4(_05096_ ), .ZN(_05315_ ) );
NAND4_X1 _12581_ ( .A1(_05054_ ), .A2(\EXU.op_i [4] ), .A3(\EXU.mepc_i [5] ), .A4(_05055_ ), .ZN(_05316_ ) );
XNOR2_X1 _12582_ ( .A(_05058_ ), .B(_04272_ ), .ZN(_05317_ ) );
INV_X1 _12583_ ( .A(_05317_ ), .ZN(_05318_ ) );
OAI21_X1 _12584_ ( .A(_05316_ ), .B1(_05318_ ), .B2(_05077_ ), .ZN(_05319_ ) );
AOI21_X1 _12585_ ( .A(_05315_ ), .B1(_05319_ ), .B2(_05051_ ), .ZN(_05320_ ) );
AND3_X1 _12586_ ( .A1(_05188_ ), .A2(_05189_ ), .A3(_05320_ ), .ZN(_05321_ ) );
OAI22_X1 _12587_ ( .A1(_05314_ ), .A2(_05321_ ), .B1(_04237_ ), .B2(_05208_ ), .ZN(_00222_ ) );
NAND4_X1 _12588_ ( .A1(_05054_ ), .A2(\EXU.op_i [4] ), .A3(\EXU.mepc_i [4] ), .A4(_05055_ ), .ZN(_05322_ ) );
XNOR2_X1 _12589_ ( .A(_05057_ ), .B(_04273_ ), .ZN(_05323_ ) );
INV_X1 _12590_ ( .A(_05323_ ), .ZN(_05324_ ) );
OAI211_X1 _12591_ ( .A(_05051_ ), .B(_05322_ ), .C1(_05077_ ), .C2(_05324_ ), .ZN(_05325_ ) );
OR2_X1 _12592_ ( .A1(_05051_ ), .A2(\EXU.mtvec_i [4] ), .ZN(_05326_ ) );
AOI211_X1 _12593_ ( .A(_05211_ ), .B(_05034_ ), .C1(_05325_ ), .C2(_05326_ ), .ZN(_05327_ ) );
XNOR2_X1 _12594_ ( .A(_04445_ ), .B(_04447_ ), .ZN(_05328_ ) );
XNOR2_X1 _12595_ ( .A(_04474_ ), .B(_05328_ ), .ZN(_05329_ ) );
OAI21_X1 _12596_ ( .A(_05135_ ), .B1(_05041_ ), .B2(_05329_ ), .ZN(_05330_ ) );
BUF_X4 _12597_ ( .A(_05087_ ), .Z(_05331_ ) );
OAI22_X1 _12598_ ( .A1(_05327_ ), .A2(_05330_ ), .B1(_04238_ ), .B2(_05331_ ), .ZN(_00223_ ) );
NAND4_X1 _12599_ ( .A1(_05054_ ), .A2(\EXU.op_i [4] ), .A3(\EXU.mepc_i [3] ), .A4(_05055_ ), .ZN(_05332_ ) );
XOR2_X1 _12600_ ( .A(\EXU.pc_i [3] ), .B(\EXU.pc_i [2] ), .Z(_05333_ ) );
INV_X1 _12601_ ( .A(_05333_ ), .ZN(_05334_ ) );
OAI211_X1 _12602_ ( .A(_05051_ ), .B(_05332_ ), .C1(_05077_ ), .C2(_05334_ ), .ZN(_05335_ ) );
OR2_X1 _12603_ ( .A1(_05051_ ), .A2(\EXU.mtvec_i [3] ), .ZN(_05336_ ) );
AOI211_X1 _12604_ ( .A(_05211_ ), .B(_05034_ ), .C1(_05335_ ), .C2(_05336_ ), .ZN(_05337_ ) );
XNOR2_X1 _12605_ ( .A(_04466_ ), .B(_04470_ ), .ZN(_05338_ ) );
OAI21_X1 _12606_ ( .A(_05135_ ), .B1(_05041_ ), .B2(_05338_ ), .ZN(_05339_ ) );
OAI22_X1 _12607_ ( .A1(_05337_ ), .A2(_05339_ ), .B1(_04230_ ), .B2(_05331_ ), .ZN(_00224_ ) );
AND4_X1 _12608_ ( .A1(\EXU.op_i [4] ), .A2(_05092_ ), .A3(\EXU.mtvec_i [2] ), .A4(_05055_ ), .ZN(_05340_ ) );
MUX2_X1 _12609_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_B_$_MUX__Y_B ), .B(\EXU.mepc_i [2] ), .S(_05077_ ), .Z(_05341_ ) );
AOI211_X1 _12610_ ( .A(_05340_ ), .B(_05049_ ), .C1(_05051_ ), .C2(_05341_ ), .ZN(_05342_ ) );
XOR2_X1 _12611_ ( .A(_04457_ ), .B(_04464_ ), .Z(_05343_ ) );
OAI21_X1 _12612_ ( .A(_05135_ ), .B1(_05041_ ), .B2(_05343_ ), .ZN(_05344_ ) );
OAI22_X1 _12613_ ( .A1(_05342_ ), .A2(_05344_ ), .B1(_04231_ ), .B2(_05331_ ), .ZN(_00225_ ) );
XNOR2_X1 _12614_ ( .A(_04631_ ), .B(_04641_ ), .ZN(_05345_ ) );
AND2_X1 _12615_ ( .A1(_05345_ ), .A2(_05049_ ), .ZN(_05346_ ) );
XOR2_X1 _12616_ ( .A(_05244_ ), .B(\EXU.pc_i [28] ), .Z(_05347_ ) );
MUX2_X1 _12617_ ( .A(\EXU.mepc_i [28] ), .B(_05347_ ), .S(_05099_ ), .Z(_05348_ ) );
MUX2_X1 _12618_ ( .A(\EXU.mtvec_i [28] ), .B(_05348_ ), .S(_04360_ ), .Z(_05349_ ) );
AOI21_X1 _12619_ ( .A(_05346_ ), .B1(_05040_ ), .B2(_05349_ ), .ZN(_05350_ ) );
NOR3_X1 _12620_ ( .A1(_05350_ ), .A2(\LSU.ls_read_done_$_OR__B_Y_$_ORNOT__A_Y_$_ANDNOT__A_Y_$_OR__A_1_B ), .A3(_05086_ ), .ZN(_05351_ ) );
MUX2_X1 _12621_ ( .A(\EXU.dnpc_o [28] ), .B(_05351_ ), .S(_05087_ ), .Z(_00226_ ) );
XOR2_X1 _12622_ ( .A(_04453_ ), .B(_04456_ ), .Z(_05352_ ) );
BUF_X2 _12623_ ( .A(_05352_ ), .Z(_05353_ ) );
INV_X1 _12624_ ( .A(_05353_ ), .ZN(_05354_ ) );
AND4_X1 _12625_ ( .A1(\EXU.op_i [4] ), .A2(_05047_ ), .A3(\EXU.mtvec_i [1] ), .A4(_05096_ ), .ZN(_05355_ ) );
MUX2_X1 _12626_ ( .A(\EXU.add_pc_4 [1] ), .B(\EXU.mepc_i [1] ), .S(_05076_ ), .Z(_05356_ ) );
AOI21_X1 _12627_ ( .A(_05355_ ), .B1(_05356_ ), .B2(_05264_ ), .ZN(_05357_ ) );
MUX2_X1 _12628_ ( .A(_05354_ ), .B(_05357_ ), .S(_05041_ ), .Z(_05358_ ) );
OAI22_X1 _12629_ ( .A1(_05358_ ), .A2(_05083_ ), .B1(_04232_ ), .B2(_05331_ ), .ZN(_00227_ ) );
XOR2_X1 _12630_ ( .A(_04454_ ), .B(_04455_ ), .Z(_05359_ ) );
AND2_X1 _12631_ ( .A1(_05359_ ), .A2(_05036_ ), .ZN(_05360_ ) );
INV_X2 _12632_ ( .A(_05359_ ), .ZN(_05361_ ) );
AOI21_X1 _12633_ ( .A(_05211_ ), .B1(_05034_ ), .B2(_05361_ ), .ZN(_05362_ ) );
INV_X1 _12634_ ( .A(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_A ), .ZN(_05363_ ) );
NAND4_X1 _12635_ ( .A1(_05092_ ), .A2(\EXU.op_i [4] ), .A3(_05363_ ), .A4(_05055_ ), .ZN(_05364_ ) );
MUX2_X1 _12636_ ( .A(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_B ), .B(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_B_$_MUX__A_B ), .S(_05077_ ), .Z(_05365_ ) );
OAI221_X1 _12637_ ( .A(_05364_ ), .B1(_05103_ ), .B2(_05365_ ), .C1(_05033_ ), .C2(_04961_ ), .ZN(_05366_ ) );
AOI21_X1 _12638_ ( .A(_05360_ ), .B1(_05362_ ), .B2(_05366_ ), .ZN(_05367_ ) );
OAI22_X1 _12639_ ( .A1(_05367_ ), .A2(_05083_ ), .B1(_04233_ ), .B2(_05331_ ), .ZN(_00228_ ) );
AOI21_X1 _12640_ ( .A(_04629_ ), .B1(_04606_ ), .B2(_04622_ ), .ZN(_05368_ ) );
OAI21_X1 _12641_ ( .A(_04624_ ), .B1(_05368_ ), .B2(_04610_ ), .ZN(_05369_ ) );
XNOR2_X1 _12642_ ( .A(_05369_ ), .B(_04614_ ), .ZN(_05370_ ) );
AND2_X1 _12643_ ( .A1(_05370_ ), .A2(_05049_ ), .ZN(_05371_ ) );
NAND3_X1 _12644_ ( .A1(_05138_ ), .A2(\EXU.pc_i [26] ), .A3(_05242_ ), .ZN(_05372_ ) );
XNOR2_X1 _12645_ ( .A(_05372_ ), .B(\EXU.pc_i [27] ), .ZN(_05373_ ) );
MUX2_X1 _12646_ ( .A(\EXU.mepc_i [27] ), .B(_05373_ ), .S(_05099_ ), .Z(_05374_ ) );
MUX2_X1 _12647_ ( .A(\EXU.mtvec_i [27] ), .B(_05374_ ), .S(_05050_ ), .Z(_05375_ ) );
AOI21_X1 _12648_ ( .A(_05371_ ), .B1(_05091_ ), .B2(_05375_ ), .ZN(_05376_ ) );
OAI22_X1 _12649_ ( .A1(_05376_ ), .A2(_05083_ ), .B1(_04246_ ), .B2(_05331_ ), .ZN(_00229_ ) );
NAND3_X1 _12650_ ( .A1(_05045_ ), .A2(\EXU.mtvec_i [26] ), .A3(_05092_ ), .ZN(_05377_ ) );
AND4_X1 _12651_ ( .A1(\EXU.op_i [4] ), .A2(_05053_ ), .A3(\EXU.mepc_i [26] ), .A4(_04340_ ), .ZN(_05378_ ) );
XOR2_X1 _12652_ ( .A(_05243_ ), .B(\EXU.pc_i [26] ), .Z(_05379_ ) );
AOI21_X1 _12653_ ( .A(_05378_ ), .B1(_05379_ ), .B2(_05100_ ), .ZN(_05380_ ) );
OAI211_X1 _12654_ ( .A(_05041_ ), .B(_05377_ ), .C1(_05104_ ), .C2(_05380_ ), .ZN(_05381_ ) );
XOR2_X1 _12655_ ( .A(_05368_ ), .B(_04610_ ), .Z(_05382_ ) );
OAI211_X1 _12656_ ( .A(_05082_ ), .B(_05381_ ), .C1(_05382_ ), .C2(_05041_ ), .ZN(_05383_ ) );
OAI21_X1 _12657_ ( .A(_05383_ ), .B1(_04247_ ), .B2(_05088_ ), .ZN(_00230_ ) );
AND4_X1 _12658_ ( .A1(\EXU.op_i [4] ), .A2(_05047_ ), .A3(\EXU.mtvec_i [25] ), .A4(_05096_ ), .ZN(_05384_ ) );
NOR3_X1 _12659_ ( .A1(_05241_ ), .A2(_04261_ ), .A3(_04262_ ), .ZN(_05385_ ) );
AND2_X1 _12660_ ( .A1(_05138_ ), .A2(_05385_ ), .ZN(_05386_ ) );
AND3_X1 _12661_ ( .A1(_05386_ ), .A2(\EXU.pc_i [23] ), .A3(\EXU.pc_i [22] ), .ZN(_05387_ ) );
NAND2_X1 _12662_ ( .A1(_05387_ ), .A2(\EXU.pc_i [24] ), .ZN(_05388_ ) );
XNOR2_X1 _12663_ ( .A(_05388_ ), .B(\EXU.pc_i [25] ), .ZN(_05389_ ) );
MUX2_X1 _12664_ ( .A(\EXU.mepc_i [25] ), .B(_05389_ ), .S(_05100_ ), .Z(_05390_ ) );
AOI21_X1 _12665_ ( .A(_05384_ ), .B1(_05390_ ), .B2(_05264_ ), .ZN(_05391_ ) );
AND2_X1 _12666_ ( .A1(_04619_ ), .A2(_04626_ ), .ZN(_05392_ ) );
AOI21_X1 _12667_ ( .A(_05392_ ), .B1(_04606_ ), .B2(_04621_ ), .ZN(_05393_ ) );
XOR2_X1 _12668_ ( .A(_05393_ ), .B(_04618_ ), .Z(_05394_ ) );
MUX2_X1 _12669_ ( .A(_05391_ ), .B(_05394_ ), .S(_05049_ ), .Z(_05395_ ) );
OAI22_X1 _12670_ ( .A1(_05395_ ), .A2(_05083_ ), .B1(_04248_ ), .B2(_05331_ ), .ZN(_00231_ ) );
XNOR2_X1 _12671_ ( .A(_04605_ ), .B(_04621_ ), .ZN(_05396_ ) );
NOR2_X1 _12672_ ( .A1(_05396_ ), .A2(_05042_ ), .ZN(_05397_ ) );
NAND4_X1 _12673_ ( .A1(_05092_ ), .A2(\EXU.op_i [4] ), .A3(\EXU.mtvec_i [24] ), .A4(_05055_ ), .ZN(_05398_ ) );
AND4_X1 _12674_ ( .A1(\EXU.op_i [4] ), .A2(_05053_ ), .A3(\EXU.mepc_i [24] ), .A4(_05119_ ), .ZN(_05399_ ) );
NAND3_X1 _12675_ ( .A1(_05386_ ), .A2(\EXU.pc_i [23] ), .A3(\EXU.pc_i [22] ), .ZN(_05400_ ) );
XNOR2_X1 _12676_ ( .A(_05400_ ), .B(\EXU.pc_i [24] ), .ZN(_05401_ ) );
AOI21_X1 _12677_ ( .A(_05399_ ), .B1(_05401_ ), .B2(_05100_ ), .ZN(_05402_ ) );
OAI21_X1 _12678_ ( .A(_05398_ ), .B1(_05402_ ), .B2(_05103_ ), .ZN(_05403_ ) );
OAI21_X1 _12679_ ( .A(_05135_ ), .B1(_05117_ ), .B2(_05403_ ), .ZN(_05404_ ) );
OAI22_X1 _12680_ ( .A1(_05397_ ), .A2(_05404_ ), .B1(_04249_ ), .B2(_05331_ ), .ZN(_00232_ ) );
AOI21_X1 _12681_ ( .A(_04600_ ), .B1(_05112_ ), .B2(_04567_ ), .ZN(_05405_ ) );
OR2_X1 _12682_ ( .A1(_05405_ ), .A2(_04553_ ), .ZN(_05406_ ) );
OAI21_X1 _12683_ ( .A(_05406_ ), .B1(_04552_ ), .B2(_04602_ ), .ZN(_05407_ ) );
XNOR2_X1 _12684_ ( .A(_04555_ ), .B(_04556_ ), .ZN(_05408_ ) );
XOR2_X1 _12685_ ( .A(_05407_ ), .B(_05408_ ), .Z(_05409_ ) );
NOR2_X1 _12686_ ( .A1(_05409_ ), .A2(_05042_ ), .ZN(_05410_ ) );
NAND3_X1 _12687_ ( .A1(_05138_ ), .A2(\EXU.pc_i [22] ), .A3(_05385_ ), .ZN(_05411_ ) );
XNOR2_X1 _12688_ ( .A(_05411_ ), .B(\EXU.pc_i [23] ), .ZN(_05412_ ) );
MUX2_X1 _12689_ ( .A(\EXU.mepc_i [23] ), .B(_05412_ ), .S(_05099_ ), .Z(_05413_ ) );
MUX2_X1 _12690_ ( .A(\EXU.mtvec_i [23] ), .B(_05413_ ), .S(_05050_ ), .Z(_05414_ ) );
OAI21_X1 _12691_ ( .A(_05082_ ), .B1(_05049_ ), .B2(_05414_ ), .ZN(_05415_ ) );
OAI22_X1 _12692_ ( .A1(_05410_ ), .A2(_05415_ ), .B1(_04253_ ), .B2(_05331_ ), .ZN(_00233_ ) );
XOR2_X1 _12693_ ( .A(_05405_ ), .B(_04553_ ), .Z(_05416_ ) );
NOR2_X1 _12694_ ( .A1(_05416_ ), .A2(_05042_ ), .ZN(_05417_ ) );
NAND4_X1 _12695_ ( .A1(_05092_ ), .A2(\EXU.op_i [4] ), .A3(\EXU.mtvec_i [22] ), .A4(_05055_ ), .ZN(_05418_ ) );
AND4_X1 _12696_ ( .A1(\EXU.op_i [4] ), .A2(_05053_ ), .A3(\EXU.mepc_i [22] ), .A4(_05119_ ), .ZN(_05419_ ) );
INV_X1 _12697_ ( .A(\EXU.pc_i [22] ), .ZN(_05420_ ) );
XNOR2_X1 _12698_ ( .A(_05386_ ), .B(_05420_ ), .ZN(_05421_ ) );
AOI21_X1 _12699_ ( .A(_05419_ ), .B1(_05421_ ), .B2(_05100_ ), .ZN(_05422_ ) );
OAI21_X1 _12700_ ( .A(_05418_ ), .B1(_05422_ ), .B2(_05103_ ), .ZN(_05423_ ) );
OAI21_X1 _12701_ ( .A(_05082_ ), .B1(_05049_ ), .B2(_05423_ ), .ZN(_05424_ ) );
OAI22_X1 _12702_ ( .A1(_05417_ ), .A2(_05424_ ), .B1(_04254_ ), .B2(_05331_ ), .ZN(_00234_ ) );
OAI211_X1 _12703_ ( .A(\EXU.state ), .B(\EXU.rd_i [3] ), .C1(_04393_ ), .C2(\LSU.ls_read_done_$_OR__B_Y_$_ORNOT__A_Y_$_ANDNOT__A_Y_$_OR__A_1_B ), .ZN(_05425_ ) );
NOR2_X1 _12704_ ( .A1(_04393_ ), .A2(\LSU.ls_read_done_$_OR__B_Y_$_ORNOT__A_Y_$_ANDNOT__A_Y_$_OR__A_1_B ), .ZN(_05426_ ) );
INV_X1 _12705_ ( .A(_05426_ ), .ZN(_05427_ ) );
INV_X1 _12706_ ( .A(\EXU.rd_o [3] ), .ZN(_05428_ ) );
OAI21_X1 _12707_ ( .A(_05425_ ), .B1(_05427_ ), .B2(_05428_ ), .ZN(_00236_ ) );
OAI211_X1 _12708_ ( .A(\EXU.state ), .B(\EXU.rd_i [2] ), .C1(_04393_ ), .C2(\LSU.ls_read_done_$_OR__B_Y_$_ORNOT__A_Y_$_ANDNOT__A_Y_$_OR__A_1_B ), .ZN(_05429_ ) );
INV_X1 _12709_ ( .A(\EXU.rd_o [2] ), .ZN(_05430_ ) );
OAI21_X1 _12710_ ( .A(_05429_ ), .B1(_05427_ ), .B2(_05430_ ), .ZN(_00237_ ) );
OAI211_X1 _12711_ ( .A(\EXU.state ), .B(\EXU.rd_i [1] ), .C1(_04393_ ), .C2(\LSU.ls_read_done_$_OR__B_Y_$_ORNOT__A_Y_$_ANDNOT__A_Y_$_OR__A_1_B ), .ZN(_05431_ ) );
INV_X1 _12712_ ( .A(\EXU.rd_o [1] ), .ZN(_05432_ ) );
OAI21_X1 _12713_ ( .A(_05431_ ), .B1(_05427_ ), .B2(_05432_ ), .ZN(_00238_ ) );
OAI211_X1 _12714_ ( .A(\EXU.state ), .B(\EXU.rd_i [0] ), .C1(_04393_ ), .C2(\LSU.ls_read_done_$_OR__B_Y_$_ORNOT__A_Y_$_ANDNOT__A_Y_$_OR__A_1_B ), .ZN(_05433_ ) );
INV_X1 _12715_ ( .A(\EXU.rd_o [0] ), .ZN(_05434_ ) );
OAI21_X1 _12716_ ( .A(_05433_ ), .B1(_05427_ ), .B2(_05434_ ), .ZN(_00239_ ) );
NOR2_X1 _12717_ ( .A1(\EXU.rd_o [3] ), .A2(\EXU.rd_o [2] ), .ZN(_05435_ ) );
AND3_X1 _12718_ ( .A1(_05435_ ), .A2(_05432_ ), .A3(_05434_ ), .ZN(_05436_ ) );
INV_X1 _12719_ ( .A(_03740_ ), .ZN(_05437_ ) );
OR4_X1 _12720_ ( .A1(\IDU.funct3 [2] ), .A2(_05437_ ), .A3(\IDU.funct3 [1] ), .A4(\IDU.funct3 [0] ), .ZN(_05438_ ) );
OR4_X1 _12721_ ( .A1(_03788_ ), .A2(_03785_ ), .A3(_03792_ ), .A4(_05438_ ), .ZN(_05439_ ) );
OR3_X2 _12722_ ( .A1(_05439_ ), .A2(_03835_ ), .A3(_03946_ ), .ZN(_05440_ ) );
INV_X1 _12723_ ( .A(_03819_ ), .ZN(_05441_ ) );
OAI211_X1 _12724_ ( .A(_03900_ ), .B(_03901_ ), .C1(\IDU.imm_$_NOR__Y_1_A_$_MUX__Y_B ), .C2(_03749_ ), .ZN(_05442_ ) );
AOI22_X1 _12725_ ( .A1(_03744_ ), .A2(_03747_ ), .B1(\IDU.imm_$_NOR__Y_2_A_$_MUX__Y_B ), .B2(\IDU.imm_$_NOR__Y_3_A_$_MUX__Y_B ), .ZN(_05443_ ) );
NOR4_X1 _12726_ ( .A1(_05440_ ), .A2(_05441_ ), .A3(_05442_ ), .A4(_05443_ ), .ZN(_05444_ ) );
NAND3_X1 _12727_ ( .A1(_03728_ ), .A2(\IDU.funct7 [6] ), .A3(_03745_ ), .ZN(_05445_ ) );
AND2_X1 _12728_ ( .A1(_03934_ ), .A2(_05445_ ), .ZN(_05446_ ) );
BUF_X4 _12729_ ( .A(_05446_ ), .Z(_05447_ ) );
BUF_X2 _12730_ ( .A(_03730_ ), .Z(_05448_ ) );
BUF_X2 _12731_ ( .A(_03735_ ), .Z(_05449_ ) );
NAND3_X1 _12732_ ( .A1(_05448_ ), .A2(\IDU.funct7 [0] ), .A3(_05449_ ), .ZN(_05450_ ) );
NAND2_X1 _12733_ ( .A1(_05447_ ), .A2(_05450_ ), .ZN(_05451_ ) );
NAND3_X1 _12734_ ( .A1(_05448_ ), .A2(\IDU.funct7 [1] ), .A3(_05449_ ), .ZN(_05452_ ) );
NAND2_X1 _12735_ ( .A1(_05447_ ), .A2(_05452_ ), .ZN(_05453_ ) );
NAND3_X1 _12736_ ( .A1(_03730_ ), .A2(\IDU.immI [4] ), .A3(_03735_ ), .ZN(_05454_ ) );
NAND2_X1 _12737_ ( .A1(_05447_ ), .A2(_05454_ ), .ZN(_05455_ ) );
NAND3_X1 _12738_ ( .A1(_03730_ ), .A2(\IDU.immI [3] ), .A3(_03735_ ), .ZN(_05456_ ) );
NAND2_X1 _12739_ ( .A1(_05446_ ), .A2(_05456_ ), .ZN(_05457_ ) );
OR4_X1 _12740_ ( .A1(_05451_ ), .A2(_05453_ ), .A3(_05455_ ), .A4(_05457_ ), .ZN(_05458_ ) );
NAND3_X1 _12741_ ( .A1(_05448_ ), .A2(\IDU.immI [1] ), .A3(_05449_ ), .ZN(_05459_ ) );
NAND2_X1 _12742_ ( .A1(_05447_ ), .A2(_05459_ ), .ZN(_05460_ ) );
NAND3_X1 _12743_ ( .A1(_05448_ ), .A2(\IDU.immI [0] ), .A3(_05449_ ), .ZN(_05461_ ) );
NAND2_X1 _12744_ ( .A1(_05447_ ), .A2(_05461_ ), .ZN(_05462_ ) );
INV_X1 _12745_ ( .A(_05447_ ), .ZN(_05463_ ) );
AND3_X1 _12746_ ( .A1(_05448_ ), .A2(\IDU.immI [2] ), .A3(_05449_ ), .ZN(_05464_ ) );
NOR2_X1 _12747_ ( .A1(_05463_ ), .A2(_05464_ ), .ZN(_05465_ ) );
INV_X1 _12748_ ( .A(_05465_ ), .ZN(_05466_ ) );
NOR4_X1 _12749_ ( .A1(_05458_ ), .A2(_05460_ ), .A3(_05462_ ), .A4(_05466_ ), .ZN(_05467_ ) );
AND3_X1 _12750_ ( .A1(_05448_ ), .A2(\IDU.funct7 [3] ), .A3(_05449_ ), .ZN(_05468_ ) );
NOR2_X1 _12751_ ( .A1(_05463_ ), .A2(_05468_ ), .ZN(_05469_ ) );
INV_X1 _12752_ ( .A(_05469_ ), .ZN(_05470_ ) );
NAND3_X1 _12753_ ( .A1(_05448_ ), .A2(\IDU.funct7 [4] ), .A3(_05449_ ), .ZN(_05471_ ) );
NAND2_X1 _12754_ ( .A1(_05447_ ), .A2(_05471_ ), .ZN(_05472_ ) );
NAND3_X1 _12755_ ( .A1(_05448_ ), .A2(\IDU.funct7 [5] ), .A3(_05449_ ), .ZN(_05473_ ) );
NAND2_X1 _12756_ ( .A1(_05447_ ), .A2(_05473_ ), .ZN(_05474_ ) );
NAND3_X1 _12757_ ( .A1(_05448_ ), .A2(\IDU.funct7 [2] ), .A3(_05449_ ), .ZN(_05475_ ) );
NAND2_X1 _12758_ ( .A1(_05447_ ), .A2(_05475_ ), .ZN(_05476_ ) );
NOR4_X1 _12759_ ( .A1(_05470_ ), .A2(_05472_ ), .A3(_05474_ ), .A4(_05476_ ), .ZN(_05477_ ) );
NAND3_X1 _12760_ ( .A1(_05448_ ), .A2(\IDU.funct7 [6] ), .A3(_05449_ ), .ZN(_05478_ ) );
NAND2_X1 _12761_ ( .A1(_05447_ ), .A2(_05478_ ), .ZN(_05479_ ) );
NOR4_X1 _12762_ ( .A1(_05479_ ), .A2(_03777_ ), .A3(_03772_ ), .A4(_03770_ ), .ZN(_05480_ ) );
NAND4_X1 _12763_ ( .A1(_05444_ ), .A2(_05467_ ), .A3(_05477_ ), .A4(_05480_ ), .ZN(_05481_ ) );
AND2_X1 _12764_ ( .A1(_03726_ ), .A2(_03743_ ), .ZN(_05482_ ) );
NAND2_X2 _12765_ ( .A1(_05481_ ), .A2(_05482_ ), .ZN(_05483_ ) );
OAI21_X1 _12766_ ( .A(\IDU.imm_$_NOR__Y_8_A_$_MUX__Y_B ), .B1(_03727_ ), .B2(_03742_ ), .ZN(_05484_ ) );
AND2_X1 _12767_ ( .A1(_05483_ ), .A2(_05484_ ), .ZN(_05485_ ) );
XNOR2_X1 _12768_ ( .A(_05485_ ), .B(\EXU.rd_o [3] ), .ZN(_05486_ ) );
OAI21_X1 _12769_ ( .A(\IDU.imm_$_NOR__Y_A_$_MUX__Y_B ), .B1(_03727_ ), .B2(_03742_ ), .ZN(_05487_ ) );
AND2_X1 _12770_ ( .A1(_05483_ ), .A2(_05487_ ), .ZN(_05488_ ) );
XNOR2_X1 _12771_ ( .A(_05488_ ), .B(\EXU.rd_o [0] ), .ZN(_05489_ ) );
OAI21_X1 _12772_ ( .A(\IDU.imm_$_NOR__Y_9_A_$_MUX__Y_B ), .B1(_03727_ ), .B2(_03742_ ), .ZN(_05490_ ) );
AND2_X1 _12773_ ( .A1(_05483_ ), .A2(_05490_ ), .ZN(_05491_ ) );
XNOR2_X1 _12774_ ( .A(_05491_ ), .B(\EXU.rd_o [2] ), .ZN(_05492_ ) );
OAI21_X1 _12775_ ( .A(\IDU.imm_$_NOR__Y_10_A_$_MUX__Y_B ), .B1(_03727_ ), .B2(_03742_ ), .ZN(_05493_ ) );
AND2_X1 _12776_ ( .A1(_05483_ ), .A2(_05493_ ), .ZN(_05494_ ) );
XNOR2_X1 _12777_ ( .A(_05494_ ), .B(\EXU.rd_o [1] ), .ZN(_05495_ ) );
NAND4_X1 _12778_ ( .A1(_05486_ ), .A2(_05489_ ), .A3(_05492_ ), .A4(_05495_ ), .ZN(_05496_ ) );
INV_X1 _12779_ ( .A(\IDU.immJ [18] ), .ZN(_05497_ ) );
NOR2_X1 _12780_ ( .A1(_03744_ ), .A2(_05497_ ), .ZN(_05498_ ) );
XNOR2_X1 _12781_ ( .A(_05498_ ), .B(\EXU.rd_o [3] ), .ZN(_05499_ ) );
NOR2_X1 _12782_ ( .A1(_03744_ ), .A2(_03949_ ), .ZN(_05500_ ) );
XNOR2_X1 _12783_ ( .A(_05500_ ), .B(\EXU.rd_o [0] ), .ZN(_05501_ ) );
INV_X1 _12784_ ( .A(\IDU.immJ [17] ), .ZN(_05502_ ) );
NOR2_X1 _12785_ ( .A1(_03744_ ), .A2(_05502_ ), .ZN(_05503_ ) );
XNOR2_X1 _12786_ ( .A(_05503_ ), .B(\EXU.rd_o [2] ), .ZN(_05504_ ) );
INV_X1 _12787_ ( .A(\IDU.immJ [16] ), .ZN(_05505_ ) );
NOR2_X1 _12788_ ( .A1(_03744_ ), .A2(_05505_ ), .ZN(_05506_ ) );
XNOR2_X1 _12789_ ( .A(_05506_ ), .B(\EXU.rd_o [1] ), .ZN(_05507_ ) );
NAND4_X1 _12790_ ( .A1(_05499_ ), .A2(_05501_ ), .A3(_05504_ ), .A4(_05507_ ), .ZN(_05508_ ) );
AOI21_X1 _12791_ ( .A(_05436_ ), .B1(_05496_ ), .B2(_05508_ ), .ZN(_05509_ ) );
INV_X1 _12792_ ( .A(\IDU.state ), .ZN(_05510_ ) );
NOR2_X1 _12793_ ( .A1(_05509_ ), .A2(_05510_ ), .ZN(_05511_ ) );
INV_X1 _12794_ ( .A(_05511_ ), .ZN(_05512_ ) );
NOR2_X1 _12795_ ( .A1(_05512_ ), .A2(\EXU.state ), .ZN(_05513_ ) );
BUF_X8 _12796_ ( .A(_05513_ ), .Z(_05514_ ) );
BUF_X2 _12797_ ( .A(_05514_ ), .Z(\IDU.updata ) );
BUF_X4 _12798_ ( .A(_04395_ ), .Z(_05515_ ) );
BUF_X4 _12799_ ( .A(_04355_ ), .Z(_05516_ ) );
AOI22_X1 _12800_ ( .A1(_05516_ ), .A2(\EXU.mstatus_i [31] ), .B1(_04336_ ), .B2(\EXU.mcause_i [31] ), .ZN(_05517_ ) );
BUF_X4 _12801_ ( .A(_04350_ ), .Z(_05518_ ) );
AOI22_X1 _12802_ ( .A1(_04353_ ), .A2(\EXU.mtvec_i [31] ), .B1(_05518_ ), .B2(\EXU.mepc_i [31] ), .ZN(_05519_ ) );
NAND2_X1 _12803_ ( .A1(_05517_ ), .A2(_05519_ ), .ZN(_05520_ ) );
INV_X1 _12804_ ( .A(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ), .ZN(_05521_ ) );
INV_X1 _12805_ ( .A(fanout_net_6 ), .ZN(_05522_ ) );
NOR2_X1 _12806_ ( .A1(_05522_ ), .A2(fanout_net_5 ), .ZN(_05523_ ) );
AND2_X1 _12807_ ( .A1(_05523_ ), .A2(fanout_net_10 ), .ZN(_05524_ ) );
BUF_X4 _12808_ ( .A(_05524_ ), .Z(_05525_ ) );
AND4_X1 _12809_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ), .A4(fanout_net_10 ), .ZN(_05526_ ) );
OAI22_X1 _12810_ ( .A1(_05520_ ), .A2(_05521_ ), .B1(_05525_ ), .B2(_05526_ ), .ZN(_05527_ ) );
BUF_X2 _12811_ ( .A(_04716_ ), .Z(_05528_ ) );
AOI22_X1 _12812_ ( .A1(_05103_ ), .A2(\EXU.pc_i [31] ), .B1(\EXU.r1_i [31] ), .B2(_05528_ ), .ZN(_05529_ ) );
NAND2_X1 _12813_ ( .A1(_05527_ ), .A2(_05529_ ), .ZN(_05530_ ) );
BUF_X4 _12814_ ( .A(_04417_ ), .Z(_05531_ ) );
NAND2_X1 _12815_ ( .A1(_04732_ ), .A2(_05531_ ), .ZN(_05532_ ) );
NOR2_X1 _12816_ ( .A1(_05532_ ), .A2(_04385_ ), .ZN(_05533_ ) );
NOR2_X1 _12817_ ( .A1(_04427_ ), .A2(_05533_ ), .ZN(_05534_ ) );
BUF_X4 _12818_ ( .A(_05534_ ), .Z(_05535_ ) );
NAND4_X1 _12819_ ( .A1(_04337_ ), .A2(_04338_ ), .A3(_04383_ ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_14_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05536_ ) );
NAND2_X4 _12820_ ( .A1(_04717_ ), .A2(_05536_ ), .ZN(_05537_ ) );
AND2_X1 _12821_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .ZN(_05538_ ) );
AND2_X1 _12822_ ( .A1(_05538_ ), .A2(_05026_ ), .ZN(_05539_ ) );
AND2_X1 _12823_ ( .A1(_05523_ ), .A2(_05026_ ), .ZN(_05540_ ) );
OAI21_X1 _12824_ ( .A(_05537_ ), .B1(_05539_ ), .B2(_05540_ ), .ZN(_05541_ ) );
INV_X1 _12825_ ( .A(_05541_ ), .ZN(_05542_ ) );
AND2_X2 _12826_ ( .A1(_04715_ ), .A2(_05026_ ), .ZN(_05543_ ) );
NAND4_X1 _12827_ ( .A1(_05543_ ), .A2(_04383_ ), .A3(_04340_ ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_14_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05544_ ) );
INV_X1 _12828_ ( .A(\EXU.funct7_i ), .ZN(_05545_ ) );
NAND4_X1 _12829_ ( .A1(_05543_ ), .A2(_05545_ ), .A3(_04387_ ), .A4(_04423_ ), .ZN(_05546_ ) );
AND2_X2 _12830_ ( .A1(_05544_ ), .A2(_05546_ ), .ZN(_05547_ ) );
INV_X2 _12831_ ( .A(_05547_ ), .ZN(_05548_ ) );
AND2_X4 _12832_ ( .A1(_05537_ ), .A2(_04716_ ), .ZN(_05549_ ) );
NOR3_X2 _12833_ ( .A1(_05542_ ), .A2(_05548_ ), .A3(_05549_ ), .ZN(_05550_ ) );
INV_X1 _12834_ ( .A(_05550_ ), .ZN(_05551_ ) );
AND3_X1 _12835_ ( .A1(_04434_ ), .A2(\EXU.funct7_i ), .A3(_04711_ ), .ZN(_05552_ ) );
INV_X1 _12836_ ( .A(_05552_ ), .ZN(_05553_ ) );
AND2_X4 _12837_ ( .A1(_05537_ ), .A2(_05540_ ), .ZN(_05554_ ) );
BUF_X8 _12838_ ( .A(_05554_ ), .Z(_05555_ ) );
INV_X4 _12839_ ( .A(_05555_ ), .ZN(_05556_ ) );
INV_X1 _12840_ ( .A(_05524_ ), .ZN(_05557_ ) );
INV_X1 _12841_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_14_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05558_ ) );
AND2_X1 _12842_ ( .A1(_05538_ ), .A2(fanout_net_10 ), .ZN(_05559_ ) );
INV_X1 _12843_ ( .A(_05559_ ), .ZN(_05560_ ) );
OAI22_X1 _12844_ ( .A1(_05557_ ), .A2(_05558_ ), .B1(_05560_ ), .B2(\EXU.funct7_i ), .ZN(_05561_ ) );
NAND2_X1 _12845_ ( .A1(_05561_ ), .A2(_04422_ ), .ZN(_05562_ ) );
OAI211_X1 _12846_ ( .A(_04387_ ), .B(_04423_ ), .C1(_05524_ ), .C2(_05559_ ), .ZN(_05563_ ) );
AND4_X4 _12847_ ( .A1(_05556_ ), .A2(_05547_ ), .A3(_05562_ ), .A4(_05563_ ), .ZN(_05564_ ) );
BUF_X4 _12848_ ( .A(_05549_ ), .Z(_05565_ ) );
OAI21_X4 _12849_ ( .A(_05553_ ), .B1(_05564_ ), .B2(_05565_ ), .ZN(_05566_ ) );
AND2_X1 _12850_ ( .A1(_05537_ ), .A2(_04711_ ), .ZN(_05567_ ) );
INV_X1 _12851_ ( .A(_05567_ ), .ZN(_05568_ ) );
AOI21_X4 _12852_ ( .A(_05551_ ), .B1(_05566_ ), .B2(_05568_ ), .ZN(_05569_ ) );
AND2_X1 _12853_ ( .A1(_04709_ ), .A2(_05026_ ), .ZN(_05570_ ) );
AND3_X1 _12854_ ( .A1(_05553_ ), .A2(_05570_ ), .A3(_05537_ ), .ZN(_05571_ ) );
BUF_X4 _12855_ ( .A(_05571_ ), .Z(_05572_ ) );
AND2_X1 _12856_ ( .A1(_05572_ ), .A2(_05568_ ), .ZN(_05573_ ) );
INV_X1 _12857_ ( .A(_05573_ ), .ZN(_05574_ ) );
INV_X1 _12858_ ( .A(_05565_ ), .ZN(_05575_ ) );
AND2_X1 _12859_ ( .A1(_05562_ ), .A2(_05563_ ), .ZN(_05576_ ) );
INV_X1 _12860_ ( .A(_05576_ ), .ZN(_05577_ ) );
NAND4_X1 _12861_ ( .A1(_05543_ ), .A2(_05558_ ), .A3(_04387_ ), .A4(_04423_ ), .ZN(_05578_ ) );
NAND4_X1 _12862_ ( .A1(_05543_ ), .A2(\EXU.funct7_i ), .A3(_04340_ ), .A4(_04383_ ), .ZN(_05579_ ) );
AND2_X1 _12863_ ( .A1(_05578_ ), .A2(_05579_ ), .ZN(_05580_ ) );
AOI21_X1 _12864_ ( .A(_05548_ ), .B1(_05541_ ), .B2(_05580_ ), .ZN(_05581_ ) );
OAI21_X1 _12865_ ( .A(_05575_ ), .B1(_05577_ ), .B2(_05581_ ), .ZN(_05582_ ) );
AND2_X1 _12866_ ( .A1(_05574_ ), .A2(_05582_ ), .ZN(_05583_ ) );
AND2_X1 _12867_ ( .A1(_05569_ ), .A2(_05583_ ), .ZN(_05584_ ) );
BUF_X4 _12868_ ( .A(_05584_ ), .Z(_05585_ ) );
NAND2_X1 _12869_ ( .A1(_04653_ ), .A2(_05585_ ), .ZN(_05586_ ) );
AND3_X4 _12870_ ( .A1(_04392_ ), .A2(_04370_ ), .A3(_04424_ ), .ZN(_05587_ ) );
INV_X2 _12871_ ( .A(_05587_ ), .ZN(_05588_ ) );
INV_X4 _12872_ ( .A(_05569_ ), .ZN(_05589_ ) );
NOR2_X2 _12873_ ( .A1(_05589_ ), .A2(_05582_ ), .ZN(_05590_ ) );
INV_X4 _12874_ ( .A(_05590_ ), .ZN(_05591_ ) );
NOR4_X4 _12875_ ( .A1(_05588_ ), .A2(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B ), .A3(_04395_ ), .A4(_05591_ ), .ZN(_05592_ ) );
AND2_X4 _12876_ ( .A1(_05590_ ), .A2(_04332_ ), .ZN(_05593_ ) );
AND3_X1 _12877_ ( .A1(_04392_ ), .A2(_04370_ ), .A3(_04436_ ), .ZN(_05594_ ) );
OAI21_X2 _12878_ ( .A(_05593_ ), .B1(_05587_ ), .B2(_05594_ ), .ZN(_05595_ ) );
AOI21_X2 _12879_ ( .A(\LSU.ls_wdata_i_$_MUX__Y_23_A_$_ANDNOT__Y_B ), .B1(_05593_ ), .B2(_05587_ ), .ZN(_05596_ ) );
NOR3_X4 _12880_ ( .A1(_05592_ ), .A2(_05595_ ), .A3(_05596_ ), .ZN(_05597_ ) );
AND2_X2 _12881_ ( .A1(_05595_ ), .A2(_04909_ ), .ZN(_05598_ ) );
NOR2_X4 _12882_ ( .A1(_05597_ ), .A2(_05598_ ), .ZN(_05599_ ) );
BUF_X8 _12883_ ( .A(_05599_ ), .Z(_05600_ ) );
BUF_X8 _12884_ ( .A(_05600_ ), .Z(_05601_ ) );
BUF_X4 _12885_ ( .A(_04902_ ), .Z(_05602_ ) );
BUF_X4 _12886_ ( .A(_05602_ ), .Z(_05603_ ) );
BUF_X4 _12887_ ( .A(_05603_ ), .Z(_05604_ ) );
NOR3_X1 _12888_ ( .A1(_05601_ ), .A2(_04725_ ), .A3(_05604_ ), .ZN(_05605_ ) );
BUF_X4 _12889_ ( .A(_04892_ ), .Z(_05606_ ) );
BUF_X4 _12890_ ( .A(_05606_ ), .Z(_05607_ ) );
AND3_X1 _12891_ ( .A1(_05605_ ), .A2(_04885_ ), .A3(_05607_ ), .ZN(_05608_ ) );
NAND3_X1 _12892_ ( .A1(_05593_ ), .A2(\EXU.imm_i [0] ), .A3(_05587_ ), .ZN(_05609_ ) );
AND2_X4 _12893_ ( .A1(_05593_ ), .A2(_05587_ ), .ZN(_05610_ ) );
BUF_X4 _12894_ ( .A(_04904_ ), .Z(_05611_ ) );
OAI21_X1 _12895_ ( .A(_05609_ ), .B1(_05610_ ), .B2(_05611_ ), .ZN(_05612_ ) );
INV_X1 _12896_ ( .A(_05612_ ), .ZN(_05613_ ) );
AND3_X1 _12897_ ( .A1(_05593_ ), .A2(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_05587_ ), .ZN(_05614_ ) );
AOI21_X1 _12898_ ( .A(_04896_ ), .B1(_05593_ ), .B2(_05587_ ), .ZN(_05615_ ) );
OR2_X2 _12899_ ( .A1(_05614_ ), .A2(_05615_ ), .ZN(_05616_ ) );
NAND3_X1 _12900_ ( .A1(_05593_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .A3(_05587_ ), .ZN(_05617_ ) );
OAI21_X4 _12901_ ( .A(_05617_ ), .B1(_05610_ ), .B2(_04888_ ), .ZN(_05618_ ) );
AND3_X2 _12902_ ( .A1(_05613_ ), .A2(_05616_ ), .A3(_05618_ ), .ZN(_05619_ ) );
NAND3_X1 _12903_ ( .A1(_05593_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_21_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_05587_ ), .ZN(_05620_ ) );
OAI21_X1 _12904_ ( .A(_05620_ ), .B1(_05610_ ), .B2(_04880_ ), .ZN(_05621_ ) );
NAND2_X4 _12905_ ( .A1(_05619_ ), .A2(_05621_ ), .ZN(_05622_ ) );
AND3_X1 _12906_ ( .A1(_05593_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_20_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_05587_ ), .ZN(_05623_ ) );
INV_X1 _12907_ ( .A(_05610_ ), .ZN(_05624_ ) );
AOI21_X1 _12908_ ( .A(_05623_ ), .B1(_05624_ ), .B2(\LSU.ls_wdata_i_$_MUX__Y_19_A_$_ANDNOT__Y_B ), .ZN(_05625_ ) );
NOR2_X4 _12909_ ( .A1(_05622_ ), .A2(_05625_ ), .ZN(_05626_ ) );
INV_X1 _12910_ ( .A(_05626_ ), .ZN(_05627_ ) );
AOI22_X1 _12911_ ( .A1(_05608_ ), .A2(_04954_ ), .B1(_05627_ ), .B2(\EXU.r1_i [31] ), .ZN(_05628_ ) );
NOR2_X1 _12912_ ( .A1(_05628_ ), .A2(_05591_ ), .ZN(_05629_ ) );
BUF_X4 _12913_ ( .A(_05568_ ), .Z(_05630_ ) );
NAND3_X1 _12914_ ( .A1(_04720_ ), .A2(\EXU.r1_i [31] ), .A3(_04723_ ), .ZN(_05631_ ) );
NAND3_X1 _12915_ ( .A1(_05572_ ), .A2(_05630_ ), .A3(_05631_ ), .ZN(_05632_ ) );
AOI21_X1 _12916_ ( .A(_04726_ ), .B1(_05632_ ), .B2(_05556_ ), .ZN(_05633_ ) );
AND2_X1 _12917_ ( .A1(_05537_ ), .A2(_05539_ ), .ZN(_05634_ ) );
INV_X2 _12918_ ( .A(_05634_ ), .ZN(_05635_ ) );
MUX2_X1 _12919_ ( .A(_04727_ ), .B(_05633_ ), .S(_05635_ ), .Z(_05636_ ) );
OR2_X1 _12920_ ( .A1(_05629_ ), .A2(_05636_ ), .ZN(_05637_ ) );
AND3_X1 _12921_ ( .A1(_05566_ ), .A2(_05550_ ), .A3(_05630_ ), .ZN(_05638_ ) );
AND2_X1 _12922_ ( .A1(_05638_ ), .A2(_05583_ ), .ZN(_05639_ ) );
INV_X1 _12923_ ( .A(_05639_ ), .ZN(_05640_ ) );
BUF_X4 _12924_ ( .A(_05640_ ), .Z(_05641_ ) );
INV_X1 _12925_ ( .A(_04661_ ), .ZN(_05642_ ) );
INV_X1 _12926_ ( .A(_04662_ ), .ZN(_05643_ ) );
OAI21_X1 _12927_ ( .A(_04654_ ), .B1(\EXU.r1_i [0] ), .B2(_04904_ ), .ZN(_05644_ ) );
OR2_X1 _12928_ ( .A1(_05000_ ), .A2(\EXU.r2_i [1] ), .ZN(_05645_ ) );
AOI211_X1 _12929_ ( .A(_05642_ ), .B(_05643_ ), .C1(_05644_ ), .C2(_05645_ ), .ZN(_05646_ ) );
NOR2_X1 _12930_ ( .A1(_04893_ ), .A2(\EXU.r2_i [2] ), .ZN(_05647_ ) );
NAND2_X1 _12931_ ( .A1(_04661_ ), .A2(_05647_ ), .ZN(_05648_ ) );
INV_X1 _12932_ ( .A(\EXU.r1_i [3] ), .ZN(_05649_ ) );
OAI21_X1 _12933_ ( .A(_05648_ ), .B1(_05649_ ), .B2(\EXU.r2_i [3] ), .ZN(_05650_ ) );
NOR2_X1 _12934_ ( .A1(_05646_ ), .A2(_05650_ ), .ZN(_05651_ ) );
INV_X1 _12935_ ( .A(_05651_ ), .ZN(_05652_ ) );
AND3_X1 _12936_ ( .A1(_05652_ ), .A2(_04669_ ), .A3(_04672_ ), .ZN(_05653_ ) );
NOR2_X1 _12937_ ( .A1(_04955_ ), .A2(\EXU.r2_i [4] ), .ZN(_05654_ ) );
NAND2_X1 _12938_ ( .A1(_04670_ ), .A2(_05654_ ), .ZN(_05655_ ) );
OAI21_X1 _12939_ ( .A(_05655_ ), .B1(_05006_ ), .B2(\EXU.r2_i [5] ), .ZN(_05656_ ) );
NAND2_X1 _12940_ ( .A1(_05656_ ), .A2(_04669_ ), .ZN(_05657_ ) );
INV_X1 _12941_ ( .A(_04667_ ), .ZN(_05658_ ) );
OR2_X1 _12942_ ( .A1(_04940_ ), .A2(\EXU.r2_i [6] ), .ZN(_05659_ ) );
OR2_X1 _12943_ ( .A1(_05658_ ), .A2(_05659_ ), .ZN(_05660_ ) );
OAI211_X1 _12944_ ( .A(_05657_ ), .B(_05660_ ), .C1(_04930_ ), .C2(\EXU.r2_i [7] ), .ZN(_05661_ ) );
OAI211_X1 _12945_ ( .A(_04687_ ), .B(_04700_ ), .C1(_05653_ ), .C2(_05661_ ), .ZN(_05662_ ) );
INV_X1 _12946_ ( .A(\EXU.r2_i [14] ), .ZN(_05663_ ) );
NAND3_X1 _12947_ ( .A1(_04680_ ), .A2(\EXU.r1_i [14] ), .A3(_05663_ ), .ZN(_05664_ ) );
NOR2_X1 _12948_ ( .A1(_04877_ ), .A2(\EXU.r2_i [12] ), .ZN(_05665_ ) );
AND2_X1 _12949_ ( .A1(_04683_ ), .A2(_05665_ ), .ZN(_05666_ ) );
INV_X1 _12950_ ( .A(\EXU.r2_i [13] ), .ZN(_05667_ ) );
AOI21_X1 _12951_ ( .A(_05666_ ), .B1(\EXU.r1_i [13] ), .B2(_05667_ ), .ZN(_05668_ ) );
OAI221_X1 _12952_ ( .A(_05664_ ), .B1(_05017_ ), .B2(\EXU.r2_i [15] ), .C1(_05668_ ), .C2(_04682_ ), .ZN(_05669_ ) );
NOR2_X1 _12953_ ( .A1(_04926_ ), .A2(\EXU.r2_i [8] ), .ZN(_05670_ ) );
AND2_X1 _12954_ ( .A1(_04697_ ), .A2(_05670_ ), .ZN(_05671_ ) );
INV_X1 _12955_ ( .A(\EXU.r2_i [9] ), .ZN(_05672_ ) );
AOI21_X1 _12956_ ( .A(_05671_ ), .B1(\EXU.r1_i [9] ), .B2(_05672_ ), .ZN(_05673_ ) );
INV_X1 _12957_ ( .A(_04696_ ), .ZN(_05674_ ) );
NOR2_X1 _12958_ ( .A1(_05673_ ), .A2(_05674_ ), .ZN(_05675_ ) );
NOR2_X1 _12959_ ( .A1(_04841_ ), .A2(\EXU.r2_i [11] ), .ZN(_05676_ ) );
NOR2_X1 _12960_ ( .A1(_04849_ ), .A2(\EXU.r2_i [10] ), .ZN(_05677_ ) );
AND2_X1 _12961_ ( .A1(_04694_ ), .A2(_05677_ ), .ZN(_05678_ ) );
NOR3_X1 _12962_ ( .A1(_05675_ ), .A2(_05676_ ), .A3(_05678_ ), .ZN(_05679_ ) );
INV_X1 _12963_ ( .A(_05679_ ), .ZN(_05680_ ) );
AOI21_X1 _12964_ ( .A(_05669_ ), .B1(_05680_ ), .B2(_04687_ ), .ZN(_05681_ ) );
NAND2_X1 _12965_ ( .A1(_05662_ ), .A2(_05681_ ), .ZN(_05682_ ) );
NAND3_X1 _12966_ ( .A1(_05682_ ), .A2(_04693_ ), .A3(_04707_ ), .ZN(_05683_ ) );
INV_X1 _12967_ ( .A(\EXU.r2_i [22] ), .ZN(_05684_ ) );
NAND3_X1 _12968_ ( .A1(_04691_ ), .A2(\EXU.r1_i [22] ), .A3(_05684_ ), .ZN(_05685_ ) );
NOR2_X1 _12969_ ( .A1(_04835_ ), .A2(\EXU.r2_i [20] ), .ZN(_05686_ ) );
AND2_X1 _12970_ ( .A1(_04688_ ), .A2(_05686_ ), .ZN(_05687_ ) );
INV_X1 _12971_ ( .A(\EXU.r2_i [21] ), .ZN(_05688_ ) );
AOI21_X1 _12972_ ( .A(_05687_ ), .B1(\EXU.r1_i [21] ), .B2(_05688_ ), .ZN(_05689_ ) );
NAND2_X1 _12973_ ( .A1(_04691_ ), .A2(_04692_ ), .ZN(_05690_ ) );
OAI221_X1 _12974_ ( .A(_05685_ ), .B1(_04792_ ), .B2(\EXU.r2_i [23] ), .C1(_05689_ ), .C2(_05690_ ), .ZN(_05691_ ) );
NOR2_X1 _12975_ ( .A1(_04764_ ), .A2(\EXU.r2_i [16] ), .ZN(_05692_ ) );
AND2_X1 _12976_ ( .A1(_04704_ ), .A2(_05692_ ), .ZN(_05693_ ) );
INV_X1 _12977_ ( .A(\EXU.r2_i [17] ), .ZN(_05694_ ) );
AOI21_X1 _12978_ ( .A(_05693_ ), .B1(\EXU.r1_i [17] ), .B2(_05694_ ), .ZN(_05695_ ) );
INV_X1 _12979_ ( .A(_04703_ ), .ZN(_05696_ ) );
OR2_X1 _12980_ ( .A1(_05695_ ), .A2(_05696_ ), .ZN(_05697_ ) );
NOR2_X1 _12981_ ( .A1(_04742_ ), .A2(\EXU.r2_i [18] ), .ZN(_05698_ ) );
AND2_X1 _12982_ ( .A1(_04701_ ), .A2(_05698_ ), .ZN(_05699_ ) );
INV_X1 _12983_ ( .A(\EXU.r2_i [19] ), .ZN(_05700_ ) );
AOI21_X1 _12984_ ( .A(_05699_ ), .B1(\EXU.r1_i [19] ), .B2(_05700_ ), .ZN(_05701_ ) );
AND2_X1 _12985_ ( .A1(_05697_ ), .A2(_05701_ ), .ZN(_05702_ ) );
INV_X1 _12986_ ( .A(_05702_ ), .ZN(_05703_ ) );
AOI21_X1 _12987_ ( .A(_05691_ ), .B1(_05703_ ), .B2(_04693_ ), .ZN(_05704_ ) );
AND2_X1 _12988_ ( .A1(_05683_ ), .A2(_05704_ ), .ZN(_05705_ ) );
INV_X1 _12989_ ( .A(_05705_ ), .ZN(_05706_ ) );
AND2_X1 _12990_ ( .A1(_05706_ ), .A2(_04678_ ), .ZN(_05707_ ) );
NOR2_X1 _12991_ ( .A1(_04814_ ), .A2(\EXU.r2_i [25] ), .ZN(_05708_ ) );
NOR2_X1 _12992_ ( .A1(_04821_ ), .A2(\EXU.r2_i [24] ), .ZN(_05709_ ) );
AOI21_X1 _12993_ ( .A(_05708_ ), .B1(_04673_ ), .B2(_05709_ ), .ZN(_05710_ ) );
INV_X1 _12994_ ( .A(_05710_ ), .ZN(_05711_ ) );
AND3_X1 _12995_ ( .A1(_05711_ ), .A2(_04676_ ), .A3(_04677_ ), .ZN(_05712_ ) );
NOR2_X1 _12996_ ( .A1(_04801_ ), .A2(\EXU.r2_i [27] ), .ZN(_05713_ ) );
INV_X1 _12997_ ( .A(\EXU.r2_i [26] ), .ZN(_05714_ ) );
AND3_X1 _12998_ ( .A1(_04676_ ), .A2(\EXU.r1_i [26] ), .A3(_05714_ ), .ZN(_05715_ ) );
OR3_X1 _12999_ ( .A1(_05712_ ), .A2(_05713_ ), .A3(_05715_ ), .ZN(_05716_ ) );
OAI211_X1 _13000_ ( .A(_04663_ ), .B(_04664_ ), .C1(_05707_ ), .C2(_05716_ ), .ZN(_05717_ ) );
NOR2_X1 _13001_ ( .A1(_04771_ ), .A2(\EXU.r2_i [29] ), .ZN(_05718_ ) );
NOR2_X1 _13002_ ( .A1(_04778_ ), .A2(\EXU.r2_i [28] ), .ZN(_05719_ ) );
AOI21_X1 _13003_ ( .A(_05718_ ), .B1(_04663_ ), .B2(_05719_ ), .ZN(_05720_ ) );
AOI21_X1 _13004_ ( .A(_04657_ ), .B1(_05717_ ), .B2(_05720_ ), .ZN(_05721_ ) );
NOR2_X1 _13005_ ( .A1(_04736_ ), .A2(\EXU.r2_i [30] ), .ZN(_05722_ ) );
OR3_X1 _13006_ ( .A1(_05721_ ), .A2(_04659_ ), .A3(_05722_ ), .ZN(_05723_ ) );
OAI21_X1 _13007_ ( .A(_04659_ ), .B1(_05721_ ), .B2(_05722_ ), .ZN(_05724_ ) );
AOI21_X1 _13008_ ( .A(_05641_ ), .B1(_05723_ ), .B2(_05724_ ), .ZN(_05725_ ) );
BUF_X4 _13009_ ( .A(_04908_ ), .Z(_05726_ ) );
NAND2_X1 _13010_ ( .A1(_05726_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05727_ ) );
BUF_X2 _13011_ ( .A(_04907_ ), .Z(_05728_ ) );
OAI211_X1 _13012_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_22_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(_05728_ ), .C1(_04984_ ), .C2(_05611_ ), .ZN(_05729_ ) );
NAND2_X1 _13013_ ( .A1(_05727_ ), .A2(_05729_ ), .ZN(_05730_ ) );
NAND2_X1 _13014_ ( .A1(_05730_ ), .A2(_05603_ ), .ZN(_05731_ ) );
NAND2_X1 _13015_ ( .A1(_05726_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_21_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05732_ ) );
OAI211_X1 _13016_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_20_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(_04907_ ), .C1(_04984_ ), .C2(_05611_ ), .ZN(_05733_ ) );
NAND2_X1 _13017_ ( .A1(_05732_ ), .A2(_05733_ ), .ZN(_05734_ ) );
BUF_X4 _13018_ ( .A(_04901_ ), .Z(_05735_ ) );
NAND2_X1 _13019_ ( .A1(_05734_ ), .A2(_05735_ ), .ZN(_05736_ ) );
NAND2_X1 _13020_ ( .A1(_05731_ ), .A2(_05736_ ), .ZN(_05737_ ) );
NOR2_X1 _13021_ ( .A1(_04908_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05738_ ) );
AOI21_X1 _13022_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_19_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_04906_ ), .B2(_04907_ ), .ZN(_05739_ ) );
OR3_X1 _13023_ ( .A1(_05738_ ), .A2(_04901_ ), .A3(_05739_ ), .ZN(_05740_ ) );
AND3_X1 _13024_ ( .A1(_04906_ ), .A2(_04854_ ), .A3(_04907_ ), .ZN(_05741_ ) );
AOI21_X1 _13025_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B1(_04906_ ), .B2(_04907_ ), .ZN(_05742_ ) );
NOR2_X1 _13026_ ( .A1(_05741_ ), .A2(_05742_ ), .ZN(_05743_ ) );
NAND2_X1 _13027_ ( .A1(_05743_ ), .A2(_05735_ ), .ZN(_05744_ ) );
NAND2_X1 _13028_ ( .A1(_05740_ ), .A2(_05744_ ), .ZN(_05745_ ) );
MUX2_X1 _13029_ ( .A(_05737_ ), .B(_05745_ ), .S(_05606_ ), .Z(_05746_ ) );
BUF_X4 _13030_ ( .A(_04885_ ), .Z(_05747_ ) );
NAND2_X1 _13031_ ( .A1(_05746_ ), .A2(_05747_ ), .ZN(_05748_ ) );
NAND2_X1 _13032_ ( .A1(_05726_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05749_ ) );
BUF_X4 _13033_ ( .A(_04908_ ), .Z(_05750_ ) );
OAI211_X1 _13034_ ( .A(_05749_ ), .B(_04901_ ), .C1(_04929_ ), .C2(_05750_ ), .ZN(_05751_ ) );
NAND2_X1 _13035_ ( .A1(_04908_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_27_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05752_ ) );
OAI211_X1 _13036_ ( .A(_05752_ ), .B(_05602_ ), .C1(_04944_ ), .C2(_05726_ ), .ZN(_05753_ ) );
AND2_X1 _13037_ ( .A1(_05751_ ), .A2(_05753_ ), .ZN(_05754_ ) );
BUF_X4 _13038_ ( .A(_04996_ ), .Z(_05755_ ) );
OR2_X1 _13039_ ( .A1(_05754_ ), .A2(_05755_ ), .ZN(_05756_ ) );
BUF_X2 _13040_ ( .A(_04886_ ), .Z(_05757_ ) );
NAND2_X1 _13041_ ( .A1(_05750_ ), .A2(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_B_$_MUX__Y_A ), .ZN(_05758_ ) );
BUF_X4 _13042_ ( .A(_04984_ ), .Z(_05759_ ) );
BUF_X4 _13043_ ( .A(_05611_ ), .Z(_05760_ ) );
OAI211_X1 _13044_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(_05728_ ), .C1(_05759_ ), .C2(_05760_ ), .ZN(_05761_ ) );
NAND2_X1 _13045_ ( .A1(_05758_ ), .A2(_05761_ ), .ZN(_05762_ ) );
MUX2_X1 _13046_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_A ), .S(_04908_ ), .Z(_05763_ ) );
MUX2_X1 _13047_ ( .A(_05762_ ), .B(_05763_ ), .S(_05603_ ), .Z(_05764_ ) );
OAI211_X1 _13048_ ( .A(_05756_ ), .B(_05757_ ), .C1(_05607_ ), .C2(_05764_ ), .ZN(_05765_ ) );
AOI21_X1 _13049_ ( .A(_04954_ ), .B1(_05748_ ), .B2(_05765_ ), .ZN(_05766_ ) );
BUF_X2 _13050_ ( .A(_05575_ ), .Z(_05767_ ) );
OR2_X1 _13051_ ( .A1(_05766_ ), .A2(_05767_ ), .ZN(_05768_ ) );
BUF_X4 _13052_ ( .A(_04954_ ), .Z(_05769_ ) );
INV_X1 _13053_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_11_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05770_ ) );
NAND2_X1 _13054_ ( .A1(_05726_ ), .A2(_05770_ ), .ZN(_05771_ ) );
OAI211_X1 _13055_ ( .A(_04825_ ), .B(_05728_ ), .C1(_04984_ ), .C2(_05611_ ), .ZN(_05772_ ) );
NAND2_X1 _13056_ ( .A1(_05771_ ), .A2(_05772_ ), .ZN(_05773_ ) );
BUF_X2 _13057_ ( .A(_05602_ ), .Z(_05774_ ) );
NAND2_X1 _13058_ ( .A1(_05773_ ), .A2(_05774_ ), .ZN(_05775_ ) );
AND3_X1 _13059_ ( .A1(_04906_ ), .A2(_04794_ ), .A3(_04907_ ), .ZN(_05776_ ) );
AOI21_X1 _13060_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ), .B1(_04906_ ), .B2(_05728_ ), .ZN(_05777_ ) );
OAI21_X1 _13061_ ( .A(_05735_ ), .B1(_05776_ ), .B2(_05777_ ), .ZN(_05778_ ) );
AOI21_X1 _13062_ ( .A(_05755_ ), .B1(_05775_ ), .B2(_05778_ ), .ZN(_05779_ ) );
NAND2_X1 _13063_ ( .A1(_05750_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05780_ ) );
BUF_X4 _13064_ ( .A(_05726_ ), .Z(_05781_ ) );
OAI211_X1 _13065_ ( .A(_05780_ ), .B(_05774_ ), .C1(_04755_ ), .C2(_05781_ ), .ZN(_05782_ ) );
NAND2_X1 _13066_ ( .A1(_05750_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_13_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05783_ ) );
BUF_X4 _13067_ ( .A(_04901_ ), .Z(_05784_ ) );
BUF_X4 _13068_ ( .A(_04907_ ), .Z(_05785_ ) );
OAI211_X1 _13069_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_12_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(_05785_ ), .C1(_05759_ ), .C2(_05760_ ), .ZN(_05786_ ) );
NAND3_X1 _13070_ ( .A1(_05783_ ), .A2(_05784_ ), .A3(_05786_ ), .ZN(_05787_ ) );
AOI21_X1 _13071_ ( .A(_05606_ ), .B1(_05782_ ), .B2(_05787_ ), .ZN(_05788_ ) );
NOR2_X1 _13072_ ( .A1(_05779_ ), .A2(_05788_ ), .ZN(_05789_ ) );
NAND2_X1 _13073_ ( .A1(_05781_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_5_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05790_ ) );
OAI211_X1 _13074_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_4_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(_05785_ ), .C1(_05759_ ), .C2(_05760_ ), .ZN(_05791_ ) );
NAND3_X1 _13075_ ( .A1(_05790_ ), .A2(_05784_ ), .A3(_05791_ ), .ZN(_05792_ ) );
NAND2_X1 _13076_ ( .A1(_05750_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ), .ZN(_05793_ ) );
OAI211_X1 _13077_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_6_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(_05728_ ), .C1(_04984_ ), .C2(_05611_ ), .ZN(_05794_ ) );
NAND3_X1 _13078_ ( .A1(_05793_ ), .A2(_05774_ ), .A3(_05794_ ), .ZN(_05795_ ) );
AND2_X1 _13079_ ( .A1(_05792_ ), .A2(_05795_ ), .ZN(_05796_ ) );
NAND2_X1 _13080_ ( .A1(_05781_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_3_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05797_ ) );
OAI211_X1 _13081_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_2_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(_05785_ ), .C1(_05759_ ), .C2(_05760_ ), .ZN(_05798_ ) );
NAND2_X1 _13082_ ( .A1(_05797_ ), .A2(_05798_ ), .ZN(_05799_ ) );
MUX2_X1 _13083_ ( .A(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_A ), .S(_05726_ ), .Z(_05800_ ) );
MUX2_X1 _13084_ ( .A(_05799_ ), .B(_05800_ ), .S(_05784_ ), .Z(_05801_ ) );
BUF_X4 _13085_ ( .A(_04892_ ), .Z(_05802_ ) );
MUX2_X1 _13086_ ( .A(_05796_ ), .B(_05801_ ), .S(_05802_ ), .Z(_05803_ ) );
BUF_X4 _13087_ ( .A(_04885_ ), .Z(_05804_ ) );
MUX2_X1 _13088_ ( .A(_05789_ ), .B(_05803_ ), .S(_05804_ ), .Z(_05805_ ) );
AOI21_X1 _13089_ ( .A(_05768_ ), .B1(_05769_ ), .B2(_05805_ ), .ZN(_05806_ ) );
BUF_X2 _13090_ ( .A(_04954_ ), .Z(_05807_ ) );
AND3_X1 _13091_ ( .A1(_05566_ ), .A2(_05551_ ), .A3(_05568_ ), .ZN(_05808_ ) );
AND2_X1 _13092_ ( .A1(_05808_ ), .A2(_05583_ ), .ZN(_05809_ ) );
AND4_X1 _13093_ ( .A1(_04427_ ), .A2(_05608_ ), .A3(_05807_ ), .A4(_05809_ ), .ZN(_05810_ ) );
NOR4_X1 _13094_ ( .A1(_05637_ ), .A2(_05725_ ), .A3(_05806_ ), .A4(_05810_ ), .ZN(_05811_ ) );
AOI21_X1 _13095_ ( .A(_05535_ ), .B1(_05586_ ), .B2(_05811_ ), .ZN(_05812_ ) );
NOR2_X1 _13096_ ( .A1(_05075_ ), .A2(_05037_ ), .ZN(_05813_ ) );
INV_X1 _13097_ ( .A(_04343_ ), .ZN(_05814_ ) );
AOI21_X1 _13098_ ( .A(_05814_ ), .B1(_05517_ ), .B2(_05519_ ), .ZN(_05815_ ) );
NAND3_X1 _13099_ ( .A1(_04387_ ), .A2(\EXU.ls_rdata_i [31] ), .A3(_04388_ ), .ZN(_05816_ ) );
AND3_X2 _13100_ ( .A1(\EXU.op_i [3] ), .A2(\EXU.op_i [2] ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B ), .ZN(_05817_ ) );
NAND3_X1 _13101_ ( .A1(_05817_ ), .A2(_05531_ ), .A3(\EXU.imm_i [31] ), .ZN(_05818_ ) );
NAND2_X1 _13102_ ( .A1(_05816_ ), .A2(_05818_ ), .ZN(_05819_ ) );
OR4_X2 _13103_ ( .A1(_05812_ ), .A2(_05813_ ), .A3(_05815_ ), .A4(_05819_ ), .ZN(_05820_ ) );
INV_X1 _13104_ ( .A(_04394_ ), .ZN(_05821_ ) );
BUF_X4 _13105_ ( .A(_05821_ ), .Z(_05822_ ) );
MUX2_X2 _13106_ ( .A(_05530_ ), .B(_05820_ ), .S(_05822_ ), .Z(_05823_ ) );
INV_X1 _13107_ ( .A(_04376_ ), .ZN(_05824_ ) );
BUF_X4 _13108_ ( .A(_05824_ ), .Z(_05825_ ) );
NAND2_X1 _13109_ ( .A1(_05823_ ), .A2(_05825_ ), .ZN(_05826_ ) );
NAND3_X1 _13110_ ( .A1(_04377_ ), .A2(_05051_ ), .A3(_05530_ ), .ZN(_05827_ ) );
AOI21_X1 _13111_ ( .A(_05515_ ), .B1(_05826_ ), .B2(_05827_ ), .ZN(_05828_ ) );
MUX2_X1 _13112_ ( .A(\EXU.xrd_o [31] ), .B(_05828_ ), .S(_04400_ ), .Z(_00241_ ) );
INV_X2 _13113_ ( .A(_04355_ ), .ZN(_05829_ ) );
BUF_X4 _13114_ ( .A(_05829_ ), .Z(_05830_ ) );
BUF_X2 _13115_ ( .A(_04349_ ), .Z(_05831_ ) );
BUF_X4 _13116_ ( .A(_05052_ ), .Z(_05832_ ) );
NAND4_X1 _13117_ ( .A1(_05831_ ), .A2(_05832_ ), .A3(\EXU.mtvec_i [30] ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05833_ ) );
NOR2_X1 _13118_ ( .A1(_04344_ ), .A2(\EXU.imm_i [0] ), .ZN(_05834_ ) );
INV_X1 _13119_ ( .A(_05834_ ), .ZN(_05835_ ) );
BUF_X2 _13120_ ( .A(_04335_ ), .Z(_05836_ ) );
BUF_X2 _13121_ ( .A(_04334_ ), .Z(_05837_ ) );
AOI22_X1 _13122_ ( .A1(_05833_ ), .A2(_05835_ ), .B1(_05836_ ), .B2(_05837_ ), .ZN(_05838_ ) );
CLKBUF_X2 _13123_ ( .A(_04335_ ), .Z(_05839_ ) );
AND3_X1 _13124_ ( .A1(_05837_ ), .A2(\EXU.mcause_i [30] ), .A3(_05839_ ), .ZN(_05840_ ) );
OAI21_X1 _13125_ ( .A(_05830_ ), .B1(_05838_ ), .B2(_05840_ ), .ZN(_05841_ ) );
AOI22_X1 _13126_ ( .A1(_05516_ ), .A2(\EXU.mstatus_i [30] ), .B1(_05518_ ), .B2(\EXU.mepc_i [30] ), .ZN(_05842_ ) );
NAND2_X1 _13127_ ( .A1(_05841_ ), .A2(_05842_ ), .ZN(_05843_ ) );
INV_X1 _13128_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_A ), .ZN(_05844_ ) );
AND4_X1 _13129_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_A ), .A4(fanout_net_10 ), .ZN(_05845_ ) );
OAI22_X1 _13130_ ( .A1(_05843_ ), .A2(_05844_ ), .B1(_05525_ ), .B2(_05845_ ), .ZN(_05846_ ) );
AOI22_X1 _13131_ ( .A1(_04359_ ), .A2(\EXU.pc_i [30] ), .B1(\EXU.r1_i [30] ), .B2(_05528_ ), .ZN(_05847_ ) );
NAND2_X1 _13132_ ( .A1(_05846_ ), .A2(_05847_ ), .ZN(_05848_ ) );
BUF_X4 _13133_ ( .A(_05534_ ), .Z(_05849_ ) );
BUF_X2 _13134_ ( .A(_05585_ ), .Z(_05850_ ) );
NAND2_X1 _13135_ ( .A1(_05089_ ), .A2(_05850_ ), .ZN(_05851_ ) );
NOR2_X2 _13136_ ( .A1(_05590_ ), .A2(_05809_ ), .ZN(_05852_ ) );
AND2_X1 _13137_ ( .A1(_05622_ ), .A2(_05625_ ), .ZN(_05853_ ) );
NOR2_X4 _13138_ ( .A1(_05853_ ), .A2(_05626_ ), .ZN(_05854_ ) );
INV_X1 _13139_ ( .A(_05854_ ), .ZN(_05855_ ) );
BUF_X4 _13140_ ( .A(_05855_ ), .Z(_05856_ ) );
NOR2_X1 _13141_ ( .A1(_05612_ ), .A2(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ), .ZN(_05857_ ) );
NOR2_X1 _13142_ ( .A1(_05592_ ), .A2(_05596_ ), .ZN(_05858_ ) );
XOR2_X1 _13143_ ( .A(_05858_ ), .B(_05616_ ), .Z(_05859_ ) );
INV_X1 _13144_ ( .A(_05859_ ), .ZN(_05860_ ) );
AOI21_X1 _13145_ ( .A(_05857_ ), .B1(_05860_ ), .B2(_05521_ ), .ZN(_05861_ ) );
AND2_X1 _13146_ ( .A1(_05613_ ), .A2(_05616_ ), .ZN(_05862_ ) );
XOR2_X2 _13147_ ( .A(_05862_ ), .B(_05618_ ), .Z(_05863_ ) );
MUX2_X1 _13148_ ( .A(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ), .B(_05861_ ), .S(_05863_ ), .Z(_05864_ ) );
XOR2_X1 _13149_ ( .A(_05619_ ), .B(_05621_ ), .Z(_05865_ ) );
BUF_X4 _13150_ ( .A(_05865_ ), .Z(_05866_ ) );
NAND2_X1 _13151_ ( .A1(_05864_ ), .A2(_05866_ ), .ZN(_05867_ ) );
OR2_X2 _13152_ ( .A1(_05866_ ), .A2(_05521_ ), .ZN(_05868_ ) );
AOI21_X1 _13153_ ( .A(_05856_ ), .B1(_05867_ ), .B2(_05868_ ), .ZN(_05869_ ) );
NOR2_X2 _13154_ ( .A1(_05854_ ), .A2(_05521_ ), .ZN(_05870_ ) );
NOR2_X2 _13155_ ( .A1(_05870_ ), .A2(_05626_ ), .ZN(_05871_ ) );
BUF_X2 _13156_ ( .A(_05590_ ), .Z(_05872_ ) );
AND2_X1 _13157_ ( .A1(_05871_ ), .A2(_05872_ ), .ZN(_05873_ ) );
INV_X1 _13158_ ( .A(_05873_ ), .ZN(_05874_ ) );
OR2_X1 _13159_ ( .A1(_05869_ ), .A2(_05874_ ), .ZN(_05875_ ) );
MUX2_X1 _13160_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_A ), .B(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ), .S(_05600_ ), .Z(_05876_ ) );
BUF_X4 _13161_ ( .A(_05603_ ), .Z(_05877_ ) );
BUF_X4 _13162_ ( .A(_05877_ ), .Z(_05878_ ) );
NOR2_X1 _13163_ ( .A1(_05876_ ), .A2(_05878_ ), .ZN(_05879_ ) );
BUF_X4 _13164_ ( .A(_05747_ ), .Z(_05880_ ) );
BUF_X4 _13165_ ( .A(_05607_ ), .Z(_05881_ ) );
AND3_X1 _13166_ ( .A1(_05879_ ), .A2(_05880_ ), .A3(_05881_ ), .ZN(_05882_ ) );
NAND2_X1 _13167_ ( .A1(_05882_ ), .A2(_05769_ ), .ZN(_05883_ ) );
AOI21_X1 _13168_ ( .A(_05852_ ), .B1(_05875_ ), .B2(_05883_ ), .ZN(_05884_ ) );
AND3_X1 _13169_ ( .A1(_05717_ ), .A2(_04657_ ), .A3(_05720_ ), .ZN(_05885_ ) );
NOR3_X1 _13170_ ( .A1(_05885_ ), .A2(_05721_ ), .A3(_05641_ ), .ZN(_05886_ ) );
BUF_X2 _13171_ ( .A(_05572_ ), .Z(_05887_ ) );
BUF_X2 _13172_ ( .A(_05630_ ), .Z(_05888_ ) );
OAI211_X1 _13173_ ( .A(_05887_ ), .B(_05888_ ), .C1(_04736_ ), .C2(_04734_ ), .ZN(_05889_ ) );
BUF_X4 _13174_ ( .A(_05556_ ), .Z(_05890_ ) );
AOI21_X1 _13175_ ( .A(_04737_ ), .B1(_05889_ ), .B2(_05890_ ), .ZN(_05891_ ) );
BUF_X2 _13176_ ( .A(_05634_ ), .Z(_05892_ ) );
AND4_X1 _13177_ ( .A1(_05844_ ), .A2(_05892_ ), .A3(_04731_ ), .A4(_04733_ ), .ZN(_05893_ ) );
OR2_X1 _13178_ ( .A1(_05891_ ), .A2(_05893_ ), .ZN(_05894_ ) );
NAND2_X1 _13179_ ( .A1(_05750_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_20_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05895_ ) );
OAI211_X1 _13180_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_19_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(_05728_ ), .C1(_04984_ ), .C2(_05611_ ), .ZN(_05896_ ) );
NAND2_X1 _13181_ ( .A1(_05895_ ), .A2(_05896_ ), .ZN(_05897_ ) );
NAND2_X1 _13182_ ( .A1(_05897_ ), .A2(_05774_ ), .ZN(_05898_ ) );
NAND2_X1 _13183_ ( .A1(_05726_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05899_ ) );
OAI211_X1 _13184_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .B(_05728_ ), .C1(_04984_ ), .C2(_05611_ ), .ZN(_05900_ ) );
NAND2_X1 _13185_ ( .A1(_05899_ ), .A2(_05900_ ), .ZN(_05901_ ) );
NAND2_X1 _13186_ ( .A1(_05901_ ), .A2(_05735_ ), .ZN(_05902_ ) );
NAND3_X1 _13187_ ( .A1(_05898_ ), .A2(_05902_ ), .A3(_05606_ ), .ZN(_05903_ ) );
NOR2_X1 _13188_ ( .A1(_04908_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_21_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05904_ ) );
AOI21_X1 _13189_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_22_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_04906_ ), .B2(_04907_ ), .ZN(_05905_ ) );
OR3_X1 _13190_ ( .A1(_05904_ ), .A2(_05602_ ), .A3(_05905_ ), .ZN(_05906_ ) );
NAND2_X1 _13191_ ( .A1(_05726_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_24_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05907_ ) );
OAI211_X1 _13192_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_05728_ ), .C1(_04984_ ), .C2(_05611_ ), .ZN(_05908_ ) );
NAND2_X1 _13193_ ( .A1(_05907_ ), .A2(_05908_ ), .ZN(_05909_ ) );
NAND2_X1 _13194_ ( .A1(_05909_ ), .A2(_05603_ ), .ZN(_05910_ ) );
NAND3_X1 _13195_ ( .A1(_05906_ ), .A2(_04996_ ), .A3(_05910_ ), .ZN(_05911_ ) );
AND2_X1 _13196_ ( .A1(_05903_ ), .A2(_05911_ ), .ZN(_05912_ ) );
OR2_X1 _13197_ ( .A1(_05912_ ), .A2(_05757_ ), .ZN(_05913_ ) );
INV_X2 _13198_ ( .A(_04954_ ), .ZN(_05914_ ) );
NAND2_X1 _13199_ ( .A1(_05750_ ), .A2(_04944_ ), .ZN(_05915_ ) );
OAI211_X1 _13200_ ( .A(_05915_ ), .B(_05735_ ), .C1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .C2(_05781_ ), .ZN(_05916_ ) );
OAI211_X1 _13201_ ( .A(_04951_ ), .B(_05785_ ), .C1(_05759_ ), .C2(_05760_ ), .ZN(_05917_ ) );
OAI211_X1 _13202_ ( .A(_05603_ ), .B(_05917_ ), .C1(_04909_ ), .C2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05918_ ) );
AOI21_X1 _13203_ ( .A(_05755_ ), .B1(_05916_ ), .B2(_05918_ ), .ZN(_05919_ ) );
NAND2_X1 _13204_ ( .A1(_05726_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05920_ ) );
OAI211_X1 _13205_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_B_$_MUX__Y_A ), .B(_05728_ ), .C1(_04984_ ), .C2(_05611_ ), .ZN(_05921_ ) );
NAND2_X1 _13206_ ( .A1(_05920_ ), .A2(_05921_ ), .ZN(_05922_ ) );
MUX2_X1 _13207_ ( .A(_04999_ ), .B(_05922_ ), .S(_05735_ ), .Z(_05923_ ) );
BUF_X4 _13208_ ( .A(_04996_ ), .Z(_05924_ ) );
AOI21_X1 _13209_ ( .A(_05919_ ), .B1(_05923_ ), .B2(_05924_ ), .ZN(_05925_ ) );
NAND2_X1 _13210_ ( .A1(_05925_ ), .A2(_05757_ ), .ZN(_05926_ ) );
AND3_X1 _13211_ ( .A1(_05913_ ), .A2(_05914_ ), .A3(_05926_ ), .ZN(_05927_ ) );
BUF_X4 _13212_ ( .A(_05750_ ), .Z(_05928_ ) );
NAND2_X1 _13213_ ( .A1(_05928_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_4_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05929_ ) );
OAI211_X1 _13214_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_3_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(_05785_ ), .C1(_05759_ ), .C2(_05760_ ), .ZN(_05930_ ) );
NAND3_X1 _13215_ ( .A1(_05929_ ), .A2(_05877_ ), .A3(_05930_ ), .ZN(_05931_ ) );
MUX2_X1 _13216_ ( .A(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_A ), .B(\EXU.xrd_o_$_SDFFCE_PP0P__Q_2_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .S(_05928_ ), .Z(_05932_ ) );
OAI211_X1 _13217_ ( .A(_05607_ ), .B(_05931_ ), .C1(_05932_ ), .C2(_05878_ ), .ZN(_05933_ ) );
BUF_X2 _13218_ ( .A(_05606_ ), .Z(_05934_ ) );
NAND2_X1 _13219_ ( .A1(_05781_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_6_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05935_ ) );
OAI211_X1 _13220_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_5_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(_05785_ ), .C1(_05759_ ), .C2(_05760_ ), .ZN(_05936_ ) );
NAND2_X1 _13221_ ( .A1(_05935_ ), .A2(_05936_ ), .ZN(_05937_ ) );
BUF_X4 _13222_ ( .A(_05735_ ), .Z(_05938_ ) );
NAND2_X1 _13223_ ( .A1(_05937_ ), .A2(_05938_ ), .ZN(_05939_ ) );
NAND2_X1 _13224_ ( .A1(_05928_ ), .A2(_04794_ ), .ZN(_05940_ ) );
OAI211_X1 _13225_ ( .A(_05940_ ), .B(_05604_ ), .C1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ), .C2(_05928_ ), .ZN(_05941_ ) );
AND2_X1 _13226_ ( .A1(_05939_ ), .A2(_05941_ ), .ZN(_05942_ ) );
OAI21_X1 _13227_ ( .A(_05933_ ), .B1(_05934_ ), .B2(_05942_ ), .ZN(_05943_ ) );
AND3_X1 _13228_ ( .A1(_04906_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_11_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A3(_05728_ ), .ZN(_05944_ ) );
AOI21_X1 _13229_ ( .A(_04752_ ), .B1(_04906_ ), .B2(_05785_ ), .ZN(_05945_ ) );
OR3_X1 _13230_ ( .A1(_05944_ ), .A2(_05945_ ), .A3(_04901_ ), .ZN(_05946_ ) );
OAI211_X1 _13231_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ), .B(_05785_ ), .C1(_05759_ ), .C2(_05760_ ), .ZN(_05947_ ) );
OAI211_X1 _13232_ ( .A(_05784_ ), .B(_05947_ ), .C1(_04909_ ), .C2(_04825_ ), .ZN(_05948_ ) );
AND3_X1 _13233_ ( .A1(_05946_ ), .A2(_05606_ ), .A3(_05948_ ), .ZN(_05949_ ) );
NAND2_X1 _13234_ ( .A1(_05781_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_16_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_05950_ ) );
OAI211_X1 _13235_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B(_05785_ ), .C1(_05759_ ), .C2(_05760_ ), .ZN(_05951_ ) );
NAND2_X1 _13236_ ( .A1(_05950_ ), .A2(_05951_ ), .ZN(_05952_ ) );
NAND2_X1 _13237_ ( .A1(_05952_ ), .A2(_05604_ ), .ZN(_05953_ ) );
NAND2_X1 _13238_ ( .A1(_05781_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05954_ ) );
OAI211_X1 _13239_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_13_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(_05785_ ), .C1(_05759_ ), .C2(_05760_ ), .ZN(_05955_ ) );
NAND2_X1 _13240_ ( .A1(_05954_ ), .A2(_05955_ ), .ZN(_05956_ ) );
NAND2_X1 _13241_ ( .A1(_05956_ ), .A2(_05938_ ), .ZN(_05957_ ) );
AOI21_X1 _13242_ ( .A(_05606_ ), .B1(_05953_ ), .B2(_05957_ ), .ZN(_05958_ ) );
OR2_X1 _13243_ ( .A1(_05949_ ), .A2(_05958_ ), .ZN(_05959_ ) );
BUF_X4 _13244_ ( .A(_04886_ ), .Z(_05960_ ) );
MUX2_X1 _13245_ ( .A(_05943_ ), .B(_05959_ ), .S(_05960_ ), .Z(_05961_ ) );
AOI211_X1 _13246_ ( .A(_05767_ ), .B(_05927_ ), .C1(_05769_ ), .C2(_05961_ ), .ZN(_05962_ ) );
NOR4_X1 _13247_ ( .A1(_05884_ ), .A2(_05886_ ), .A3(_05894_ ), .A4(_05962_ ), .ZN(_05963_ ) );
AOI21_X1 _13248_ ( .A(_05849_ ), .B1(_05851_ ), .B2(_05963_ ), .ZN(_05964_ ) );
AND2_X1 _13249_ ( .A1(_05098_ ), .A2(_05039_ ), .ZN(_05965_ ) );
NAND2_X1 _13250_ ( .A1(_05843_ ), .A2(_05044_ ), .ZN(_05966_ ) );
BUF_X2 _13251_ ( .A(_05817_ ), .Z(_05967_ ) );
BUF_X2 _13252_ ( .A(_05531_ ), .Z(_05968_ ) );
NAND3_X1 _13253_ ( .A1(_05967_ ), .A2(_05968_ ), .A3(\EXU.imm_i [30] ), .ZN(_05969_ ) );
BUF_X2 _13254_ ( .A(_04387_ ), .Z(_05970_ ) );
BUF_X2 _13255_ ( .A(_04388_ ), .Z(_05971_ ) );
NAND3_X1 _13256_ ( .A1(_05970_ ), .A2(\EXU.ls_rdata_i [30] ), .A3(_05971_ ), .ZN(_05972_ ) );
NAND3_X1 _13257_ ( .A1(_05966_ ), .A2(_05969_ ), .A3(_05972_ ), .ZN(_05973_ ) );
OR3_X2 _13258_ ( .A1(_05964_ ), .A2(_05965_ ), .A3(_05973_ ), .ZN(_05974_ ) );
MUX2_X2 _13259_ ( .A(_05848_ ), .B(_05974_ ), .S(_05822_ ), .Z(_05975_ ) );
NAND2_X1 _13260_ ( .A1(_05975_ ), .A2(_05825_ ), .ZN(_05976_ ) );
BUF_X4 _13261_ ( .A(_05050_ ), .Z(_05977_ ) );
NAND3_X1 _13262_ ( .A1(_04377_ ), .A2(_05977_ ), .A3(_05848_ ), .ZN(_05978_ ) );
AOI21_X1 _13263_ ( .A(_05515_ ), .B1(_05976_ ), .B2(_05978_ ), .ZN(_05979_ ) );
MUX2_X1 _13264_ ( .A(\EXU.xrd_o [30] ), .B(_05979_ ), .S(_04400_ ), .Z(_00242_ ) );
INV_X1 _13265_ ( .A(_04336_ ), .ZN(_05980_ ) );
BUF_X4 _13266_ ( .A(_05980_ ), .Z(_05981_ ) );
OR2_X1 _13267_ ( .A1(_04353_ ), .A2(\EXU.imm_i [11] ), .ZN(_05982_ ) );
NAND2_X1 _13268_ ( .A1(_05982_ ), .A2(_05980_ ), .ZN(_05983_ ) );
BUF_X2 _13269_ ( .A(_04349_ ), .Z(_05984_ ) );
AND3_X1 _13270_ ( .A1(_04352_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_10_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05984_ ), .ZN(_05985_ ) );
OAI221_X1 _13271_ ( .A(_05829_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_10_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05981_ ), .C1(_05983_ ), .C2(_05985_ ), .ZN(_05986_ ) );
BUF_X4 _13272_ ( .A(_05832_ ), .Z(_05987_ ) );
BUF_X4 _13273_ ( .A(_04345_ ), .Z(_05988_ ) );
BUF_X4 _13274_ ( .A(_05988_ ), .Z(_05989_ ) );
NAND4_X1 _13275_ ( .A1(_05987_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_10_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_05989_ ), .ZN(_05990_ ) );
NAND2_X1 _13276_ ( .A1(_05986_ ), .A2(_05990_ ), .ZN(_05991_ ) );
INV_X1 _13277_ ( .A(_04350_ ), .ZN(_05992_ ) );
BUF_X4 _13278_ ( .A(_05992_ ), .Z(_05993_ ) );
MUX2_X1 _13279_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_10_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ), .B(_05991_ ), .S(_05993_ ), .Z(_05994_ ) );
BUF_X4 _13280_ ( .A(_05557_ ), .Z(_05995_ ) );
BUF_X4 _13281_ ( .A(_05995_ ), .Z(_05996_ ) );
NAND4_X1 _13282_ ( .A1(_04973_ ), .A2(fanout_net_6 ), .A3(fanout_net_5 ), .A4(fanout_net_10 ), .ZN(_05997_ ) );
AOI22_X1 _13283_ ( .A1(_05994_ ), .A2(_04973_ ), .B1(_05996_ ), .B2(_05997_ ), .ZN(_05998_ ) );
BUF_X4 _13284_ ( .A(_05046_ ), .Z(_05999_ ) );
NAND3_X1 _13285_ ( .A1(_05045_ ), .A2(\EXU.pc_i [21] ), .A3(_05999_ ), .ZN(_06000_ ) );
INV_X1 _13286_ ( .A(_04716_ ), .ZN(_06001_ ) );
BUF_X4 _13287_ ( .A(_06001_ ), .Z(_06002_ ) );
BUF_X4 _13288_ ( .A(_06002_ ), .Z(_06003_ ) );
OAI21_X1 _13289_ ( .A(_06000_ ), .B1(_04973_ ), .B2(_06003_ ), .ZN(_06004_ ) );
OAI211_X1 _13290_ ( .A(_04371_ ), .B(_04374_ ), .C1(_05998_ ), .C2(_06004_ ), .ZN(_06005_ ) );
BUF_X2 _13291_ ( .A(_04389_ ), .Z(_06006_ ) );
BUF_X2 _13292_ ( .A(_06006_ ), .Z(_06007_ ) );
AND2_X1 _13293_ ( .A1(_05817_ ), .A2(_05531_ ), .ZN(_06008_ ) );
BUF_X4 _13294_ ( .A(_06008_ ), .Z(_06009_ ) );
AOI22_X1 _13295_ ( .A1(_06007_ ), .A2(\EXU.ls_rdata_i [21] ), .B1(_06009_ ), .B2(\EXU.imm_i [21] ), .ZN(_06010_ ) );
BUF_X4 _13296_ ( .A(_05814_ ), .Z(_06011_ ) );
BUF_X4 _13297_ ( .A(_06011_ ), .Z(_06012_ ) );
OAI21_X1 _13298_ ( .A(_06010_ ), .B1(_05994_ ), .B2(_06012_ ), .ZN(_06013_ ) );
BUF_X4 _13299_ ( .A(_05535_ ), .Z(_06014_ ) );
BUF_X4 _13300_ ( .A(_05585_ ), .Z(_06015_ ) );
NAND2_X1 _13301_ ( .A1(_05114_ ), .A2(_06015_ ), .ZN(_06016_ ) );
INV_X1 _13302_ ( .A(_04689_ ), .ZN(_06017_ ) );
AND2_X1 _13303_ ( .A1(_05682_ ), .A2(_04707_ ), .ZN(_06018_ ) );
INV_X1 _13304_ ( .A(_06018_ ), .ZN(_06019_ ) );
AOI21_X1 _13305_ ( .A(_06017_ ), .B1(_06019_ ), .B2(_05702_ ), .ZN(_06020_ ) );
NOR2_X1 _13306_ ( .A1(_06020_ ), .A2(_05686_ ), .ZN(_06021_ ) );
XNOR2_X1 _13307_ ( .A(_06021_ ), .B(_04688_ ), .ZN(_06022_ ) );
BUF_X2 _13308_ ( .A(_05639_ ), .Z(_06023_ ) );
NAND2_X1 _13309_ ( .A1(_06022_ ), .A2(_06023_ ), .ZN(_06024_ ) );
AOI21_X1 _13310_ ( .A(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ), .B1(_05863_ ), .B2(_05859_ ), .ZN(_06025_ ) );
INV_X1 _13311_ ( .A(_05866_ ), .ZN(_06026_ ) );
BUF_X2 _13312_ ( .A(_06026_ ), .Z(_06027_ ) );
AND2_X1 _13313_ ( .A1(_06025_ ), .A2(_06027_ ), .ZN(_06028_ ) );
OAI211_X1 _13314_ ( .A(_05871_ ), .B(_05872_ ), .C1(_06028_ ), .C2(_05856_ ), .ZN(_06029_ ) );
BUF_X4 _13315_ ( .A(_05802_ ), .Z(_06030_ ) );
NOR2_X1 _13316_ ( .A1(_05601_ ), .A2(\EXU.r1_i [25] ), .ZN(_06031_ ) );
BUF_X8 _13317_ ( .A(_05597_ ), .Z(_06032_ ) );
BUF_X8 _13318_ ( .A(_06032_ ), .Z(_06033_ ) );
BUF_X8 _13319_ ( .A(_05598_ ), .Z(_06034_ ) );
BUF_X8 _13320_ ( .A(_06034_ ), .Z(_06035_ ) );
NOR3_X1 _13321_ ( .A1(_06033_ ), .A2(\EXU.r1_i [26] ), .A3(_06035_ ), .ZN(_06036_ ) );
OR3_X1 _13322_ ( .A1(_06031_ ), .A2(_05877_ ), .A3(_06036_ ), .ZN(_06037_ ) );
OR3_X1 _13323_ ( .A1(_06033_ ), .A2(\EXU.r1_i [28] ), .A3(_06035_ ), .ZN(_06038_ ) );
BUF_X4 _13324_ ( .A(_05604_ ), .Z(_06039_ ) );
BUF_X4 _13325_ ( .A(_05601_ ), .Z(_06040_ ) );
OAI211_X1 _13326_ ( .A(_06038_ ), .B(_06039_ ), .C1(\EXU.r1_i [27] ), .C2(_06040_ ), .ZN(_06041_ ) );
AOI21_X1 _13327_ ( .A(_06030_ ), .B1(_06037_ ), .B2(_06041_ ), .ZN(_06042_ ) );
NOR2_X1 _13328_ ( .A1(_05600_ ), .A2(\EXU.r1_i [23] ), .ZN(_06043_ ) );
NOR3_X1 _13329_ ( .A1(_06033_ ), .A2(\EXU.r1_i [24] ), .A3(_06035_ ), .ZN(_06044_ ) );
OAI21_X1 _13330_ ( .A(_06039_ ), .B1(_06043_ ), .B2(_06044_ ), .ZN(_06045_ ) );
BUF_X8 _13331_ ( .A(_06033_ ), .Z(_06046_ ) );
BUF_X2 _13332_ ( .A(_06034_ ), .Z(_06047_ ) );
OR3_X1 _13333_ ( .A1(_06046_ ), .A2(_04785_ ), .A3(_06047_ ), .ZN(_06048_ ) );
BUF_X4 _13334_ ( .A(_05784_ ), .Z(_06049_ ) );
BUF_X8 _13335_ ( .A(_06035_ ), .Z(_06050_ ) );
OAI21_X1 _13336_ ( .A(\EXU.r1_i [21] ), .B1(_06046_ ), .B2(_06050_ ), .ZN(_06051_ ) );
NAND3_X1 _13337_ ( .A1(_06048_ ), .A2(_06049_ ), .A3(_06051_ ), .ZN(_06052_ ) );
AND3_X1 _13338_ ( .A1(_06045_ ), .A2(_05934_ ), .A3(_06052_ ), .ZN(_06053_ ) );
OAI21_X1 _13339_ ( .A(_05880_ ), .B1(_06042_ ), .B2(_06053_ ), .ZN(_06054_ ) );
OAI211_X1 _13340_ ( .A(\EXU.r1_i [31] ), .B(_05877_ ), .C1(_06046_ ), .C2(_06050_ ), .ZN(_06055_ ) );
OR3_X1 _13341_ ( .A1(_06032_ ), .A2(_05844_ ), .A3(_06034_ ), .ZN(_06056_ ) );
OAI21_X1 _13342_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_2_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_06033_ ), .B2(_06035_ ), .ZN(_06057_ ) );
NAND2_X1 _13343_ ( .A1(_06056_ ), .A2(_06057_ ), .ZN(_06058_ ) );
OAI21_X1 _13344_ ( .A(_06055_ ), .B1(_06058_ ), .B2(_06039_ ), .ZN(_06059_ ) );
BUF_X2 _13345_ ( .A(_05757_ ), .Z(_06060_ ) );
NAND3_X1 _13346_ ( .A1(_06059_ ), .A2(_06060_ ), .A3(_05881_ ), .ZN(_06061_ ) );
AND2_X1 _13347_ ( .A1(_06054_ ), .A2(_06061_ ), .ZN(_06062_ ) );
BUF_X2 _13348_ ( .A(_05914_ ), .Z(_06063_ ) );
OAI21_X1 _13349_ ( .A(_06029_ ), .B1(_06062_ ), .B2(_06063_ ), .ZN(_06064_ ) );
INV_X1 _13350_ ( .A(_05852_ ), .ZN(_06065_ ) );
BUF_X4 _13351_ ( .A(_06065_ ), .Z(_06066_ ) );
NAND2_X1 _13352_ ( .A1(_06064_ ), .A2(_06066_ ), .ZN(_06067_ ) );
NAND3_X1 _13353_ ( .A1(_04824_ ), .A2(\EXU.r1_i [21] ), .A3(_04826_ ), .ZN(_06068_ ) );
AND3_X1 _13354_ ( .A1(_05887_ ), .A2(_05888_ ), .A3(_06068_ ), .ZN(_06069_ ) );
OAI22_X1 _13355_ ( .A1(_06069_ ), .A2(_05555_ ), .B1(\EXU.r1_i [21] ), .B2(_04829_ ), .ZN(_06070_ ) );
BUF_X4 _13356_ ( .A(_05635_ ), .Z(_06071_ ) );
MUX2_X1 _13357_ ( .A(_04827_ ), .B(_06070_ ), .S(_06071_ ), .Z(_06072_ ) );
NAND2_X1 _13358_ ( .A1(_05773_ ), .A2(_05735_ ), .ZN(_06073_ ) );
NAND3_X1 _13359_ ( .A1(_05783_ ), .A2(_05603_ ), .A3(_05786_ ), .ZN(_06074_ ) );
NAND3_X1 _13360_ ( .A1(_06073_ ), .A2(_06030_ ), .A3(_06074_ ), .ZN(_06075_ ) );
OAI211_X1 _13361_ ( .A(_05780_ ), .B(_05784_ ), .C1(_04755_ ), .C2(_05928_ ), .ZN(_06076_ ) );
BUF_X4 _13362_ ( .A(_05924_ ), .Z(_06077_ ) );
OAI21_X1 _13363_ ( .A(_05604_ ), .B1(_05741_ ), .B2(_05742_ ), .ZN(_06078_ ) );
NAND3_X1 _13364_ ( .A1(_06076_ ), .A2(_06077_ ), .A3(_06078_ ), .ZN(_06079_ ) );
AOI211_X1 _13365_ ( .A(_05914_ ), .B(_06060_ ), .C1(_06075_ ), .C2(_06079_ ), .ZN(_06080_ ) );
BUF_X2 _13366_ ( .A(_05960_ ), .Z(_06081_ ) );
NAND2_X1 _13367_ ( .A1(_05730_ ), .A2(_05784_ ), .ZN(_06082_ ) );
NAND2_X1 _13368_ ( .A1(_05750_ ), .A2(_04936_ ), .ZN(_06083_ ) );
OAI211_X1 _13369_ ( .A(_06083_ ), .B(_05603_ ), .C1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_24_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .C2(_05781_ ), .ZN(_06084_ ) );
NAND2_X1 _13370_ ( .A1(_06082_ ), .A2(_06084_ ), .ZN(_06085_ ) );
OAI21_X1 _13371_ ( .A(_05784_ ), .B1(_05738_ ), .B2(_05739_ ), .ZN(_06086_ ) );
NAND3_X1 _13372_ ( .A1(_05732_ ), .A2(_05603_ ), .A3(_05733_ ), .ZN(_06087_ ) );
AND2_X1 _13373_ ( .A1(_06086_ ), .A2(_06087_ ), .ZN(_06088_ ) );
MUX2_X1 _13374_ ( .A(_06085_ ), .B(_06088_ ), .S(_05802_ ), .Z(_06089_ ) );
AOI211_X1 _13375_ ( .A(_05767_ ), .B(_06080_ ), .C1(_06081_ ), .C2(_06089_ ), .ZN(_06090_ ) );
BUF_X2 _13376_ ( .A(_05807_ ), .Z(_06091_ ) );
NAND2_X1 _13377_ ( .A1(_05762_ ), .A2(_05774_ ), .ZN(_06092_ ) );
NAND2_X1 _13378_ ( .A1(_05750_ ), .A2(_04951_ ), .ZN(_06093_ ) );
OAI211_X1 _13379_ ( .A(_06093_ ), .B(_05735_ ), .C1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_26_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .C2(_05781_ ), .ZN(_06094_ ) );
AND3_X1 _13380_ ( .A1(_06092_ ), .A2(_05606_ ), .A3(_06094_ ), .ZN(_06095_ ) );
BUF_X4 _13381_ ( .A(_05755_ ), .Z(_06096_ ) );
NOR2_X1 _13382_ ( .A1(_05763_ ), .A2(_06039_ ), .ZN(_06097_ ) );
AOI21_X1 _13383_ ( .A(_06095_ ), .B1(_06096_ ), .B2(_06097_ ), .ZN(_06098_ ) );
BUF_X4 _13384_ ( .A(_05960_ ), .Z(_06099_ ) );
BUF_X4 _13385_ ( .A(_06099_ ), .Z(_06100_ ) );
NOR2_X1 _13386_ ( .A1(_06098_ ), .A2(_06100_ ), .ZN(_06101_ ) );
OAI21_X1 _13387_ ( .A(_06090_ ), .B1(_06091_ ), .B2(_06101_ ), .ZN(_06102_ ) );
AND4_X1 _13388_ ( .A1(_06024_ ), .A2(_06067_ ), .A3(_06072_ ), .A4(_06102_ ), .ZN(_06103_ ) );
AOI21_X1 _13389_ ( .A(_06014_ ), .B1(_06016_ ), .B2(_06103_ ), .ZN(_06104_ ) );
AOI211_X1 _13390_ ( .A(_06013_ ), .B(_06104_ ), .C1(_05211_ ), .C2(_05129_ ), .ZN(_06105_ ) );
BUF_X4 _13391_ ( .A(_04394_ ), .Z(_06106_ ) );
OAI21_X1 _13392_ ( .A(_06005_ ), .B1(_06105_ ), .B2(_06106_ ), .ZN(_06107_ ) );
NAND2_X1 _13393_ ( .A1(_06107_ ), .A2(_05825_ ), .ZN(_06108_ ) );
BUF_X4 _13394_ ( .A(_04376_ ), .Z(_06109_ ) );
OAI211_X1 _13395_ ( .A(_06109_ ), .B(_05290_ ), .C1(_05998_ ), .C2(_06004_ ), .ZN(_06110_ ) );
AOI21_X1 _13396_ ( .A(_05515_ ), .B1(_06108_ ), .B2(_06110_ ), .ZN(_06111_ ) );
MUX2_X1 _13397_ ( .A(\EXU.xrd_o [21] ), .B(_06111_ ), .S(_04400_ ), .Z(_00243_ ) );
AND4_X1 _13398_ ( .A1(\EXU.mtvec_i [20] ), .A2(_04349_ ), .A3(_05052_ ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_06112_ ) );
OAI21_X1 _13399_ ( .A(_05981_ ), .B1(_06112_ ), .B2(_05834_ ), .ZN(_06113_ ) );
AND3_X1 _13400_ ( .A1(_04334_ ), .A2(\EXU.mcause_i [20] ), .A3(_05839_ ), .ZN(_06114_ ) );
INV_X1 _13401_ ( .A(_06114_ ), .ZN(_06115_ ) );
AOI21_X1 _13402_ ( .A(_05516_ ), .B1(_06113_ ), .B2(_06115_ ), .ZN(_06116_ ) );
AND3_X1 _13403_ ( .A1(_05836_ ), .A2(_05831_ ), .A3(\EXU.mepc_i [20] ), .ZN(_06117_ ) );
BUF_X2 _13404_ ( .A(_04352_ ), .Z(_06118_ ) );
AND3_X1 _13405_ ( .A1(_06118_ ), .A2(\EXU.mstatus_i [20] ), .A3(_05988_ ), .ZN(_06119_ ) );
NOR3_X1 _13406_ ( .A1(_06116_ ), .A2(_06117_ ), .A3(_06119_ ), .ZN(_06120_ ) );
NAND4_X1 _13407_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_11_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_06121_ ) );
AOI22_X1 _13408_ ( .A1(_06120_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_11_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_05995_ ), .B2(_06121_ ), .ZN(_06122_ ) );
BUF_X2 _13409_ ( .A(_04343_ ), .Z(_06123_ ) );
NAND3_X1 _13410_ ( .A1(_06123_ ), .A2(\EXU.pc_i [20] ), .A3(_05046_ ), .ZN(_06124_ ) );
OAI21_X1 _13411_ ( .A(_06124_ ), .B1(_04835_ ), .B2(_06002_ ), .ZN(_06125_ ) );
OR2_X1 _13412_ ( .A1(_06122_ ), .A2(_06125_ ), .ZN(_06126_ ) );
NAND2_X1 _13413_ ( .A1(_05133_ ), .A2(_05850_ ), .ZN(_06127_ ) );
NOR3_X1 _13414_ ( .A1(_05774_ ), .A2(_04911_ ), .A3(_05781_ ), .ZN(_06128_ ) );
INV_X1 _13415_ ( .A(_06128_ ), .ZN(_06129_ ) );
NAND2_X1 _13416_ ( .A1(_05922_ ), .A2(_05774_ ), .ZN(_06130_ ) );
OAI211_X1 _13417_ ( .A(_05735_ ), .B(_05917_ ), .C1(_04909_ ), .C2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_06131_ ) );
NAND2_X1 _13418_ ( .A1(_06130_ ), .A2(_06131_ ), .ZN(_06132_ ) );
MUX2_X1 _13419_ ( .A(_06129_ ), .B(_06132_ ), .S(_05606_ ), .Z(_06133_ ) );
OAI21_X1 _13420_ ( .A(_05914_ ), .B1(_06133_ ), .B2(_06060_ ), .ZN(_06134_ ) );
AND2_X1 _13421_ ( .A1(_06134_ ), .A2(_05565_ ), .ZN(_06135_ ) );
NAND2_X1 _13422_ ( .A1(_05928_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_26_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_06136_ ) );
OAI211_X1 _13423_ ( .A(_06136_ ), .B(_05877_ ), .C1(_04936_ ), .C2(_05928_ ), .ZN(_06137_ ) );
OAI211_X1 _13424_ ( .A(_06137_ ), .B(_05924_ ), .C1(_05878_ ), .C2(_05909_ ), .ZN(_06138_ ) );
NAND3_X1 _13425_ ( .A1(_05895_ ), .A2(_05938_ ), .A3(_05896_ ), .ZN(_06139_ ) );
NOR2_X1 _13426_ ( .A1(_05904_ ), .A2(_05905_ ), .ZN(_06140_ ) );
OAI211_X1 _13427_ ( .A(_05802_ ), .B(_06139_ ), .C1(_06140_ ), .C2(_06049_ ), .ZN(_06141_ ) );
AND2_X1 _13428_ ( .A1(_06138_ ), .A2(_06141_ ), .ZN(_06142_ ) );
OR3_X1 _13429_ ( .A1(_05944_ ), .A2(_05774_ ), .A3(_05945_ ), .ZN(_06143_ ) );
BUF_X4 _13430_ ( .A(_05938_ ), .Z(_06144_ ) );
OAI211_X1 _13431_ ( .A(_06143_ ), .B(_05802_ ), .C1(_06144_ ), .C2(_05956_ ), .ZN(_06145_ ) );
NAND3_X1 _13432_ ( .A1(_05950_ ), .A2(_05938_ ), .A3(_05951_ ), .ZN(_06146_ ) );
OAI211_X1 _13433_ ( .A(_06146_ ), .B(_05924_ ), .C1(_05901_ ), .C2(_06049_ ), .ZN(_06147_ ) );
AND2_X1 _13434_ ( .A1(_06145_ ), .A2(_06147_ ), .ZN(_06148_ ) );
MUX2_X1 _13435_ ( .A(_06142_ ), .B(_06148_ ), .S(_05804_ ), .Z(_06149_ ) );
OAI21_X1 _13436_ ( .A(_06135_ ), .B1(_06063_ ), .B2(_06149_ ), .ZN(_06150_ ) );
INV_X1 _13437_ ( .A(_05857_ ), .ZN(_06151_ ) );
NOR2_X1 _13438_ ( .A1(_05859_ ), .A2(_06151_ ), .ZN(_06152_ ) );
INV_X1 _13439_ ( .A(_05863_ ), .ZN(_06153_ ) );
AOI21_X1 _13440_ ( .A(_06152_ ), .B1(_06153_ ), .B2(_05521_ ), .ZN(_06154_ ) );
NOR2_X1 _13441_ ( .A1(_06154_ ), .A2(_05866_ ), .ZN(_06155_ ) );
OAI211_X2 _13442_ ( .A(_05872_ ), .B(_05871_ ), .C1(_06155_ ), .C2(_05856_ ), .ZN(_06156_ ) );
NAND2_X1 _13443_ ( .A1(_05876_ ), .A2(_05877_ ), .ZN(_06157_ ) );
INV_X1 _13444_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_2_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_06158_ ) );
OR3_X4 _13445_ ( .A1(_06033_ ), .A2(_06158_ ), .A3(_06035_ ), .ZN(_06159_ ) );
BUF_X4 _13446_ ( .A(_06032_ ), .Z(_06160_ ) );
OAI21_X1 _13447_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_3_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_06160_ ), .B2(_06047_ ), .ZN(_06161_ ) );
NAND2_X2 _13448_ ( .A1(_06159_ ), .A2(_06161_ ), .ZN(_06162_ ) );
NAND2_X2 _13449_ ( .A1(_06162_ ), .A2(_06049_ ), .ZN(_06163_ ) );
AND4_X1 _13450_ ( .A1(_05757_ ), .A2(_06157_ ), .A3(_05607_ ), .A4(_06163_ ), .ZN(_06164_ ) );
NOR2_X4 _13451_ ( .A1(_05600_ ), .A2(\EXU.r1_i [26] ), .ZN(_06165_ ) );
NOR3_X2 _13452_ ( .A1(_06032_ ), .A2(\EXU.r1_i [27] ), .A3(_06034_ ), .ZN(_06166_ ) );
OAI21_X1 _13453_ ( .A(_05602_ ), .B1(_06165_ ), .B2(_06166_ ), .ZN(_06167_ ) );
OR3_X1 _13454_ ( .A1(_05597_ ), .A2(_04814_ ), .A3(_05598_ ), .ZN(_06168_ ) );
OAI21_X1 _13455_ ( .A(\EXU.r1_i [24] ), .B1(_06032_ ), .B2(_06034_ ), .ZN(_06169_ ) );
NAND3_X1 _13456_ ( .A1(_06168_ ), .A2(_04901_ ), .A3(_06169_ ), .ZN(_06170_ ) );
AND2_X2 _13457_ ( .A1(_06167_ ), .A2(_06170_ ), .ZN(_06171_ ) );
NOR2_X1 _13458_ ( .A1(_05599_ ), .A2(\EXU.r1_i [20] ), .ZN(_06172_ ) );
NOR3_X2 _13459_ ( .A1(_06032_ ), .A2(\EXU.r1_i [21] ), .A3(_06034_ ), .ZN(_06173_ ) );
OR3_X4 _13460_ ( .A1(_06172_ ), .A2(_05602_ ), .A3(_06173_ ), .ZN(_06174_ ) );
OAI21_X1 _13461_ ( .A(_04785_ ), .B1(_06032_ ), .B2(_06034_ ), .ZN(_06175_ ) );
INV_X4 _13462_ ( .A(_05600_ ), .ZN(_06176_ ) );
OAI211_X2 _13463_ ( .A(_05602_ ), .B(_06175_ ), .C1(_06176_ ), .C2(\EXU.r1_i [23] ), .ZN(_06177_ ) );
NAND2_X2 _13464_ ( .A1(_06174_ ), .A2(_06177_ ), .ZN(_06178_ ) );
MUX2_X2 _13465_ ( .A(_06171_ ), .B(_06178_ ), .S(_04892_ ), .Z(_06179_ ) );
AOI21_X1 _13466_ ( .A(_06164_ ), .B1(_06179_ ), .B2(_05880_ ), .ZN(_06180_ ) );
BUF_X2 _13467_ ( .A(_05914_ ), .Z(_06181_ ) );
OAI21_X1 _13468_ ( .A(_06156_ ), .B1(_06180_ ), .B2(_06181_ ), .ZN(_06182_ ) );
NAND2_X1 _13469_ ( .A1(_06182_ ), .A2(_06066_ ), .ZN(_06183_ ) );
OAI211_X1 _13470_ ( .A(_05887_ ), .B(_05888_ ), .C1(_04835_ ), .C2(_04833_ ), .ZN(_06184_ ) );
AOI21_X1 _13471_ ( .A(_04836_ ), .B1(_06184_ ), .B2(_05890_ ), .ZN(_06185_ ) );
BUF_X4 _13472_ ( .A(_05892_ ), .Z(_06186_ ) );
AOI21_X1 _13473_ ( .A(_06185_ ), .B1(_04834_ ), .B2(_06186_ ), .ZN(_06187_ ) );
NOR3_X1 _13474_ ( .A1(_06018_ ), .A2(_04689_ ), .A3(_05703_ ), .ZN(_06188_ ) );
OR3_X1 _13475_ ( .A1(_06020_ ), .A2(_05640_ ), .A3(_06188_ ), .ZN(_06189_ ) );
AND4_X2 _13476_ ( .A1(_06150_ ), .A2(_06183_ ), .A3(_06187_ ), .A4(_06189_ ), .ZN(_06190_ ) );
AOI21_X1 _13477_ ( .A(_05849_ ), .B1(_06127_ ), .B2(_06190_ ), .ZN(_06191_ ) );
AND2_X1 _13478_ ( .A1(_05140_ ), .A2(_05039_ ), .ZN(_06192_ ) );
AOI22_X1 _13479_ ( .A1(_06006_ ), .A2(\EXU.ls_rdata_i [20] ), .B1(_06009_ ), .B2(\EXU.imm_i [20] ), .ZN(_06193_ ) );
OAI21_X1 _13480_ ( .A(_06193_ ), .B1(_06120_ ), .B2(_06011_ ), .ZN(_06194_ ) );
OR3_X2 _13481_ ( .A1(_06191_ ), .A2(_06192_ ), .A3(_06194_ ), .ZN(_06195_ ) );
MUX2_X1 _13482_ ( .A(_06126_ ), .B(_06195_ ), .S(_05822_ ), .Z(_06196_ ) );
NAND2_X1 _13483_ ( .A1(_06196_ ), .A2(_05825_ ), .ZN(_06197_ ) );
NAND3_X1 _13484_ ( .A1(_04377_ ), .A2(_05977_ ), .A3(_06126_ ), .ZN(_06198_ ) );
AOI21_X1 _13485_ ( .A(_05515_ ), .B1(_06197_ ), .B2(_06198_ ), .ZN(_06199_ ) );
MUX2_X1 _13486_ ( .A(\EXU.xrd_o [20] ), .B(_06199_ ), .S(_04400_ ), .Z(_00244_ ) );
NAND2_X1 _13487_ ( .A1(\EXU.imm_i [11] ), .A2(\EXU.imm_i [0] ), .ZN(_06200_ ) );
NOR2_X1 _13488_ ( .A1(_04353_ ), .A2(_06200_ ), .ZN(_06201_ ) );
NOR2_X1 _13489_ ( .A1(_06201_ ), .A2(_04350_ ), .ZN(_06202_ ) );
BUF_X2 _13490_ ( .A(_04334_ ), .Z(_06203_ ) );
BUF_X2 _13491_ ( .A(_04335_ ), .Z(_06204_ ) );
NAND3_X1 _13492_ ( .A1(_06203_ ), .A2(\EXU.mcause_i [19] ), .A3(_06204_ ), .ZN(_06205_ ) );
BUF_X4 _13493_ ( .A(_04352_ ), .Z(_06206_ ) );
NAND3_X1 _13494_ ( .A1(_06206_ ), .A2(\EXU.mstatus_i [19] ), .A3(_05988_ ), .ZN(_06207_ ) );
BUF_X4 _13495_ ( .A(_05984_ ), .Z(_06208_ ) );
NAND3_X1 _13496_ ( .A1(_06118_ ), .A2(\EXU.mtvec_i [19] ), .A3(_06208_ ), .ZN(_06209_ ) );
NAND4_X1 _13497_ ( .A1(_06202_ ), .A2(_06205_ ), .A3(_06207_ ), .A4(_06209_ ), .ZN(_06210_ ) );
OAI21_X1 _13498_ ( .A(_06210_ ), .B1(\EXU.mepc_i [19] ), .B2(_05992_ ), .ZN(_06211_ ) );
NAND4_X1 _13499_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_12_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_06212_ ) );
AOI22_X1 _13500_ ( .A1(_06211_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_12_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_05995_ ), .B2(_06212_ ), .ZN(_06213_ ) );
NAND3_X1 _13501_ ( .A1(_06123_ ), .A2(\EXU.pc_i [19] ), .A3(_05046_ ), .ZN(_06214_ ) );
OAI21_X1 _13502_ ( .A(_06214_ ), .B1(_04750_ ), .B2(_06002_ ), .ZN(_06215_ ) );
OR2_X1 _13503_ ( .A1(_06213_ ), .A2(_06215_ ), .ZN(_06216_ ) );
NAND2_X1 _13504_ ( .A1(_05147_ ), .A2(_05850_ ), .ZN(_06217_ ) );
NAND4_X1 _13505_ ( .A1(_06176_ ), .A2(\EXU.r1_i [31] ), .A3(_06096_ ), .A4(_06144_ ), .ZN(_06218_ ) );
MUX2_X1 _13506_ ( .A(\EXU.r1_i [29] ), .B(\EXU.r1_i [30] ), .S(_05600_ ), .Z(_06219_ ) );
NAND2_X1 _13507_ ( .A1(_06219_ ), .A2(_06039_ ), .ZN(_06220_ ) );
OAI211_X1 _13508_ ( .A(_06038_ ), .B(_05938_ ), .C1(\EXU.r1_i [27] ), .C2(_06040_ ), .ZN(_06221_ ) );
AND2_X1 _13509_ ( .A1(_06220_ ), .A2(_06221_ ), .ZN(_06222_ ) );
OAI211_X1 _13510_ ( .A(_05960_ ), .B(_06218_ ), .C1(_06222_ ), .C2(_06077_ ), .ZN(_06223_ ) );
OR3_X1 _13511_ ( .A1(_06031_ ), .A2(_05784_ ), .A3(_06036_ ), .ZN(_06224_ ) );
OR3_X1 _13512_ ( .A1(_06043_ ), .A2(_05774_ ), .A3(_06044_ ), .ZN(_06225_ ) );
NAND3_X1 _13513_ ( .A1(_06224_ ), .A2(_06225_ ), .A3(_05924_ ), .ZN(_06226_ ) );
NOR2_X1 _13514_ ( .A1(_05601_ ), .A2(\EXU.r1_i [19] ), .ZN(_06227_ ) );
NOR3_X1 _13515_ ( .A1(_06033_ ), .A2(\EXU.r1_i [20] ), .A3(_06035_ ), .ZN(_06228_ ) );
OR3_X1 _13516_ ( .A1(_06227_ ), .A2(_05774_ ), .A3(_06228_ ), .ZN(_06229_ ) );
OAI21_X1 _13517_ ( .A(_04973_ ), .B1(_06160_ ), .B2(_06050_ ), .ZN(_06230_ ) );
OAI211_X1 _13518_ ( .A(_05877_ ), .B(_06230_ ), .C1(_06176_ ), .C2(\EXU.r1_i [22] ), .ZN(_06231_ ) );
NAND3_X1 _13519_ ( .A1(_06229_ ), .A2(_05607_ ), .A3(_06231_ ), .ZN(_06232_ ) );
AND2_X1 _13520_ ( .A1(_06226_ ), .A2(_06232_ ), .ZN(_06233_ ) );
OAI21_X1 _13521_ ( .A(_06223_ ), .B1(_06060_ ), .B2(_06233_ ), .ZN(_06234_ ) );
OR2_X1 _13522_ ( .A1(_06234_ ), .A2(_06181_ ), .ZN(_06235_ ) );
NOR2_X1 _13523_ ( .A1(_05863_ ), .A2(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ), .ZN(_06236_ ) );
AND2_X1 _13524_ ( .A1(_06236_ ), .A2(_06027_ ), .ZN(_06237_ ) );
OAI211_X1 _13525_ ( .A(_05871_ ), .B(_05872_ ), .C1(_05856_ ), .C2(_06237_ ), .ZN(_06238_ ) );
AOI21_X1 _13526_ ( .A(_05852_ ), .B1(_06235_ ), .B2(_06238_ ), .ZN(_06239_ ) );
INV_X1 _13527_ ( .A(_04702_ ), .ZN(_06240_ ) );
NAND2_X1 _13528_ ( .A1(_05682_ ), .A2(_04706_ ), .ZN(_06241_ ) );
AOI21_X1 _13529_ ( .A(_06240_ ), .B1(_06241_ ), .B2(_05695_ ), .ZN(_06242_ ) );
NOR2_X1 _13530_ ( .A1(_06242_ ), .A2(_05698_ ), .ZN(_06243_ ) );
XNOR2_X1 _13531_ ( .A(_06243_ ), .B(_04701_ ), .ZN(_06244_ ) );
AND2_X1 _13532_ ( .A1(_06244_ ), .A2(_06023_ ), .ZN(_06245_ ) );
NAND3_X1 _13533_ ( .A1(_04746_ ), .A2(\EXU.r1_i [19] ), .A3(_04748_ ), .ZN(_06246_ ) );
AOI21_X1 _13534_ ( .A(_05555_ ), .B1(_05573_ ), .B2(_06246_ ), .ZN(_06247_ ) );
OAI21_X1 _13535_ ( .A(_05635_ ), .B1(_06247_ ), .B2(_04751_ ), .ZN(_06248_ ) );
OAI21_X1 _13536_ ( .A(_05892_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_12_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B2(_04749_ ), .ZN(_06249_ ) );
AND3_X1 _13537_ ( .A1(_06248_ ), .A2(_04427_ ), .A3(_06249_ ), .ZN(_06250_ ) );
NOR3_X1 _13538_ ( .A1(_05764_ ), .A2(_04886_ ), .A3(_05924_ ), .ZN(_06251_ ) );
OAI21_X1 _13539_ ( .A(_05565_ ), .B1(_06251_ ), .B2(_04954_ ), .ZN(_06252_ ) );
MUX2_X1 _13540_ ( .A(_05737_ ), .B(_05754_ ), .S(_05755_ ), .Z(_06253_ ) );
AND2_X1 _13541_ ( .A1(_04954_ ), .A2(_04885_ ), .ZN(_06254_ ) );
AND3_X1 _13542_ ( .A1(_05740_ ), .A2(_05744_ ), .A3(_05755_ ), .ZN(_06255_ ) );
AOI21_X1 _13543_ ( .A(_05755_ ), .B1(_05782_ ), .B2(_05787_ ), .ZN(_06256_ ) );
NOR2_X1 _13544_ ( .A1(_06255_ ), .A2(_06256_ ), .ZN(_06257_ ) );
AOI221_X4 _13545_ ( .A(_06252_ ), .B1(_05960_ ), .B2(_06253_ ), .C1(_06254_ ), .C2(_06257_ ), .ZN(_06258_ ) );
NOR4_X1 _13546_ ( .A1(_06239_ ), .A2(_06245_ ), .A3(_06250_ ), .A4(_06258_ ), .ZN(_06259_ ) );
AOI21_X1 _13547_ ( .A(_05849_ ), .B1(_06217_ ), .B2(_06259_ ), .ZN(_06260_ ) );
AND2_X1 _13548_ ( .A1(_05152_ ), .A2(_05039_ ), .ZN(_06261_ ) );
AOI22_X1 _13549_ ( .A1(_06006_ ), .A2(\EXU.ls_rdata_i [19] ), .B1(_06008_ ), .B2(\EXU.imm_i [19] ), .ZN(_06262_ ) );
OAI21_X1 _13550_ ( .A(_06262_ ), .B1(_06211_ ), .B2(_06011_ ), .ZN(_06263_ ) );
OR3_X2 _13551_ ( .A1(_06260_ ), .A2(_06261_ ), .A3(_06263_ ), .ZN(_06264_ ) );
MUX2_X2 _13552_ ( .A(_06216_ ), .B(_06264_ ), .S(_05822_ ), .Z(_06265_ ) );
NAND2_X1 _13553_ ( .A1(_06265_ ), .A2(_05825_ ), .ZN(_06266_ ) );
NAND3_X1 _13554_ ( .A1(_04377_ ), .A2(_05977_ ), .A3(_06216_ ), .ZN(_06267_ ) );
AOI21_X1 _13555_ ( .A(_05515_ ), .B1(_06266_ ), .B2(_06267_ ), .ZN(_06268_ ) );
MUX2_X1 _13556_ ( .A(\EXU.xrd_o [19] ), .B(_06268_ ), .S(_04400_ ), .Z(_00245_ ) );
NAND3_X1 _13557_ ( .A1(_06203_ ), .A2(\EXU.mcause_i [18] ), .A3(_06204_ ), .ZN(_06269_ ) );
NAND3_X1 _13558_ ( .A1(_06206_ ), .A2(\EXU.mstatus_i [18] ), .A3(_05989_ ), .ZN(_06270_ ) );
NAND3_X1 _13559_ ( .A1(_06206_ ), .A2(\EXU.mtvec_i [18] ), .A3(_06208_ ), .ZN(_06271_ ) );
NAND4_X1 _13560_ ( .A1(_06202_ ), .A2(_06269_ ), .A3(_06270_ ), .A4(_06271_ ), .ZN(_06272_ ) );
OR2_X1 _13561_ ( .A1(_05992_ ), .A2(\EXU.mepc_i [18] ), .ZN(_06273_ ) );
NAND2_X1 _13562_ ( .A1(_06272_ ), .A2(_06273_ ), .ZN(_06274_ ) );
NAND4_X1 _13563_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_13_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_06275_ ) );
AOI22_X1 _13564_ ( .A1(_06274_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_13_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_05995_ ), .B2(_06275_ ), .ZN(_06276_ ) );
NAND3_X1 _13565_ ( .A1(_06123_ ), .A2(\EXU.pc_i [18] ), .A3(_05046_ ), .ZN(_06277_ ) );
OAI21_X1 _13566_ ( .A(_06277_ ), .B1(_04742_ ), .B2(_06002_ ), .ZN(_06278_ ) );
OR2_X1 _13567_ ( .A1(_06276_ ), .A2(_06278_ ), .ZN(_06279_ ) );
NAND2_X1 _13568_ ( .A1(_05157_ ), .A2(_05850_ ), .ZN(_06280_ ) );
NAND3_X1 _13569_ ( .A1(_05906_ ), .A2(_05607_ ), .A3(_05910_ ), .ZN(_06281_ ) );
NAND3_X1 _13570_ ( .A1(_05916_ ), .A2(_05918_ ), .A3(_05924_ ), .ZN(_06282_ ) );
NAND2_X1 _13571_ ( .A1(_06281_ ), .A2(_06282_ ), .ZN(_06283_ ) );
AOI21_X1 _13572_ ( .A(_05802_ ), .B1(_05898_ ), .B2(_05902_ ), .ZN(_06284_ ) );
AOI21_X1 _13573_ ( .A(_05924_ ), .B1(_05953_ ), .B2(_05957_ ), .ZN(_06285_ ) );
NOR2_X1 _13574_ ( .A1(_06284_ ), .A2(_06285_ ), .ZN(_06286_ ) );
MUX2_X1 _13575_ ( .A(_06283_ ), .B(_06286_ ), .S(_05804_ ), .Z(_06287_ ) );
AND2_X1 _13576_ ( .A1(_06287_ ), .A2(_05807_ ), .ZN(_06288_ ) );
BUF_X4 _13577_ ( .A(_06077_ ), .Z(_06289_ ) );
NOR4_X1 _13578_ ( .A1(_05923_ ), .A2(_05807_ ), .A3(_06099_ ), .A4(_06289_ ), .ZN(_06290_ ) );
OAI21_X1 _13579_ ( .A(_05565_ ), .B1(_06288_ ), .B2(_06290_ ), .ZN(_06291_ ) );
NOR2_X1 _13580_ ( .A1(_05861_ ), .A2(_05863_ ), .ZN(_06292_ ) );
AND2_X1 _13581_ ( .A1(_06292_ ), .A2(_06026_ ), .ZN(_06293_ ) );
OAI211_X1 _13582_ ( .A(_05871_ ), .B(_05872_ ), .C1(_06293_ ), .C2(_05856_ ), .ZN(_06294_ ) );
OR3_X1 _13583_ ( .A1(_06165_ ), .A2(_05604_ ), .A3(_06166_ ), .ZN(_06295_ ) );
NOR2_X1 _13584_ ( .A1(_05601_ ), .A2(_04778_ ), .ZN(_06296_ ) );
NOR3_X4 _13585_ ( .A1(_06046_ ), .A2(_04771_ ), .A3(_06050_ ), .ZN(_06297_ ) );
OAI21_X1 _13586_ ( .A(_05877_ ), .B1(_06296_ ), .B2(_06297_ ), .ZN(_06298_ ) );
NAND3_X1 _13587_ ( .A1(_06295_ ), .A2(_05607_ ), .A3(_06298_ ), .ZN(_06299_ ) );
OAI21_X1 _13588_ ( .A(_06299_ ), .B1(_05879_ ), .B2(_05934_ ), .ZN(_06300_ ) );
OR3_X1 _13589_ ( .A1(_06172_ ), .A2(_05784_ ), .A3(_06173_ ), .ZN(_06301_ ) );
OR3_X1 _13590_ ( .A1(_06160_ ), .A2(\EXU.r1_i [19] ), .A3(_06047_ ), .ZN(_06302_ ) );
OAI211_X1 _13591_ ( .A(_06302_ ), .B(_05938_ ), .C1(\EXU.r1_i [18] ), .C2(_06040_ ), .ZN(_06303_ ) );
AOI21_X1 _13592_ ( .A(_06096_ ), .B1(_06301_ ), .B2(_06303_ ), .ZN(_06304_ ) );
OR3_X1 _13593_ ( .A1(_06160_ ), .A2(\EXU.r1_i [25] ), .A3(_06047_ ), .ZN(_06305_ ) );
OAI211_X1 _13594_ ( .A(_06305_ ), .B(_05877_ ), .C1(\EXU.r1_i [24] ), .C2(_06040_ ), .ZN(_06306_ ) );
OAI211_X1 _13595_ ( .A(_05938_ ), .B(_06175_ ), .C1(_06176_ ), .C2(\EXU.r1_i [23] ), .ZN(_06307_ ) );
AOI21_X1 _13596_ ( .A(_05802_ ), .B1(_06306_ ), .B2(_06307_ ), .ZN(_06308_ ) );
NOR2_X1 _13597_ ( .A1(_06304_ ), .A2(_06308_ ), .ZN(_06309_ ) );
MUX2_X1 _13598_ ( .A(_06300_ ), .B(_06309_ ), .S(_05804_ ), .Z(_06310_ ) );
OAI21_X1 _13599_ ( .A(_06294_ ), .B1(_06310_ ), .B2(_06063_ ), .ZN(_06311_ ) );
NAND2_X1 _13600_ ( .A1(_06311_ ), .A2(_06066_ ), .ZN(_06312_ ) );
BUF_X4 _13601_ ( .A(_05572_ ), .Z(_06313_ ) );
BUF_X4 _13602_ ( .A(_05630_ ), .Z(_06314_ ) );
OAI211_X1 _13603_ ( .A(_06313_ ), .B(_06314_ ), .C1(_04742_ ), .C2(_04741_ ), .ZN(_06315_ ) );
BUF_X4 _13604_ ( .A(_05890_ ), .Z(_06316_ ) );
AOI21_X1 _13605_ ( .A(_04743_ ), .B1(_06315_ ), .B2(_06316_ ), .ZN(_06317_ ) );
AOI21_X1 _13606_ ( .A(_06317_ ), .B1(_04744_ ), .B2(_06186_ ), .ZN(_06318_ ) );
AND3_X1 _13607_ ( .A1(_06241_ ), .A2(_06240_ ), .A3(_05695_ ), .ZN(_06319_ ) );
OR3_X1 _13608_ ( .A1(_06319_ ), .A2(_05640_ ), .A3(_06242_ ), .ZN(_06320_ ) );
AND4_X1 _13609_ ( .A1(_06291_ ), .A2(_06312_ ), .A3(_06318_ ), .A4(_06320_ ), .ZN(_06321_ ) );
AOI21_X1 _13610_ ( .A(_05849_ ), .B1(_06280_ ), .B2(_06321_ ), .ZN(_06322_ ) );
NAND2_X1 _13611_ ( .A1(_05161_ ), .A2(_05039_ ), .ZN(_06323_ ) );
AOI22_X1 _13612_ ( .A1(_06007_ ), .A2(\EXU.ls_rdata_i [18] ), .B1(_06009_ ), .B2(\EXU.imm_i [18] ), .ZN(_06324_ ) );
OAI211_X1 _13613_ ( .A(_06323_ ), .B(_06324_ ), .C1(_06011_ ), .C2(_06274_ ), .ZN(_06325_ ) );
OR2_X1 _13614_ ( .A1(_06322_ ), .A2(_06325_ ), .ZN(_06326_ ) );
MUX2_X1 _13615_ ( .A(_06279_ ), .B(_06326_ ), .S(_05822_ ), .Z(_06327_ ) );
NAND2_X1 _13616_ ( .A1(_06327_ ), .A2(_05825_ ), .ZN(_06328_ ) );
NAND3_X1 _13617_ ( .A1(_04377_ ), .A2(_05977_ ), .A3(_06279_ ), .ZN(_06329_ ) );
AOI21_X1 _13618_ ( .A(_05515_ ), .B1(_06328_ ), .B2(_06329_ ), .ZN(_06330_ ) );
MUX2_X1 _13619_ ( .A(\EXU.xrd_o [18] ), .B(_06330_ ), .S(_04400_ ), .Z(_00246_ ) );
AND3_X1 _13620_ ( .A1(_04352_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_14_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05984_ ), .ZN(_06331_ ) );
OAI221_X1 _13621_ ( .A(_05829_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_14_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05981_ ), .C1(_05983_ ), .C2(_06331_ ), .ZN(_06332_ ) );
NAND4_X1 _13622_ ( .A1(_05987_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_14_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_05989_ ), .ZN(_06333_ ) );
NAND2_X1 _13623_ ( .A1(_06332_ ), .A2(_06333_ ), .ZN(_06334_ ) );
MUX2_X1 _13624_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_14_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ), .B(_06334_ ), .S(_05993_ ), .Z(_06335_ ) );
NAND4_X1 _13625_ ( .A1(_04756_ ), .A2(fanout_net_6 ), .A3(fanout_net_5 ), .A4(fanout_net_10 ), .ZN(_06336_ ) );
AOI22_X1 _13626_ ( .A1(_06335_ ), .A2(_04756_ ), .B1(_05996_ ), .B2(_06336_ ), .ZN(_06337_ ) );
NAND3_X1 _13627_ ( .A1(_05045_ ), .A2(\EXU.pc_i [17] ), .A3(_05999_ ), .ZN(_06338_ ) );
OAI21_X1 _13628_ ( .A(_06338_ ), .B1(_04756_ ), .B2(_06003_ ), .ZN(_06339_ ) );
OAI211_X1 _13629_ ( .A(_04371_ ), .B(_04374_ ), .C1(_06337_ ), .C2(_06339_ ), .ZN(_06340_ ) );
AOI22_X1 _13630_ ( .A1(_06007_ ), .A2(\EXU.ls_rdata_i [17] ), .B1(_06009_ ), .B2(\EXU.imm_i [17] ), .ZN(_06341_ ) );
OAI21_X1 _13631_ ( .A(_06341_ ), .B1(_06335_ ), .B2(_06012_ ), .ZN(_06342_ ) );
NAND2_X1 _13632_ ( .A1(_05178_ ), .A2(_06015_ ), .ZN(_06343_ ) );
NAND2_X1 _13633_ ( .A1(_06219_ ), .A2(_06144_ ), .ZN(_06344_ ) );
NAND3_X1 _13634_ ( .A1(_06176_ ), .A2(_05521_ ), .A3(_05878_ ), .ZN(_06345_ ) );
AOI21_X1 _13635_ ( .A(_06030_ ), .B1(_06344_ ), .B2(_06345_ ), .ZN(_06346_ ) );
AOI21_X1 _13636_ ( .A(_06096_ ), .B1(_06037_ ), .B2(_06041_ ), .ZN(_06347_ ) );
OR3_X1 _13637_ ( .A1(_06346_ ), .A2(_05804_ ), .A3(_06347_ ), .ZN(_06348_ ) );
OR3_X1 _13638_ ( .A1(_06227_ ), .A2(_06049_ ), .A3(_06228_ ), .ZN(_06349_ ) );
OR3_X1 _13639_ ( .A1(_06033_ ), .A2(_04742_ ), .A3(_06035_ ), .ZN(_06350_ ) );
OAI21_X1 _13640_ ( .A(\EXU.r1_i [17] ), .B1(_06046_ ), .B2(_06050_ ), .ZN(_06351_ ) );
NAND2_X1 _13641_ ( .A1(_06350_ ), .A2(_06351_ ), .ZN(_06352_ ) );
NAND2_X1 _13642_ ( .A1(_06352_ ), .A2(_06144_ ), .ZN(_06353_ ) );
NAND2_X1 _13643_ ( .A1(_06349_ ), .A2(_06353_ ), .ZN(_06354_ ) );
NAND2_X1 _13644_ ( .A1(_06354_ ), .A2(_05881_ ), .ZN(_06355_ ) );
BUF_X2 _13645_ ( .A(_05747_ ), .Z(_06356_ ) );
BUF_X2 _13646_ ( .A(_05924_ ), .Z(_06357_ ) );
NAND3_X1 _13647_ ( .A1(_06045_ ), .A2(_06357_ ), .A3(_06052_ ), .ZN(_06358_ ) );
NAND3_X1 _13648_ ( .A1(_06355_ ), .A2(_06356_ ), .A3(_06358_ ), .ZN(_06359_ ) );
AND2_X2 _13649_ ( .A1(_06348_ ), .A2(_06359_ ), .ZN(_06360_ ) );
BUF_X4 _13650_ ( .A(_05769_ ), .Z(_06361_ ) );
NAND2_X1 _13651_ ( .A1(_06360_ ), .A2(_06361_ ), .ZN(_06362_ ) );
NOR3_X1 _13652_ ( .A1(_05863_ ), .A2(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ), .A3(_05859_ ), .ZN(_06363_ ) );
AND2_X1 _13653_ ( .A1(_06363_ ), .A2(_06027_ ), .ZN(_06364_ ) );
OAI211_X1 _13654_ ( .A(_05871_ ), .B(_05872_ ), .C1(_06364_ ), .C2(_05856_ ), .ZN(_06365_ ) );
AOI21_X1 _13655_ ( .A(_05852_ ), .B1(_06362_ ), .B2(_06365_ ), .ZN(_06366_ ) );
AOI21_X1 _13656_ ( .A(_05692_ ), .B1(_05682_ ), .B2(_04705_ ), .ZN(_06367_ ) );
XNOR2_X1 _13657_ ( .A(_06367_ ), .B(_04704_ ), .ZN(_06368_ ) );
AND2_X1 _13658_ ( .A1(_06368_ ), .A2(_06023_ ), .ZN(_06369_ ) );
NAND3_X1 _13659_ ( .A1(_04757_ ), .A2(\EXU.r1_i [17] ), .A3(_04758_ ), .ZN(_06370_ ) );
AOI21_X1 _13660_ ( .A(_05555_ ), .B1(_05573_ ), .B2(_06370_ ), .ZN(_06371_ ) );
AND2_X1 _13661_ ( .A1(_04759_ ), .A2(_04756_ ), .ZN(_06372_ ) );
OR3_X1 _13662_ ( .A1(_06371_ ), .A2(_06372_ ), .A3(_05892_ ), .ZN(_06373_ ) );
NAND4_X1 _13663_ ( .A1(_06186_ ), .A2(_04755_ ), .A3(_04757_ ), .A4(_04758_ ), .ZN(_06374_ ) );
NAND2_X1 _13664_ ( .A1(_06373_ ), .A2(_06374_ ), .ZN(_06375_ ) );
NAND3_X1 _13665_ ( .A1(_06082_ ), .A2(_05606_ ), .A3(_06084_ ), .ZN(_06376_ ) );
NAND3_X1 _13666_ ( .A1(_06092_ ), .A2(_04996_ ), .A3(_06094_ ), .ZN(_06377_ ) );
AND3_X1 _13667_ ( .A1(_06376_ ), .A2(_06377_ ), .A3(_06060_ ), .ZN(_06378_ ) );
NAND3_X1 _13668_ ( .A1(_06086_ ), .A2(_05755_ ), .A3(_06087_ ), .ZN(_06379_ ) );
NAND3_X1 _13669_ ( .A1(_06076_ ), .A2(_05802_ ), .A3(_06078_ ), .ZN(_06380_ ) );
AOI21_X1 _13670_ ( .A(_06099_ ), .B1(_06379_ ), .B2(_06380_ ), .ZN(_06381_ ) );
OAI21_X1 _13671_ ( .A(_05769_ ), .B1(_06378_ ), .B2(_06381_ ), .ZN(_06382_ ) );
BUF_X2 _13672_ ( .A(_06039_ ), .Z(_06383_ ) );
NOR3_X1 _13673_ ( .A1(_05763_ ), .A2(_06357_ ), .A3(_06383_ ), .ZN(_06384_ ) );
NAND2_X1 _13674_ ( .A1(_06384_ ), .A2(_06356_ ), .ZN(_06385_ ) );
AOI21_X1 _13675_ ( .A(_05767_ ), .B1(_06385_ ), .B2(_06063_ ), .ZN(_06386_ ) );
AND2_X1 _13676_ ( .A1(_06382_ ), .A2(_06386_ ), .ZN(_06387_ ) );
NOR4_X1 _13677_ ( .A1(_06366_ ), .A2(_06369_ ), .A3(_06375_ ), .A4(_06387_ ), .ZN(_06388_ ) );
AOI21_X1 _13678_ ( .A(_06014_ ), .B1(_06343_ ), .B2(_06388_ ), .ZN(_06389_ ) );
AOI211_X1 _13679_ ( .A(_06342_ ), .B(_06389_ ), .C1(_05211_ ), .C2(_05172_ ), .ZN(_06390_ ) );
OAI21_X1 _13680_ ( .A(_06340_ ), .B1(_06390_ ), .B2(_06106_ ), .ZN(_06391_ ) );
NAND2_X1 _13681_ ( .A1(_06391_ ), .A2(_05825_ ), .ZN(_06392_ ) );
OAI211_X1 _13682_ ( .A(_06109_ ), .B(_05290_ ), .C1(_06337_ ), .C2(_06339_ ), .ZN(_06393_ ) );
AOI21_X1 _13683_ ( .A(_05515_ ), .B1(_06392_ ), .B2(_06393_ ), .ZN(_06394_ ) );
BUF_X4 _13684_ ( .A(_04399_ ), .Z(_06395_ ) );
MUX2_X1 _13685_ ( .A(\EXU.xrd_o [17] ), .B(_06394_ ), .S(_06395_ ), .Z(_00247_ ) );
AND3_X1 _13686_ ( .A1(_04352_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_15_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05984_ ), .ZN(_06396_ ) );
OAI221_X1 _13687_ ( .A(_05829_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_15_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05981_ ), .C1(_05983_ ), .C2(_06396_ ), .ZN(_06397_ ) );
NAND4_X1 _13688_ ( .A1(_05987_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_15_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_05988_ ), .ZN(_06398_ ) );
NAND2_X1 _13689_ ( .A1(_06397_ ), .A2(_06398_ ), .ZN(_06399_ ) );
MUX2_X1 _13690_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_15_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ), .B(_06399_ ), .S(_05993_ ), .Z(_06400_ ) );
NAND4_X1 _13691_ ( .A1(_04764_ ), .A2(fanout_net_6 ), .A3(fanout_net_5 ), .A4(fanout_net_10 ), .ZN(_06401_ ) );
AOI22_X1 _13692_ ( .A1(_06400_ ), .A2(_04764_ ), .B1(_05996_ ), .B2(_06401_ ), .ZN(_06402_ ) );
NAND3_X1 _13693_ ( .A1(_05045_ ), .A2(\EXU.pc_i [16] ), .A3(_05999_ ), .ZN(_06403_ ) );
OAI21_X1 _13694_ ( .A(_06403_ ), .B1(_04764_ ), .B2(_06003_ ), .ZN(_06404_ ) );
OAI211_X1 _13695_ ( .A(_04371_ ), .B(_04374_ ), .C1(_06402_ ), .C2(_06404_ ), .ZN(_06405_ ) );
AOI22_X1 _13696_ ( .A1(_06007_ ), .A2(\EXU.ls_rdata_i [16] ), .B1(_06009_ ), .B2(\EXU.imm_i [16] ), .ZN(_06406_ ) );
OAI21_X1 _13697_ ( .A(_06406_ ), .B1(_06400_ ), .B2(_06012_ ), .ZN(_06407_ ) );
NAND2_X1 _13698_ ( .A1(_05187_ ), .A2(_06015_ ), .ZN(_06408_ ) );
NAND2_X1 _13699_ ( .A1(_06153_ ), .A2(_06152_ ), .ZN(_06409_ ) );
NOR2_X1 _13700_ ( .A1(_06409_ ), .A2(_05866_ ), .ZN(_06410_ ) );
OAI211_X1 _13701_ ( .A(_05871_ ), .B(_05872_ ), .C1(_05856_ ), .C2(_06410_ ), .ZN(_06411_ ) );
OR3_X4 _13702_ ( .A1(_06296_ ), .A2(_05878_ ), .A3(_06297_ ), .ZN(_06412_ ) );
MUX2_X1 _13703_ ( .A(\EXU.r1_i [30] ), .B(\EXU.r1_i [31] ), .S(_06040_ ), .Z(_06413_ ) );
BUF_X2 _13704_ ( .A(_06049_ ), .Z(_06414_ ) );
OAI211_X1 _13705_ ( .A(_06412_ ), .B(_06357_ ), .C1(_06413_ ), .C2(_06414_ ), .ZN(_06415_ ) );
NAND3_X1 _13706_ ( .A1(_06167_ ), .A2(_05881_ ), .A3(_06170_ ), .ZN(_06416_ ) );
NAND3_X1 _13707_ ( .A1(_06415_ ), .A2(_06416_ ), .A3(_06099_ ), .ZN(_06417_ ) );
AND3_X1 _13708_ ( .A1(_06174_ ), .A2(_06077_ ), .A3(_06177_ ), .ZN(_06418_ ) );
OR3_X1 _13709_ ( .A1(_05597_ ), .A2(_04756_ ), .A3(_05598_ ), .ZN(_06419_ ) );
OAI211_X1 _13710_ ( .A(_06419_ ), .B(_04901_ ), .C1(_04764_ ), .C2(_05600_ ), .ZN(_06420_ ) );
OR3_X1 _13711_ ( .A1(_05597_ ), .A2(_04750_ ), .A3(_05598_ ), .ZN(_06421_ ) );
OAI211_X1 _13712_ ( .A(_06421_ ), .B(_05602_ ), .C1(_04742_ ), .C2(_05600_ ), .ZN(_06422_ ) );
AOI21_X1 _13713_ ( .A(_06357_ ), .B1(_06420_ ), .B2(_06422_ ), .ZN(_06423_ ) );
NOR2_X1 _13714_ ( .A1(_06418_ ), .A2(_06423_ ), .ZN(_06424_ ) );
OAI21_X1 _13715_ ( .A(_06417_ ), .B1(_06424_ ), .B2(_06081_ ), .ZN(_06425_ ) );
OAI21_X1 _13716_ ( .A(_06411_ ), .B1(_06425_ ), .B2(_06063_ ), .ZN(_06426_ ) );
AND2_X1 _13717_ ( .A1(_06426_ ), .A2(_06066_ ), .ZN(_06427_ ) );
XNOR2_X1 _13718_ ( .A(_05682_ ), .B(_04705_ ), .ZN(_06428_ ) );
NOR2_X1 _13719_ ( .A1(_05641_ ), .A2(_06428_ ), .ZN(_06429_ ) );
OAI211_X1 _13720_ ( .A(_06313_ ), .B(_06314_ ), .C1(_04764_ ), .C2(_04763_ ), .ZN(_06430_ ) );
AOI21_X1 _13721_ ( .A(_04765_ ), .B1(_06430_ ), .B2(_06316_ ), .ZN(_06431_ ) );
AND2_X1 _13722_ ( .A1(_04766_ ), .A2(_05892_ ), .ZN(_06432_ ) );
OR2_X1 _13723_ ( .A1(_06431_ ), .A2(_06432_ ), .ZN(_06433_ ) );
AND3_X1 _13724_ ( .A1(_04998_ ), .A2(_06030_ ), .A3(_06414_ ), .ZN(_06434_ ) );
AND2_X1 _13725_ ( .A1(_06434_ ), .A2(_06356_ ), .ZN(_06435_ ) );
OAI21_X1 _13726_ ( .A(_05565_ ), .B1(_06435_ ), .B2(_05769_ ), .ZN(_06436_ ) );
OAI211_X1 _13727_ ( .A(_06139_ ), .B(_06096_ ), .C1(_06140_ ), .C2(_06144_ ), .ZN(_06437_ ) );
OAI211_X1 _13728_ ( .A(_06146_ ), .B(_05934_ ), .C1(_05901_ ), .C2(_06144_ ), .ZN(_06438_ ) );
NAND2_X1 _13729_ ( .A1(_06437_ ), .A2(_06438_ ), .ZN(_06439_ ) );
NAND2_X1 _13730_ ( .A1(_06132_ ), .A2(_06077_ ), .ZN(_06440_ ) );
OAI211_X1 _13731_ ( .A(_06137_ ), .B(_05934_ ), .C1(_05909_ ), .C2(_05878_ ), .ZN(_06441_ ) );
NAND2_X1 _13732_ ( .A1(_06440_ ), .A2(_06441_ ), .ZN(_06442_ ) );
MUX2_X1 _13733_ ( .A(_06439_ ), .B(_06442_ ), .S(_06081_ ), .Z(_06443_ ) );
AOI21_X1 _13734_ ( .A(_06436_ ), .B1(_06443_ ), .B2(_06091_ ), .ZN(_06444_ ) );
NOR4_X2 _13735_ ( .A1(_06427_ ), .A2(_06429_ ), .A3(_06433_ ), .A4(_06444_ ), .ZN(_06445_ ) );
AOI21_X1 _13736_ ( .A(_06014_ ), .B1(_06408_ ), .B2(_06445_ ), .ZN(_06446_ ) );
AOI211_X1 _13737_ ( .A(_06407_ ), .B(_06446_ ), .C1(_05211_ ), .C2(_05183_ ), .ZN(_06447_ ) );
OAI21_X1 _13738_ ( .A(_06405_ ), .B1(_06447_ ), .B2(_06106_ ), .ZN(_06448_ ) );
NAND2_X1 _13739_ ( .A1(_06448_ ), .A2(_05825_ ), .ZN(_06449_ ) );
OAI211_X1 _13740_ ( .A(_06109_ ), .B(_05290_ ), .C1(_06402_ ), .C2(_06404_ ), .ZN(_06450_ ) );
AOI21_X1 _13741_ ( .A(_05515_ ), .B1(_06449_ ), .B2(_06450_ ), .ZN(_06451_ ) );
MUX2_X1 _13742_ ( .A(\EXU.xrd_o [16] ), .B(_06451_ ), .S(_06395_ ), .Z(_00248_ ) );
NAND3_X1 _13743_ ( .A1(_06203_ ), .A2(\EXU.mcause_i [15] ), .A3(_05836_ ), .ZN(_06452_ ) );
NAND3_X1 _13744_ ( .A1(_06118_ ), .A2(\EXU.mstatus_i [15] ), .A3(_05988_ ), .ZN(_06453_ ) );
NAND3_X1 _13745_ ( .A1(_06118_ ), .A2(\EXU.mtvec_i [15] ), .A3(_06208_ ), .ZN(_06454_ ) );
NAND4_X1 _13746_ ( .A1(_06202_ ), .A2(_06452_ ), .A3(_06453_ ), .A4(_06454_ ), .ZN(_06455_ ) );
OAI21_X1 _13747_ ( .A(_06455_ ), .B1(\EXU.mepc_i [15] ), .B2(_05992_ ), .ZN(_06456_ ) );
NAND4_X1 _13748_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_16_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_06457_ ) );
AOI22_X1 _13749_ ( .A1(_06456_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_16_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_05995_ ), .B2(_06457_ ), .ZN(_06458_ ) );
NAND3_X1 _13750_ ( .A1(_06123_ ), .A2(\EXU.pc_i [15] ), .A3(_04348_ ), .ZN(_06459_ ) );
OAI21_X1 _13751_ ( .A(_06459_ ), .B1(_05017_ ), .B2(_06002_ ), .ZN(_06460_ ) );
OR2_X1 _13752_ ( .A1(_06458_ ), .A2(_06460_ ), .ZN(_06461_ ) );
NAND2_X1 _13753_ ( .A1(_05198_ ), .A2(_05850_ ), .ZN(_06462_ ) );
OAI21_X1 _13754_ ( .A(_06065_ ), .B1(_05608_ ), .B2(_05769_ ), .ZN(_06463_ ) );
NAND3_X1 _13755_ ( .A1(_06220_ ), .A2(_06357_ ), .A3(_06221_ ), .ZN(_06464_ ) );
NAND3_X1 _13756_ ( .A1(_06224_ ), .A2(_06225_ ), .A3(_06030_ ), .ZN(_06465_ ) );
NAND2_X1 _13757_ ( .A1(_06464_ ), .A2(_06465_ ), .ZN(_06466_ ) );
NAND2_X1 _13758_ ( .A1(_06466_ ), .A2(_06081_ ), .ZN(_06467_ ) );
NAND3_X1 _13759_ ( .A1(_06229_ ), .A2(_06096_ ), .A3(_06231_ ), .ZN(_06468_ ) );
NOR2_X1 _13760_ ( .A1(_05601_ ), .A2(\EXU.r1_i [15] ), .ZN(_06469_ ) );
NOR3_X1 _13761_ ( .A1(_06160_ ), .A2(\EXU.r1_i [16] ), .A3(_06047_ ), .ZN(_06470_ ) );
OR3_X1 _13762_ ( .A1(_06469_ ), .A2(_05604_ ), .A3(_06470_ ), .ZN(_06471_ ) );
NAND2_X1 _13763_ ( .A1(_06352_ ), .A2(_06039_ ), .ZN(_06472_ ) );
NAND3_X1 _13764_ ( .A1(_06471_ ), .A2(_05607_ ), .A3(_06472_ ), .ZN(_06473_ ) );
AND2_X1 _13765_ ( .A1(_06468_ ), .A2(_06473_ ), .ZN(_06474_ ) );
OAI21_X1 _13766_ ( .A(_06467_ ), .B1(_06100_ ), .B2(_06474_ ), .ZN(_06475_ ) );
AOI21_X1 _13767_ ( .A(_06463_ ), .B1(_06475_ ), .B2(_06091_ ), .ZN(_06476_ ) );
NOR3_X1 _13768_ ( .A1(_05589_ ), .A2(_04725_ ), .A3(_05582_ ), .ZN(_06477_ ) );
NAND3_X1 _13769_ ( .A1(_05622_ ), .A2(_05625_ ), .A3(_06477_ ), .ZN(_06478_ ) );
INV_X1 _13770_ ( .A(_04681_ ), .ZN(_06479_ ) );
NOR2_X1 _13771_ ( .A1(_05653_ ), .A2(_05661_ ), .ZN(_06480_ ) );
INV_X1 _13772_ ( .A(_06480_ ), .ZN(_06481_ ) );
AND2_X1 _13773_ ( .A1(_06481_ ), .A2(_04700_ ), .ZN(_06482_ ) );
NOR2_X1 _13774_ ( .A1(_06482_ ), .A2(_05680_ ), .ZN(_06483_ ) );
NOR3_X1 _13775_ ( .A1(_06483_ ), .A2(_04684_ ), .A3(_04686_ ), .ZN(_06484_ ) );
INV_X1 _13776_ ( .A(_06484_ ), .ZN(_06485_ ) );
AOI21_X1 _13777_ ( .A(_06479_ ), .B1(_06485_ ), .B2(_05668_ ), .ZN(_06486_ ) );
AOI21_X1 _13778_ ( .A(_06486_ ), .B1(\EXU.r1_i [14] ), .B2(_05663_ ), .ZN(_06487_ ) );
XNOR2_X1 _13779_ ( .A(_06487_ ), .B(_04680_ ), .ZN(_06488_ ) );
NAND2_X1 _13780_ ( .A1(_06488_ ), .A2(_06023_ ), .ZN(_06489_ ) );
NAND3_X1 _13781_ ( .A1(_04853_ ), .A2(\EXU.r1_i [15] ), .A3(_04855_ ), .ZN(_06490_ ) );
AND3_X1 _13782_ ( .A1(_05572_ ), .A2(_05630_ ), .A3(_06490_ ), .ZN(_06491_ ) );
OAI22_X1 _13783_ ( .A1(_06491_ ), .A2(_05555_ ), .B1(\EXU.r1_i [15] ), .B2(_04858_ ), .ZN(_06492_ ) );
MUX2_X1 _13784_ ( .A(_04856_ ), .B(_06492_ ), .S(_05635_ ), .Z(_06493_ ) );
AOI22_X1 _13785_ ( .A1(_04950_ ), .A2(_04952_ ), .B1(_04437_ ), .B2(_04730_ ), .ZN(_06494_ ) );
AND2_X2 _13786_ ( .A1(_06494_ ), .A2(_05565_ ), .ZN(_06495_ ) );
NAND3_X1 _13787_ ( .A1(_05748_ ), .A2(_05765_ ), .A3(_06495_ ), .ZN(_06496_ ) );
NAND4_X1 _13788_ ( .A1(_06478_ ), .A2(_06489_ ), .A3(_06493_ ), .A4(_06496_ ), .ZN(_06497_ ) );
NOR2_X1 _13789_ ( .A1(_06476_ ), .A2(_06497_ ), .ZN(_06498_ ) );
AOI21_X1 _13790_ ( .A(_05849_ ), .B1(_06462_ ), .B2(_06498_ ), .ZN(_06499_ ) );
CLKBUF_X2 _13791_ ( .A(_05038_ ), .Z(_06500_ ) );
AND2_X1 _13792_ ( .A1(_05203_ ), .A2(_06500_ ), .ZN(_06501_ ) );
AOI22_X1 _13793_ ( .A1(_06006_ ), .A2(\EXU.ls_rdata_i [15] ), .B1(_06008_ ), .B2(\EXU.imm_i [15] ), .ZN(_06502_ ) );
OAI21_X1 _13794_ ( .A(_06502_ ), .B1(_06456_ ), .B2(_05814_ ), .ZN(_06503_ ) );
OR3_X1 _13795_ ( .A1(_06499_ ), .A2(_06501_ ), .A3(_06503_ ), .ZN(_06504_ ) );
MUX2_X1 _13796_ ( .A(_06461_ ), .B(_06504_ ), .S(_05822_ ), .Z(_06505_ ) );
NAND2_X1 _13797_ ( .A1(_06505_ ), .A2(_05825_ ), .ZN(_06506_ ) );
NAND3_X1 _13798_ ( .A1(_04377_ ), .A2(_05977_ ), .A3(_06461_ ), .ZN(_06507_ ) );
AOI21_X1 _13799_ ( .A(_05515_ ), .B1(_06506_ ), .B2(_06507_ ), .ZN(_06508_ ) );
MUX2_X1 _13800_ ( .A(\EXU.xrd_o [15] ), .B(_06508_ ), .S(_06395_ ), .Z(_00249_ ) );
AND3_X1 _13801_ ( .A1(_06118_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_17_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05831_ ), .ZN(_06509_ ) );
OAI221_X1 _13802_ ( .A(_05829_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_17_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05981_ ), .C1(_05983_ ), .C2(_06509_ ), .ZN(_06510_ ) );
NAND4_X1 _13803_ ( .A1(_05987_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_17_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_05989_ ), .ZN(_06511_ ) );
NAND2_X1 _13804_ ( .A1(_06510_ ), .A2(_06511_ ), .ZN(_06512_ ) );
MUX2_X1 _13805_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_17_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ), .B(_06512_ ), .S(_05993_ ), .Z(_06513_ ) );
NAND4_X1 _13806_ ( .A1(_04864_ ), .A2(fanout_net_6 ), .A3(fanout_net_5 ), .A4(fanout_net_10 ), .ZN(_06514_ ) );
AOI22_X1 _13807_ ( .A1(_06513_ ), .A2(_04864_ ), .B1(_05996_ ), .B2(_06514_ ), .ZN(_06515_ ) );
BUF_X2 _13808_ ( .A(_05044_ ), .Z(_06516_ ) );
NAND3_X1 _13809_ ( .A1(_06516_ ), .A2(\EXU.pc_i [14] ), .A3(_05999_ ), .ZN(_06517_ ) );
OAI21_X1 _13810_ ( .A(_06517_ ), .B1(_04864_ ), .B2(_06003_ ), .ZN(_06518_ ) );
OAI211_X1 _13811_ ( .A(_04371_ ), .B(_04374_ ), .C1(_06515_ ), .C2(_06518_ ), .ZN(_06519_ ) );
NAND2_X1 _13812_ ( .A1(_05209_ ), .A2(_06015_ ), .ZN(_06520_ ) );
NAND3_X1 _13813_ ( .A1(_06301_ ), .A2(_06303_ ), .A3(_06289_ ), .ZN(_06521_ ) );
OR3_X1 _13814_ ( .A1(_05597_ ), .A2(_05017_ ), .A3(_05598_ ), .ZN(_06522_ ) );
OAI21_X2 _13815_ ( .A(\EXU.r1_i [14] ), .B1(_06032_ ), .B2(_06034_ ), .ZN(_06523_ ) );
NAND2_X1 _13816_ ( .A1(_06522_ ), .A2(_06523_ ), .ZN(_06524_ ) );
NAND2_X1 _13817_ ( .A1(_06524_ ), .A2(_06414_ ), .ZN(_06525_ ) );
BUF_X4 _13818_ ( .A(_06030_ ), .Z(_06526_ ) );
BUF_X2 _13819_ ( .A(_06160_ ), .Z(_06527_ ) );
BUF_X2 _13820_ ( .A(_06047_ ), .Z(_06528_ ) );
OR3_X1 _13821_ ( .A1(_06527_ ), .A2(\EXU.r1_i [17] ), .A3(_06528_ ), .ZN(_06529_ ) );
OAI211_X1 _13822_ ( .A(_06529_ ), .B(_06383_ ), .C1(\EXU.r1_i [16] ), .C2(_06040_ ), .ZN(_06530_ ) );
NAND3_X1 _13823_ ( .A1(_06525_ ), .A2(_06526_ ), .A3(_06530_ ), .ZN(_06531_ ) );
BUF_X4 _13824_ ( .A(_05880_ ), .Z(_06532_ ) );
NAND3_X1 _13825_ ( .A1(_06521_ ), .A2(_06531_ ), .A3(_06532_ ), .ZN(_06533_ ) );
AOI21_X1 _13826_ ( .A(_05934_ ), .B1(_06295_ ), .B2(_06298_ ), .ZN(_06534_ ) );
AOI21_X1 _13827_ ( .A(_06096_ ), .B1(_06306_ ), .B2(_06307_ ), .ZN(_06535_ ) );
NOR2_X1 _13828_ ( .A1(_06534_ ), .A2(_06535_ ), .ZN(_06536_ ) );
OAI211_X1 _13829_ ( .A(_06091_ ), .B(_06533_ ), .C1(_06536_ ), .C2(_06532_ ), .ZN(_06537_ ) );
BUF_X4 _13830_ ( .A(_06066_ ), .Z(_06538_ ) );
OAI211_X1 _13831_ ( .A(_06537_ ), .B(_06538_ ), .C1(_06361_ ), .C2(_05882_ ), .ZN(_06539_ ) );
AND3_X1 _13832_ ( .A1(_06485_ ), .A2(_06479_ ), .A3(_05668_ ), .ZN(_06540_ ) );
NOR3_X1 _13833_ ( .A1(_06540_ ), .A2(_06486_ ), .A3(_05641_ ), .ZN(_06541_ ) );
INV_X1 _13834_ ( .A(_06495_ ), .ZN(_06542_ ) );
AOI21_X1 _13835_ ( .A(_06542_ ), .B1(_05913_ ), .B2(_05926_ ), .ZN(_06543_ ) );
NAND3_X1 _13836_ ( .A1(_04860_ ), .A2(\EXU.r1_i [14] ), .A3(_04861_ ), .ZN(_06544_ ) );
NAND3_X1 _13837_ ( .A1(_06313_ ), .A2(_06314_ ), .A3(_06544_ ), .ZN(_06545_ ) );
AOI21_X1 _13838_ ( .A(_04865_ ), .B1(_06545_ ), .B2(_06316_ ), .ZN(_06546_ ) );
MUX2_X1 _13839_ ( .A(_04863_ ), .B(_06546_ ), .S(_06071_ ), .Z(_06547_ ) );
NOR3_X1 _13840_ ( .A1(_06541_ ), .A2(_06543_ ), .A3(_06547_ ), .ZN(_06548_ ) );
AND2_X1 _13841_ ( .A1(_05853_ ), .A2(_05590_ ), .ZN(_06549_ ) );
BUF_X2 _13842_ ( .A(_06549_ ), .Z(_06550_ ) );
NAND3_X1 _13843_ ( .A1(_05867_ ), .A2(_05868_ ), .A3(_06550_ ), .ZN(_06551_ ) );
AND3_X1 _13844_ ( .A1(_06539_ ), .A2(_06548_ ), .A3(_06551_ ), .ZN(_06552_ ) );
AOI21_X1 _13845_ ( .A(_06014_ ), .B1(_06520_ ), .B2(_06552_ ), .ZN(_06553_ ) );
NOR2_X1 _13846_ ( .A1(_05214_ ), .A2(_05189_ ), .ZN(_06554_ ) );
NAND3_X1 _13847_ ( .A1(_05967_ ), .A2(_05968_ ), .A3(\EXU.imm_i [14] ), .ZN(_06555_ ) );
INV_X1 _13848_ ( .A(\EXU.ls_rdata_i [14] ), .ZN(_06556_ ) );
OAI221_X1 _13849_ ( .A(_06555_ ), .B1(_06556_ ), .B2(_04414_ ), .C1(_06513_ ), .C2(_06012_ ), .ZN(_06557_ ) );
NOR3_X1 _13850_ ( .A1(_06553_ ), .A2(_06554_ ), .A3(_06557_ ), .ZN(_06558_ ) );
OAI21_X1 _13851_ ( .A(_06519_ ), .B1(_06558_ ), .B2(_06106_ ), .ZN(_06559_ ) );
NAND2_X1 _13852_ ( .A1(_06559_ ), .A2(_05825_ ), .ZN(_06560_ ) );
OAI211_X1 _13853_ ( .A(_06109_ ), .B(_05290_ ), .C1(_06515_ ), .C2(_06518_ ), .ZN(_06561_ ) );
AOI21_X1 _13854_ ( .A(_05515_ ), .B1(_06560_ ), .B2(_06561_ ), .ZN(_06562_ ) );
MUX2_X1 _13855_ ( .A(\EXU.xrd_o [14] ), .B(_06562_ ), .S(_06395_ ), .Z(_00250_ ) );
BUF_X4 _13856_ ( .A(_04395_ ), .Z(_06563_ ) );
AND3_X1 _13857_ ( .A1(_06118_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_18_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05831_ ), .ZN(_06564_ ) );
OAI221_X1 _13858_ ( .A(_05830_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_18_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05981_ ), .C1(_05983_ ), .C2(_06564_ ), .ZN(_06565_ ) );
NAND4_X1 _13859_ ( .A1(_05987_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_18_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_05989_ ), .ZN(_06566_ ) );
NAND2_X1 _13860_ ( .A1(_06565_ ), .A2(_06566_ ), .ZN(_06567_ ) );
MUX2_X1 _13861_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_18_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ), .B(_06567_ ), .S(_05993_ ), .Z(_06568_ ) );
NAND4_X1 _13862_ ( .A1(_05020_ ), .A2(fanout_net_6 ), .A3(fanout_net_5 ), .A4(fanout_net_10 ), .ZN(_06569_ ) );
AOI22_X1 _13863_ ( .A1(_06568_ ), .A2(_05020_ ), .B1(_05996_ ), .B2(_06569_ ), .ZN(_06570_ ) );
NAND3_X1 _13864_ ( .A1(_06516_ ), .A2(\EXU.pc_i [13] ), .A3(_05999_ ), .ZN(_06571_ ) );
OAI21_X1 _13865_ ( .A(_06571_ ), .B1(_05020_ ), .B2(_06003_ ), .ZN(_06572_ ) );
OAI211_X1 _13866_ ( .A(_04371_ ), .B(_04374_ ), .C1(_06570_ ), .C2(_06572_ ), .ZN(_06573_ ) );
NAND2_X1 _13867_ ( .A1(_05228_ ), .A2(_06015_ ), .ZN(_06574_ ) );
NOR2_X1 _13868_ ( .A1(_05600_ ), .A2(\EXU.r1_i [13] ), .ZN(_06575_ ) );
NOR3_X2 _13869_ ( .A1(_06033_ ), .A2(\EXU.r1_i [14] ), .A3(_06035_ ), .ZN(_06576_ ) );
OAI21_X1 _13870_ ( .A(_06144_ ), .B1(_06575_ ), .B2(_06576_ ), .ZN(_06577_ ) );
OAI21_X1 _13871_ ( .A(_06039_ ), .B1(_06469_ ), .B2(_06470_ ), .ZN(_06578_ ) );
AND2_X1 _13872_ ( .A1(_06577_ ), .A2(_06578_ ), .ZN(_06579_ ) );
MUX2_X1 _13873_ ( .A(_06579_ ), .B(_06354_ ), .S(_06289_ ), .Z(_06580_ ) );
NAND2_X1 _13874_ ( .A1(_06580_ ), .A2(_06532_ ), .ZN(_06581_ ) );
OAI21_X1 _13875_ ( .A(_06100_ ), .B1(_06042_ ), .B2(_06053_ ), .ZN(_06582_ ) );
AND3_X1 _13876_ ( .A1(_06581_ ), .A2(_06091_ ), .A3(_06582_ ), .ZN(_06583_ ) );
AND3_X1 _13877_ ( .A1(_06059_ ), .A2(_05747_ ), .A3(_06030_ ), .ZN(_06584_ ) );
OAI21_X1 _13878_ ( .A(_06538_ ), .B1(_06584_ ), .B2(_06361_ ), .ZN(_06585_ ) );
NOR2_X1 _13879_ ( .A1(_06583_ ), .A2(_06585_ ), .ZN(_06586_ ) );
NOR2_X1 _13880_ ( .A1(_06483_ ), .A2(_04686_ ), .ZN(_06587_ ) );
OR3_X1 _13881_ ( .A1(_06587_ ), .A2(_04684_ ), .A3(_05665_ ), .ZN(_06588_ ) );
OAI21_X1 _13882_ ( .A(_04684_ ), .B1(_06587_ ), .B2(_05665_ ), .ZN(_06589_ ) );
AOI21_X1 _13883_ ( .A(_05641_ ), .B1(_06588_ ), .B2(_06589_ ), .ZN(_06590_ ) );
OAI21_X1 _13884_ ( .A(_06186_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_04869_ ), .ZN(_06591_ ) );
NAND3_X1 _13885_ ( .A1(_04867_ ), .A2(\EXU.r1_i [13] ), .A3(_04868_ ), .ZN(_06592_ ) );
NAND3_X1 _13886_ ( .A1(_06313_ ), .A2(_06314_ ), .A3(_06592_ ), .ZN(_06593_ ) );
AOI22_X1 _13887_ ( .A1(_06593_ ), .A2(_06316_ ), .B1(_05020_ ), .B2(_04869_ ), .ZN(_06594_ ) );
OAI211_X1 _13888_ ( .A(_04427_ ), .B(_06591_ ), .C1(_06594_ ), .C2(_06186_ ), .ZN(_06595_ ) );
NOR2_X1 _13889_ ( .A1(_06089_ ), .A2(_05960_ ), .ZN(_06596_ ) );
NOR2_X1 _13890_ ( .A1(_06098_ ), .A2(_05804_ ), .ZN(_06597_ ) );
NOR2_X1 _13891_ ( .A1(_06596_ ), .A2(_06597_ ), .ZN(_06598_ ) );
OAI21_X1 _13892_ ( .A(_06595_ ), .B1(_06598_ ), .B2(_06542_ ), .ZN(_06599_ ) );
OR2_X2 _13893_ ( .A1(_06025_ ), .A2(_06026_ ), .ZN(_06600_ ) );
AND3_X1 _13894_ ( .A1(_06600_ ), .A2(_05868_ ), .A3(_06550_ ), .ZN(_06601_ ) );
NOR4_X1 _13895_ ( .A1(_06586_ ), .A2(_06590_ ), .A3(_06599_ ), .A4(_06601_ ), .ZN(_06602_ ) );
AOI21_X1 _13896_ ( .A(_06014_ ), .B1(_06574_ ), .B2(_06602_ ), .ZN(_06603_ ) );
NOR2_X1 _13897_ ( .A1(_05222_ ), .A2(_05189_ ), .ZN(_06604_ ) );
NAND3_X1 _13898_ ( .A1(_05967_ ), .A2(_05968_ ), .A3(\EXU.imm_i [13] ), .ZN(_06605_ ) );
NAND3_X1 _13899_ ( .A1(_05970_ ), .A2(\EXU.ls_rdata_i [13] ), .A3(_05971_ ), .ZN(_06606_ ) );
OAI211_X1 _13900_ ( .A(_06605_ ), .B(_06606_ ), .C1(_06568_ ), .C2(_06012_ ), .ZN(_06607_ ) );
NOR3_X1 _13901_ ( .A1(_06603_ ), .A2(_06604_ ), .A3(_06607_ ), .ZN(_06608_ ) );
OAI21_X1 _13902_ ( .A(_06573_ ), .B1(_06608_ ), .B2(_06106_ ), .ZN(_06609_ ) );
BUF_X4 _13903_ ( .A(_05824_ ), .Z(_06610_ ) );
NAND2_X1 _13904_ ( .A1(_06609_ ), .A2(_06610_ ), .ZN(_06611_ ) );
OAI211_X1 _13905_ ( .A(_06109_ ), .B(_05290_ ), .C1(_06570_ ), .C2(_06572_ ), .ZN(_06612_ ) );
AOI21_X1 _13906_ ( .A(_06563_ ), .B1(_06611_ ), .B2(_06612_ ), .ZN(_06613_ ) );
MUX2_X1 _13907_ ( .A(\EXU.xrd_o [13] ), .B(_06613_ ), .S(_06395_ ), .Z(_00251_ ) );
NAND4_X1 _13908_ ( .A1(_05831_ ), .A2(_05832_ ), .A3(\EXU.mtvec_i [12] ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_06614_ ) );
AOI22_X1 _13909_ ( .A1(_06614_ ), .A2(_05835_ ), .B1(_05836_ ), .B2(_06203_ ), .ZN(_06615_ ) );
AND3_X1 _13910_ ( .A1(_06203_ ), .A2(\EXU.mcause_i [12] ), .A3(_05836_ ), .ZN(_06616_ ) );
OAI21_X1 _13911_ ( .A(_05830_ ), .B1(_06615_ ), .B2(_06616_ ), .ZN(_06617_ ) );
NAND3_X1 _13912_ ( .A1(_06204_ ), .A2(_06208_ ), .A3(\EXU.mepc_i [12] ), .ZN(_06618_ ) );
NAND3_X1 _13913_ ( .A1(_06206_ ), .A2(\EXU.mstatus_i [12] ), .A3(_05989_ ), .ZN(_06619_ ) );
AND3_X1 _13914_ ( .A1(_06617_ ), .A2(_06618_ ), .A3(_06619_ ), .ZN(_06620_ ) );
NAND4_X1 _13915_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_19_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_06621_ ) );
AOI22_X1 _13916_ ( .A1(_06620_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_19_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_05996_ ), .B2(_06621_ ), .ZN(_06622_ ) );
NAND3_X1 _13917_ ( .A1(_06516_ ), .A2(\EXU.pc_i [12] ), .A3(_05999_ ), .ZN(_06623_ ) );
OAI21_X1 _13918_ ( .A(_06623_ ), .B1(_04877_ ), .B2(_06003_ ), .ZN(_06624_ ) );
OAI211_X1 _13919_ ( .A(_04374_ ), .B(_04370_ ), .C1(_06622_ ), .C2(_06624_ ), .ZN(_06625_ ) );
INV_X1 _13920_ ( .A(_05849_ ), .ZN(_06626_ ) );
AOI211_X1 _13921_ ( .A(_04685_ ), .B(_05680_ ), .C1(_06481_ ), .C2(_04700_ ), .ZN(_06627_ ) );
NOR3_X1 _13922_ ( .A1(_06587_ ), .A2(_05641_ ), .A3(_06627_ ), .ZN(_06628_ ) );
AND2_X1 _13923_ ( .A1(_06420_ ), .A2(_06422_ ), .ZN(_06629_ ) );
NOR2_X4 _13924_ ( .A1(_05600_ ), .A2(\EXU.r1_i [12] ), .ZN(_06630_ ) );
NOR3_X1 _13925_ ( .A1(_05597_ ), .A2(\EXU.r1_i [13] ), .A3(_05598_ ), .ZN(_06631_ ) );
OR3_X4 _13926_ ( .A1(_06630_ ), .A2(_05602_ ), .A3(_06631_ ), .ZN(_06632_ ) );
NAND2_X2 _13927_ ( .A1(_06524_ ), .A2(_05603_ ), .ZN(_06633_ ) );
NAND2_X1 _13928_ ( .A1(_06632_ ), .A2(_06633_ ), .ZN(_06634_ ) );
MUX2_X1 _13929_ ( .A(_06629_ ), .B(_06634_ ), .S(_04892_ ), .Z(_06635_ ) );
NAND2_X2 _13930_ ( .A1(_06635_ ), .A2(_04885_ ), .ZN(_06636_ ) );
NAND2_X2 _13931_ ( .A1(_06179_ ), .A2(_05757_ ), .ZN(_06637_ ) );
AOI21_X2 _13932_ ( .A(_05914_ ), .B1(_06636_ ), .B2(_06637_ ), .ZN(_06638_ ) );
NAND2_X1 _13933_ ( .A1(_06157_ ), .A2(_06163_ ), .ZN(_06639_ ) );
NOR4_X1 _13934_ ( .A1(_06639_ ), .A2(_04954_ ), .A3(_05757_ ), .A4(_06096_ ), .ZN(_06640_ ) );
NOR2_X2 _13935_ ( .A1(_06638_ ), .A2(_06640_ ), .ZN(_06641_ ) );
OAI221_X1 _13936_ ( .A(_05866_ ), .B1(_06151_ ), .B2(_05859_ ), .C1(_05863_ ), .C2(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ), .ZN(_06642_ ) );
NAND3_X1 _13937_ ( .A1(_06642_ ), .A2(_05853_ ), .A3(_05868_ ), .ZN(_06643_ ) );
AOI21_X1 _13938_ ( .A(_05591_ ), .B1(_06641_ ), .B2(_06643_ ), .ZN(_06644_ ) );
OAI211_X1 _13939_ ( .A(_05887_ ), .B(_05888_ ), .C1(_04877_ ), .C2(_04875_ ), .ZN(_06645_ ) );
AOI21_X1 _13940_ ( .A(_04878_ ), .B1(_06645_ ), .B2(_05890_ ), .ZN(_06646_ ) );
AND2_X1 _13941_ ( .A1(_04876_ ), .A2(_05892_ ), .ZN(_06647_ ) );
OR3_X2 _13942_ ( .A1(_06644_ ), .A2(_06646_ ), .A3(_06647_ ), .ZN(_06648_ ) );
INV_X1 _13943_ ( .A(_05809_ ), .ZN(_06649_ ) );
NOR3_X1 _13944_ ( .A1(_06641_ ), .A2(_04425_ ), .A3(_06649_ ), .ZN(_06650_ ) );
NOR2_X1 _13945_ ( .A1(_06133_ ), .A2(_05804_ ), .ZN(_06651_ ) );
AOI21_X1 _13946_ ( .A(_06651_ ), .B1(_05880_ ), .B2(_06142_ ), .ZN(_06652_ ) );
NOR4_X1 _13947_ ( .A1(_06652_ ), .A2(_04425_ ), .A3(_06181_ ), .A4(_05767_ ), .ZN(_06653_ ) );
OR4_X2 _13948_ ( .A1(_06628_ ), .A2(_06648_ ), .A3(_06650_ ), .A4(_06653_ ), .ZN(_06654_ ) );
AND2_X1 _13949_ ( .A1(_05236_ ), .A2(_05850_ ), .ZN(_06655_ ) );
OAI21_X2 _13950_ ( .A(_06626_ ), .B1(_06654_ ), .B2(_06655_ ), .ZN(_06656_ ) );
NAND2_X1 _13951_ ( .A1(_05232_ ), .A2(_05039_ ), .ZN(_06657_ ) );
OR2_X1 _13952_ ( .A1(_06620_ ), .A2(_06011_ ), .ZN(_06658_ ) );
AND3_X1 _13953_ ( .A1(_05970_ ), .A2(\EXU.ls_rdata_i [12] ), .A3(_05971_ ), .ZN(_06659_ ) );
AND3_X1 _13954_ ( .A1(_05967_ ), .A2(_05968_ ), .A3(\EXU.imm_i [12] ), .ZN(_06660_ ) );
NOR2_X1 _13955_ ( .A1(_06659_ ), .A2(_06660_ ), .ZN(_06661_ ) );
AND4_X4 _13956_ ( .A1(_06656_ ), .A2(_06657_ ), .A3(_06658_ ), .A4(_06661_ ), .ZN(_06662_ ) );
OAI21_X2 _13957_ ( .A(_06625_ ), .B1(_06662_ ), .B2(_06106_ ), .ZN(_06663_ ) );
NAND2_X1 _13958_ ( .A1(_06663_ ), .A2(_06610_ ), .ZN(_06664_ ) );
OAI211_X1 _13959_ ( .A(_06109_ ), .B(_05290_ ), .C1(_06622_ ), .C2(_06624_ ), .ZN(_06665_ ) );
AOI21_X1 _13960_ ( .A(_06563_ ), .B1(_06664_ ), .B2(_06665_ ), .ZN(_06666_ ) );
MUX2_X1 _13961_ ( .A(\EXU.xrd_o [12] ), .B(_06666_ ), .S(_06395_ ), .Z(_00252_ ) );
NAND4_X1 _13962_ ( .A1(_05984_ ), .A2(_05832_ ), .A3(\EXU.mtvec_i [29] ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_06667_ ) );
AOI22_X1 _13963_ ( .A1(_06667_ ), .A2(_05835_ ), .B1(_05836_ ), .B2(_05837_ ), .ZN(_06668_ ) );
AND3_X1 _13964_ ( .A1(_04334_ ), .A2(\EXU.mcause_i [29] ), .A3(_05839_ ), .ZN(_06669_ ) );
OAI21_X1 _13965_ ( .A(_05830_ ), .B1(_06668_ ), .B2(_06669_ ), .ZN(_06670_ ) );
AOI22_X1 _13966_ ( .A1(_05516_ ), .A2(\EXU.mstatus_i [29] ), .B1(_05518_ ), .B2(\EXU.mepc_i [29] ), .ZN(_06671_ ) );
NAND2_X1 _13967_ ( .A1(_06670_ ), .A2(_06671_ ), .ZN(_06672_ ) );
AND4_X1 _13968_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_2_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_06673_ ) );
OAI22_X1 _13969_ ( .A1(_06672_ ), .A2(_06158_ ), .B1(_05525_ ), .B2(_06673_ ), .ZN(_06674_ ) );
AOI22_X1 _13970_ ( .A1(_04359_ ), .A2(\EXU.pc_i [29] ), .B1(\EXU.r1_i [29] ), .B2(_05528_ ), .ZN(_06675_ ) );
NAND2_X1 _13971_ ( .A1(_06674_ ), .A2(_06675_ ), .ZN(_06676_ ) );
NAND2_X1 _13972_ ( .A1(_05250_ ), .A2(_05850_ ), .ZN(_06677_ ) );
AOI21_X1 _13973_ ( .A(_05767_ ), .B1(_06598_ ), .B2(_06181_ ), .ZN(_06678_ ) );
AOI21_X1 _13974_ ( .A(_05804_ ), .B1(_06075_ ), .B2(_06079_ ), .ZN(_06679_ ) );
NAND2_X1 _13975_ ( .A1(_05790_ ), .A2(_05791_ ), .ZN(_06680_ ) );
MUX2_X1 _13976_ ( .A(_06680_ ), .B(_05799_ ), .S(_06049_ ), .Z(_06681_ ) );
NOR3_X1 _13977_ ( .A1(_05776_ ), .A2(_05777_ ), .A3(_04901_ ), .ZN(_06682_ ) );
AOI21_X1 _13978_ ( .A(_05602_ ), .B1(_05793_ ), .B2(_05794_ ), .ZN(_06683_ ) );
OR2_X1 _13979_ ( .A1(_06682_ ), .A2(_06683_ ), .ZN(_06684_ ) );
MUX2_X1 _13980_ ( .A(_06681_ ), .B(_06684_ ), .S(_06077_ ), .Z(_06685_ ) );
AOI21_X1 _13981_ ( .A(_06679_ ), .B1(_06685_ ), .B2(_06356_ ), .ZN(_06686_ ) );
OAI21_X1 _13982_ ( .A(_06678_ ), .B1(_06063_ ), .B2(_06686_ ), .ZN(_06687_ ) );
AOI21_X1 _13983_ ( .A(_05855_ ), .B1(_06600_ ), .B2(_05868_ ), .ZN(_06688_ ) );
NOR4_X1 _13984_ ( .A1(_06688_ ), .A2(_05591_ ), .A3(_05626_ ), .A4(_05870_ ), .ZN(_06689_ ) );
AND2_X1 _13985_ ( .A1(_06584_ ), .A2(_05807_ ), .ZN(_06690_ ) );
OAI21_X1 _13986_ ( .A(_06066_ ), .B1(_06689_ ), .B2(_06690_ ), .ZN(_06691_ ) );
AND4_X1 _13987_ ( .A1(_06158_ ), .A2(_05892_ ), .A3(_04768_ ), .A4(_04769_ ), .ZN(_06692_ ) );
OAI211_X1 _13988_ ( .A(_06313_ ), .B(_06314_ ), .C1(_04771_ ), .C2(_04770_ ), .ZN(_06693_ ) );
NAND2_X1 _13989_ ( .A1(_06693_ ), .A2(_06316_ ), .ZN(_06694_ ) );
AOI21_X1 _13990_ ( .A(_06692_ ), .B1(_06694_ ), .B2(_04772_ ), .ZN(_06695_ ) );
INV_X1 _13991_ ( .A(_04664_ ), .ZN(_06696_ ) );
NAND2_X1 _13992_ ( .A1(_05706_ ), .A2(_04678_ ), .ZN(_06697_ ) );
NOR3_X1 _13993_ ( .A1(_05712_ ), .A2(_05713_ ), .A3(_05715_ ), .ZN(_06698_ ) );
AOI21_X1 _13994_ ( .A(_06696_ ), .B1(_06697_ ), .B2(_06698_ ), .ZN(_06699_ ) );
OR2_X1 _13995_ ( .A1(_06699_ ), .A2(_05719_ ), .ZN(_06700_ ) );
AOI21_X1 _13996_ ( .A(_05640_ ), .B1(_06700_ ), .B2(_04663_ ), .ZN(_06701_ ) );
OAI21_X1 _13997_ ( .A(_06701_ ), .B1(_04663_ ), .B2(_06700_ ), .ZN(_06702_ ) );
AND4_X2 _13998_ ( .A1(_06687_ ), .A2(_06691_ ), .A3(_06695_ ), .A4(_06702_ ), .ZN(_06703_ ) );
AOI21_X1 _13999_ ( .A(_05849_ ), .B1(_06677_ ), .B2(_06703_ ), .ZN(_06704_ ) );
AND2_X1 _14000_ ( .A1(_05246_ ), .A2(_06500_ ), .ZN(_06705_ ) );
NAND2_X1 _14001_ ( .A1(_06672_ ), .A2(_05044_ ), .ZN(_06706_ ) );
NAND3_X1 _14002_ ( .A1(_05967_ ), .A2(_05968_ ), .A3(\EXU.imm_i [29] ), .ZN(_06707_ ) );
NAND3_X1 _14003_ ( .A1(_05970_ ), .A2(\EXU.ls_rdata_i [29] ), .A3(_05971_ ), .ZN(_06708_ ) );
NAND3_X1 _14004_ ( .A1(_06706_ ), .A2(_06707_ ), .A3(_06708_ ), .ZN(_06709_ ) );
OR3_X2 _14005_ ( .A1(_06704_ ), .A2(_06705_ ), .A3(_06709_ ), .ZN(_06710_ ) );
MUX2_X1 _14006_ ( .A(_06676_ ), .B(_06710_ ), .S(_05822_ ), .Z(_06711_ ) );
NAND2_X1 _14007_ ( .A1(_06711_ ), .A2(_06610_ ), .ZN(_06712_ ) );
NAND3_X1 _14008_ ( .A1(_04377_ ), .A2(_05977_ ), .A3(_06676_ ), .ZN(_06713_ ) );
AOI21_X1 _14009_ ( .A(_06563_ ), .B1(_06712_ ), .B2(_06713_ ), .ZN(_06714_ ) );
MUX2_X1 _14010_ ( .A(\EXU.xrd_o [29] ), .B(_06714_ ), .S(_06395_ ), .Z(_00253_ ) );
NAND2_X1 _14011_ ( .A1(_05258_ ), .A2(_06015_ ), .ZN(_06715_ ) );
OAI21_X1 _14012_ ( .A(_04699_ ), .B1(_05653_ ), .B2(_05661_ ), .ZN(_06716_ ) );
NAND2_X1 _14013_ ( .A1(_06716_ ), .A2(_05673_ ), .ZN(_06717_ ) );
AOI21_X1 _14014_ ( .A(_05677_ ), .B1(_06717_ ), .B2(_04695_ ), .ZN(_06718_ ) );
XNOR2_X1 _14015_ ( .A(_06718_ ), .B(_04694_ ), .ZN(_06719_ ) );
NAND2_X1 _14016_ ( .A1(_06719_ ), .A2(_06023_ ), .ZN(_06720_ ) );
OAI211_X1 _14017_ ( .A(_06550_ ), .B(_05521_ ), .C1(_06027_ ), .C2(_06153_ ), .ZN(_06721_ ) );
INV_X1 _14018_ ( .A(_05605_ ), .ZN(_06722_ ) );
INV_X1 _14019_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_3_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_06723_ ) );
OR3_X1 _14020_ ( .A1(_06032_ ), .A2(_06723_ ), .A3(_06034_ ), .ZN(_06724_ ) );
OAI21_X1 _14021_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_4_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_06033_ ), .B2(_06035_ ), .ZN(_06725_ ) );
NAND2_X1 _14022_ ( .A1(_06724_ ), .A2(_06725_ ), .ZN(_06726_ ) );
MUX2_X1 _14023_ ( .A(_06726_ ), .B(_06058_ ), .S(_05604_ ), .Z(_06727_ ) );
MUX2_X1 _14024_ ( .A(_06722_ ), .B(_06727_ ), .S(_05802_ ), .Z(_06728_ ) );
OR2_X1 _14025_ ( .A1(_06728_ ), .A2(_06060_ ), .ZN(_06729_ ) );
OAI21_X1 _14026_ ( .A(_06721_ ), .B1(_06729_ ), .B2(_06091_ ), .ZN(_06730_ ) );
BUF_X2 _14027_ ( .A(_06181_ ), .Z(_06731_ ) );
AOI21_X1 _14028_ ( .A(_06030_ ), .B1(_06471_ ), .B2(_06472_ ), .ZN(_06732_ ) );
NOR2_X2 _14029_ ( .A1(_05601_ ), .A2(\EXU.r1_i [11] ), .ZN(_06733_ ) );
NOR3_X1 _14030_ ( .A1(_06160_ ), .A2(\EXU.r1_i [12] ), .A3(_06047_ ), .ZN(_06734_ ) );
NOR2_X1 _14031_ ( .A1(_06733_ ), .A2(_06734_ ), .ZN(_06735_ ) );
NOR2_X1 _14032_ ( .A1(_06575_ ), .A2(_06576_ ), .ZN(_06736_ ) );
MUX2_X2 _14033_ ( .A(_06735_ ), .B(_06736_ ), .S(_05604_ ), .Z(_06737_ ) );
AOI21_X1 _14034_ ( .A(_06732_ ), .B1(_06526_ ), .B2(_06737_ ), .ZN(_06738_ ) );
OR2_X1 _14035_ ( .A1(_06738_ ), .A2(_06081_ ), .ZN(_06739_ ) );
NAND3_X1 _14036_ ( .A1(_06226_ ), .A2(_06232_ ), .A3(_06081_ ), .ZN(_06740_ ) );
AOI21_X1 _14037_ ( .A(_06731_ ), .B1(_06739_ ), .B2(_06740_ ), .ZN(_06741_ ) );
OAI21_X1 _14038_ ( .A(_06538_ ), .B1(_06730_ ), .B2(_06741_ ), .ZN(_06742_ ) );
NOR2_X1 _14039_ ( .A1(_06253_ ), .A2(_05960_ ), .ZN(_06743_ ) );
NOR3_X1 _14040_ ( .A1(_05764_ ), .A2(_05747_ ), .A3(_06077_ ), .ZN(_06744_ ) );
OAI21_X1 _14041_ ( .A(_06495_ ), .B1(_06743_ ), .B2(_06744_ ), .ZN(_06745_ ) );
NAND4_X1 _14042_ ( .A1(_04427_ ), .A2(_04840_ ), .A3(_04842_ ), .A4(_04843_ ), .ZN(_06746_ ) );
NAND3_X1 _14043_ ( .A1(_04842_ ), .A2(\EXU.r1_i [11] ), .A3(_04843_ ), .ZN(_06747_ ) );
AOI21_X1 _14044_ ( .A(_05555_ ), .B1(_05573_ ), .B2(_06747_ ), .ZN(_06748_ ) );
AND2_X1 _14045_ ( .A1(_04844_ ), .A2(_04841_ ), .ZN(_06749_ ) );
OR2_X1 _14046_ ( .A1(_06748_ ), .A2(_06749_ ), .ZN(_06750_ ) );
MUX2_X1 _14047_ ( .A(_06746_ ), .B(_06750_ ), .S(_06071_ ), .Z(_06751_ ) );
AND4_X1 _14048_ ( .A1(_06720_ ), .A2(_06742_ ), .A3(_06745_ ), .A4(_06751_ ), .ZN(_06752_ ) );
AOI21_X1 _14049_ ( .A(_06014_ ), .B1(_06715_ ), .B2(_06752_ ), .ZN(_06753_ ) );
AND2_X1 _14050_ ( .A1(_05262_ ), .A2(_05039_ ), .ZN(_06754_ ) );
NAND4_X1 _14051_ ( .A1(_05984_ ), .A2(_05832_ ), .A3(\EXU.mtvec_i [11] ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_06755_ ) );
AOI22_X1 _14052_ ( .A1(_06755_ ), .A2(_05835_ ), .B1(_05839_ ), .B2(_05837_ ), .ZN(_06756_ ) );
AND3_X1 _14053_ ( .A1(_04334_ ), .A2(\EXU.mcause_i [11] ), .A3(_05839_ ), .ZN(_06757_ ) );
OAI21_X1 _14054_ ( .A(_05829_ ), .B1(_06756_ ), .B2(_06757_ ), .ZN(_06758_ ) );
NAND3_X1 _14055_ ( .A1(_06204_ ), .A2(_06208_ ), .A3(\EXU.mepc_i [11] ), .ZN(_06759_ ) );
NAND3_X1 _14056_ ( .A1(_06206_ ), .A2(\EXU.mstatus_i [11] ), .A3(_05988_ ), .ZN(_06760_ ) );
AND3_X1 _14057_ ( .A1(_06758_ ), .A2(_06759_ ), .A3(_06760_ ), .ZN(_06761_ ) );
OR2_X1 _14058_ ( .A1(_06761_ ), .A2(_06011_ ), .ZN(_06762_ ) );
INV_X1 _14059_ ( .A(_06008_ ), .ZN(_06763_ ) );
INV_X1 _14060_ ( .A(\EXU.ls_rdata_i [11] ), .ZN(_06764_ ) );
OAI221_X1 _14061_ ( .A(_06762_ ), .B1(_04344_ ), .B2(_06763_ ), .C1(_06764_ ), .C2(_04414_ ), .ZN(_06765_ ) );
OR3_X1 _14062_ ( .A1(_06753_ ), .A2(_06754_ ), .A3(_06765_ ), .ZN(_06766_ ) );
XNOR2_X1 _14063_ ( .A(_04371_ ), .B(_04372_ ), .ZN(_06767_ ) );
NAND2_X1 _14064_ ( .A1(_06766_ ), .A2(_06767_ ), .ZN(_06768_ ) );
AOI21_X1 _14065_ ( .A(_05995_ ), .B1(_06761_ ), .B2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_20_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_06769_ ) );
NOR3_X1 _14066_ ( .A1(_06761_ ), .A2(_04840_ ), .A3(_05560_ ), .ZN(_06770_ ) );
AOI211_X1 _14067_ ( .A(_06769_ ), .B(_06770_ ), .C1(\EXU.r1_i [11] ), .C2(_05528_ ), .ZN(_06771_ ) );
NAND3_X1 _14068_ ( .A1(_05045_ ), .A2(\EXU.pc_i [11] ), .A3(_05092_ ), .ZN(_06772_ ) );
NAND2_X1 _14069_ ( .A1(_06771_ ), .A2(_06772_ ), .ZN(_06773_ ) );
AND2_X1 _14070_ ( .A1(_04376_ ), .A2(_05050_ ), .ZN(_06774_ ) );
OAI21_X1 _14071_ ( .A(_06773_ ), .B1(_06774_ ), .B2(_06106_ ), .ZN(_06775_ ) );
AOI21_X1 _14072_ ( .A(_06563_ ), .B1(_06768_ ), .B2(_06775_ ), .ZN(_06776_ ) );
MUX2_X1 _14073_ ( .A(\EXU.xrd_o [11] ), .B(_06776_ ), .S(_06395_ ), .Z(_00254_ ) );
XOR2_X1 _14074_ ( .A(_06717_ ), .B(_04695_ ), .Z(_06777_ ) );
AND2_X1 _14075_ ( .A1(_06777_ ), .A2(_06023_ ), .ZN(_06778_ ) );
NOR3_X1 _14076_ ( .A1(_05923_ ), .A2(_05747_ ), .A3(_06077_ ), .ZN(_06779_ ) );
AOI21_X1 _14077_ ( .A(_06779_ ), .B1(_05880_ ), .B2(_06283_ ), .ZN(_06780_ ) );
NOR2_X1 _14078_ ( .A1(_06780_ ), .A2(_06542_ ), .ZN(_06781_ ) );
OAI211_X1 _14079_ ( .A(_06313_ ), .B(_06314_ ), .C1(_04849_ ), .C2(_04848_ ), .ZN(_06782_ ) );
NAND2_X1 _14080_ ( .A1(_06782_ ), .A2(_06316_ ), .ZN(_06783_ ) );
AND2_X1 _14081_ ( .A1(_06783_ ), .A2(_04850_ ), .ZN(_06784_ ) );
NOR3_X1 _14082_ ( .A1(_06071_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_21_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A3(_04848_ ), .ZN(_06785_ ) );
NOR4_X1 _14083_ ( .A1(_06778_ ), .A2(_06781_ ), .A3(_06784_ ), .A4(_06785_ ), .ZN(_06786_ ) );
INV_X1 _14084_ ( .A(_05584_ ), .ZN(_06787_ ) );
OAI21_X1 _14085_ ( .A(_06786_ ), .B1(_05270_ ), .B2(_06787_ ), .ZN(_06788_ ) );
NAND3_X1 _14086_ ( .A1(_06525_ ), .A2(_06289_ ), .A3(_06530_ ), .ZN(_06789_ ) );
OAI21_X1 _14087_ ( .A(_05878_ ), .B1(_06630_ ), .B2(_06631_ ), .ZN(_06790_ ) );
OR3_X1 _14088_ ( .A1(_06046_ ), .A2(_04841_ ), .A3(_06050_ ), .ZN(_06791_ ) );
OAI21_X1 _14089_ ( .A(\EXU.r1_i [10] ), .B1(_06527_ ), .B2(_06528_ ), .ZN(_06792_ ) );
NAND3_X1 _14090_ ( .A1(_06791_ ), .A2(_06414_ ), .A3(_06792_ ), .ZN(_06793_ ) );
AND2_X1 _14091_ ( .A1(_06790_ ), .A2(_06793_ ), .ZN(_06794_ ) );
OAI21_X1 _14092_ ( .A(_06789_ ), .B1(_06794_ ), .B2(_06289_ ), .ZN(_06795_ ) );
MUX2_X1 _14093_ ( .A(_06795_ ), .B(_06309_ ), .S(_06100_ ), .Z(_06796_ ) );
OR2_X1 _14094_ ( .A1(_06796_ ), .A2(_06731_ ), .ZN(_06797_ ) );
OAI21_X1 _14095_ ( .A(_05866_ ), .B1(_05861_ ), .B2(_05863_ ), .ZN(_06798_ ) );
AND3_X1 _14096_ ( .A1(_06798_ ), .A2(_05868_ ), .A3(_06550_ ), .ZN(_06799_ ) );
NOR2_X1 _14097_ ( .A1(_05601_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_5_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_06800_ ) );
NOR3_X1 _14098_ ( .A1(_06160_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_4_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A3(_06047_ ), .ZN(_06801_ ) );
NOR2_X1 _14099_ ( .A1(_06800_ ), .A2(_06801_ ), .ZN(_06802_ ) );
MUX2_X1 _14100_ ( .A(_06162_ ), .B(_06802_ ), .S(_05938_ ), .Z(_06803_ ) );
AND2_X1 _14101_ ( .A1(_06803_ ), .A2(_05934_ ), .ZN(_06804_ ) );
OAI21_X1 _14102_ ( .A(_05747_ ), .B1(_05879_ ), .B2(_05934_ ), .ZN(_06805_ ) );
NOR2_X1 _14103_ ( .A1(_06804_ ), .A2(_06805_ ), .ZN(_06806_ ) );
AOI21_X1 _14104_ ( .A(_06799_ ), .B1(_06806_ ), .B2(_06731_ ), .ZN(_06807_ ) );
AOI21_X1 _14105_ ( .A(_05852_ ), .B1(_06797_ ), .B2(_06807_ ), .ZN(_06808_ ) );
OAI21_X1 _14106_ ( .A(_06626_ ), .B1(_06788_ ), .B2(_06808_ ), .ZN(_06809_ ) );
INV_X1 _14107_ ( .A(\EXU.ls_rdata_i [10] ), .ZN(_06810_ ) );
OAI22_X1 _14108_ ( .A1(_04414_ ), .A2(_06810_ ), .B1(_06763_ ), .B2(_05545_ ), .ZN(_06811_ ) );
AOI22_X1 _14109_ ( .A1(_05516_ ), .A2(\EXU.mstatus_i [10] ), .B1(_05518_ ), .B2(\EXU.mepc_i [10] ), .ZN(_06812_ ) );
NAND3_X1 _14110_ ( .A1(_06206_ ), .A2(\EXU.mtvec_i [10] ), .A3(_06208_ ), .ZN(_06813_ ) );
NAND3_X1 _14111_ ( .A1(_06203_ ), .A2(\EXU.mcause_i [10] ), .A3(_06204_ ), .ZN(_06814_ ) );
AND3_X1 _14112_ ( .A1(_06812_ ), .A2(_06813_ ), .A3(_06814_ ), .ZN(_06815_ ) );
NOR2_X1 _14113_ ( .A1(_06815_ ), .A2(_06012_ ), .ZN(_06816_ ) );
AOI211_X1 _14114_ ( .A(_06811_ ), .B(_06816_ ), .C1(_05211_ ), .C2(_05272_ ), .ZN(_06817_ ) );
NAND2_X1 _14115_ ( .A1(_06809_ ), .A2(_06817_ ), .ZN(_06818_ ) );
NAND2_X1 _14116_ ( .A1(_06818_ ), .A2(_06767_ ), .ZN(_06819_ ) );
NAND4_X1 _14117_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_21_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_06820_ ) );
AOI22_X1 _14118_ ( .A1(_06815_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_21_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_05996_ ), .B2(_06820_ ), .ZN(_06821_ ) );
NAND3_X1 _14119_ ( .A1(_05045_ ), .A2(\EXU.pc_i [10] ), .A3(_05047_ ), .ZN(_06822_ ) );
OAI21_X1 _14120_ ( .A(_06822_ ), .B1(_04849_ ), .B2(_06003_ ), .ZN(_06823_ ) );
OAI22_X1 _14121_ ( .A1(_06774_ ), .A2(_06106_ ), .B1(_06821_ ), .B2(_06823_ ), .ZN(_06824_ ) );
AOI21_X1 _14122_ ( .A(_06563_ ), .B1(_06819_ ), .B2(_06824_ ), .ZN(_06825_ ) );
MUX2_X1 _14123_ ( .A(\EXU.xrd_o [10] ), .B(_06825_ ), .S(_06395_ ), .Z(_00255_ ) );
NAND3_X1 _14124_ ( .A1(_06203_ ), .A2(\EXU.mcause_i [9] ), .A3(_05836_ ), .ZN(_06826_ ) );
NAND3_X1 _14125_ ( .A1(_06118_ ), .A2(\EXU.mstatus_i [9] ), .A3(_05988_ ), .ZN(_06827_ ) );
NAND3_X1 _14126_ ( .A1(_06118_ ), .A2(\EXU.mtvec_i [9] ), .A3(_05831_ ), .ZN(_06828_ ) );
NAND4_X1 _14127_ ( .A1(_06202_ ), .A2(_06826_ ), .A3(_06827_ ), .A4(_06828_ ), .ZN(_06829_ ) );
OR2_X1 _14128_ ( .A1(_05992_ ), .A2(\EXU.mepc_i [9] ), .ZN(_06830_ ) );
NAND2_X1 _14129_ ( .A1(_06829_ ), .A2(_06830_ ), .ZN(_06831_ ) );
NAND4_X1 _14130_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_22_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_06832_ ) );
AOI22_X1 _14131_ ( .A1(_06831_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_22_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_05557_ ), .B2(_06832_ ), .ZN(_06833_ ) );
NAND3_X1 _14132_ ( .A1(_06123_ ), .A2(\EXU.pc_i [9] ), .A3(_04348_ ), .ZN(_06834_ ) );
OAI21_X1 _14133_ ( .A(_06834_ ), .B1(_04918_ ), .B2(_06002_ ), .ZN(_06835_ ) );
OR2_X1 _14134_ ( .A1(_06833_ ), .A2(_06835_ ), .ZN(_06836_ ) );
AOI21_X1 _14135_ ( .A(_05670_ ), .B1(_06481_ ), .B2(_04698_ ), .ZN(_06837_ ) );
XNOR2_X1 _14136_ ( .A(_06837_ ), .B(_04697_ ), .ZN(_06838_ ) );
NAND2_X1 _14137_ ( .A1(_06838_ ), .A2(_05639_ ), .ZN(_06839_ ) );
NAND3_X1 _14138_ ( .A1(_04915_ ), .A2(\EXU.r1_i [9] ), .A3(_04916_ ), .ZN(_06840_ ) );
AOI21_X1 _14139_ ( .A(_05555_ ), .B1(_05573_ ), .B2(_06840_ ), .ZN(_06841_ ) );
OR2_X1 _14140_ ( .A1(_06841_ ), .A2(_04919_ ), .ZN(_06842_ ) );
NAND2_X1 _14141_ ( .A1(_04920_ ), .A2(_06186_ ), .ZN(_06843_ ) );
AOI21_X1 _14142_ ( .A(_04886_ ), .B1(_06376_ ), .B2(_06377_ ), .ZN(_06844_ ) );
NOR4_X1 _14143_ ( .A1(_05763_ ), .A2(_04885_ ), .A3(_04996_ ), .A4(_05604_ ), .ZN(_06845_ ) );
OAI21_X1 _14144_ ( .A(_06495_ ), .B1(_06844_ ), .B2(_06845_ ), .ZN(_06846_ ) );
NAND4_X1 _14145_ ( .A1(_06839_ ), .A2(_06842_ ), .A3(_06843_ ), .A4(_06846_ ), .ZN(_06847_ ) );
AOI21_X1 _14146_ ( .A(_06847_ ), .B1(_05280_ ), .B2(_05585_ ), .ZN(_06848_ ) );
AOI21_X1 _14147_ ( .A(_06049_ ), .B1(_06724_ ), .B2(_06725_ ), .ZN(_06849_ ) );
MUX2_X1 _14148_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_6_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B(\EXU.xrd_o_$_SDFFCE_PP0P__Q_5_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .S(_06040_ ), .Z(_06850_ ) );
AOI211_X1 _14149_ ( .A(_06096_ ), .B(_06849_ ), .C1(_06850_ ), .C2(_06144_ ), .ZN(_06851_ ) );
AND2_X1 _14150_ ( .A1(_06059_ ), .A2(_06077_ ), .ZN(_06852_ ) );
OAI211_X1 _14151_ ( .A(_06063_ ), .B(_06356_ ), .C1(_06851_ ), .C2(_06852_ ), .ZN(_06853_ ) );
NOR2_X1 _14152_ ( .A1(_05865_ ), .A2(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ), .ZN(_06854_ ) );
OAI21_X1 _14153_ ( .A(_06549_ ), .B1(_06363_ ), .B2(_06854_ ), .ZN(_06855_ ) );
AOI21_X1 _14154_ ( .A(_06356_ ), .B1(_06355_ ), .B2(_06358_ ), .ZN(_06856_ ) );
OR3_X1 _14155_ ( .A1(_06032_ ), .A2(_04849_ ), .A3(_06034_ ), .ZN(_06857_ ) );
OAI21_X1 _14156_ ( .A(\EXU.r1_i [9] ), .B1(_06160_ ), .B2(_06047_ ), .ZN(_06858_ ) );
NAND2_X1 _14157_ ( .A1(_06857_ ), .A2(_06858_ ), .ZN(_06859_ ) );
MUX2_X1 _14158_ ( .A(_06859_ ), .B(_06735_ ), .S(_06039_ ), .Z(_06860_ ) );
MUX2_X1 _14159_ ( .A(_06579_ ), .B(_06860_ ), .S(_05881_ ), .Z(_06861_ ) );
AOI21_X1 _14160_ ( .A(_06856_ ), .B1(_06861_ ), .B2(_06532_ ), .ZN(_06862_ ) );
OAI211_X1 _14161_ ( .A(_06853_ ), .B(_06855_ ), .C1(_06862_ ), .C2(_06731_ ), .ZN(_06863_ ) );
NAND2_X1 _14162_ ( .A1(_06863_ ), .A2(_06066_ ), .ZN(_06864_ ) );
AOI21_X1 _14163_ ( .A(_05535_ ), .B1(_06848_ ), .B2(_06864_ ), .ZN(_06865_ ) );
AND2_X1 _14164_ ( .A1(_05284_ ), .A2(_06500_ ), .ZN(_06866_ ) );
AND3_X1 _14165_ ( .A1(_06829_ ), .A2(_05044_ ), .A3(_06830_ ), .ZN(_06867_ ) );
NAND3_X1 _14166_ ( .A1(_04387_ ), .A2(\EXU.ls_rdata_i [9] ), .A3(_04388_ ), .ZN(_06868_ ) );
OAI21_X1 _14167_ ( .A(_06868_ ), .B1(_06763_ ), .B2(_04346_ ), .ZN(_06869_ ) );
OR4_X1 _14168_ ( .A1(_06865_ ), .A2(_06866_ ), .A3(_06867_ ), .A4(_06869_ ), .ZN(_06870_ ) );
MUX2_X1 _14169_ ( .A(_06836_ ), .B(_06870_ ), .S(_05822_ ), .Z(_06871_ ) );
NAND2_X1 _14170_ ( .A1(_06871_ ), .A2(_06610_ ), .ZN(_06872_ ) );
NAND3_X1 _14171_ ( .A1(_04377_ ), .A2(_05977_ ), .A3(_06836_ ), .ZN(_06873_ ) );
AOI21_X1 _14172_ ( .A(_06563_ ), .B1(_06872_ ), .B2(_06873_ ), .ZN(_06874_ ) );
MUX2_X1 _14173_ ( .A(\EXU.xrd_o [9] ), .B(_06874_ ), .S(_06395_ ), .Z(_00256_ ) );
AND3_X1 _14174_ ( .A1(_06118_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_23_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05831_ ), .ZN(_06875_ ) );
OAI221_X1 _14175_ ( .A(_05830_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_23_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05981_ ), .C1(_05983_ ), .C2(_06875_ ), .ZN(_06876_ ) );
NAND4_X1 _14176_ ( .A1(_05987_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_23_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_05989_ ), .ZN(_06877_ ) );
NAND2_X1 _14177_ ( .A1(_06876_ ), .A2(_06877_ ), .ZN(_06878_ ) );
MUX2_X1 _14178_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_23_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ), .B(_06878_ ), .S(_05993_ ), .Z(_06879_ ) );
NAND4_X1 _14179_ ( .A1(_04926_ ), .A2(fanout_net_6 ), .A3(fanout_net_5 ), .A4(fanout_net_10 ), .ZN(_06880_ ) );
AOI22_X1 _14180_ ( .A1(_06879_ ), .A2(_04926_ ), .B1(_05996_ ), .B2(_06880_ ), .ZN(_06881_ ) );
NAND3_X1 _14181_ ( .A1(_06516_ ), .A2(\EXU.pc_i [8] ), .A3(_05999_ ), .ZN(_06882_ ) );
OAI21_X1 _14182_ ( .A(_06882_ ), .B1(_04926_ ), .B2(_06003_ ), .ZN(_06883_ ) );
OAI211_X1 _14183_ ( .A(_04371_ ), .B(_04374_ ), .C1(_06881_ ), .C2(_06883_ ), .ZN(_06884_ ) );
AND3_X1 _14184_ ( .A1(_06632_ ), .A2(_06357_ ), .A3(_06633_ ), .ZN(_06885_ ) );
OR3_X1 _14185_ ( .A1(_06527_ ), .A2(_04918_ ), .A3(_06528_ ), .ZN(_06886_ ) );
OAI21_X1 _14186_ ( .A(\EXU.r1_i [8] ), .B1(_06527_ ), .B2(_06528_ ), .ZN(_06887_ ) );
NAND3_X1 _14187_ ( .A1(_06886_ ), .A2(_06414_ ), .A3(_06887_ ), .ZN(_06888_ ) );
NAND3_X1 _14188_ ( .A1(_06791_ ), .A2(_05878_ ), .A3(_06792_ ), .ZN(_06889_ ) );
AOI21_X1 _14189_ ( .A(_06357_ ), .B1(_06888_ ), .B2(_06889_ ), .ZN(_06890_ ) );
NOR2_X1 _14190_ ( .A1(_06885_ ), .A2(_06890_ ), .ZN(_06891_ ) );
MUX2_X1 _14191_ ( .A(_06424_ ), .B(_06891_ ), .S(_06532_ ), .Z(_06892_ ) );
NAND2_X1 _14192_ ( .A1(_06892_ ), .A2(_06361_ ), .ZN(_06893_ ) );
NAND2_X1 _14193_ ( .A1(_06409_ ), .A2(_05866_ ), .ZN(_06894_ ) );
NAND3_X1 _14194_ ( .A1(_06894_ ), .A2(_05868_ ), .A3(_06550_ ), .ZN(_06895_ ) );
MUX2_X1 _14195_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ), .B(\EXU.xrd_o_$_SDFFCE_PP0P__Q_6_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .S(_05601_ ), .Z(_06896_ ) );
MUX2_X1 _14196_ ( .A(_06802_ ), .B(_06896_ ), .S(_06049_ ), .Z(_06897_ ) );
MUX2_X1 _14197_ ( .A(_06639_ ), .B(_06897_ ), .S(_05934_ ), .Z(_06898_ ) );
OR2_X1 _14198_ ( .A1(_06898_ ), .A2(_06099_ ), .ZN(_06899_ ) );
OAI211_X1 _14199_ ( .A(_06893_ ), .B(_06895_ ), .C1(_06899_ ), .C2(_06361_ ), .ZN(_06900_ ) );
NAND2_X1 _14200_ ( .A1(_06900_ ), .A2(_06538_ ), .ZN(_06901_ ) );
XNOR2_X1 _14201_ ( .A(_06480_ ), .B(_04698_ ), .ZN(_06902_ ) );
AND3_X1 _14202_ ( .A1(_06902_ ), .A2(_05583_ ), .A3(_05638_ ), .ZN(_06903_ ) );
NAND4_X1 _14203_ ( .A1(_04998_ ), .A2(_05960_ ), .A3(_06030_ ), .A4(_06414_ ), .ZN(_06904_ ) );
OAI21_X1 _14204_ ( .A(_06904_ ), .B1(_06442_ ), .B2(_06060_ ), .ZN(_06905_ ) );
AND2_X1 _14205_ ( .A1(_06905_ ), .A2(_06495_ ), .ZN(_06906_ ) );
OAI211_X1 _14206_ ( .A(_05887_ ), .B(_05888_ ), .C1(_04926_ ), .C2(_04924_ ), .ZN(_06907_ ) );
NAND2_X1 _14207_ ( .A1(_06907_ ), .A2(_05890_ ), .ZN(_06908_ ) );
AND2_X1 _14208_ ( .A1(_06908_ ), .A2(_04927_ ), .ZN(_06909_ ) );
NOR2_X1 _14209_ ( .A1(_04925_ ), .A2(_06071_ ), .ZN(_06910_ ) );
OR4_X1 _14210_ ( .A1(_06903_ ), .A2(_06906_ ), .A3(_06909_ ), .A4(_06910_ ), .ZN(_06911_ ) );
AOI21_X1 _14211_ ( .A(_06911_ ), .B1(_05295_ ), .B2(_06015_ ), .ZN(_06912_ ) );
AOI21_X1 _14212_ ( .A(_06014_ ), .B1(_06901_ ), .B2(_06912_ ), .ZN(_06913_ ) );
NOR2_X1 _14213_ ( .A1(_06879_ ), .A2(_06012_ ), .ZN(_06914_ ) );
AND2_X1 _14214_ ( .A1(_05292_ ), .A2(_05039_ ), .ZN(_06915_ ) );
NAND3_X1 _14215_ ( .A1(_05967_ ), .A2(_05968_ ), .A3(\EXU.imm_i [8] ), .ZN(_06916_ ) );
INV_X1 _14216_ ( .A(\EXU.ls_rdata_i [8] ), .ZN(_06917_ ) );
OAI21_X1 _14217_ ( .A(_06916_ ), .B1(_04414_ ), .B2(_06917_ ), .ZN(_06918_ ) );
NOR4_X1 _14218_ ( .A1(_06913_ ), .A2(_06914_ ), .A3(_06915_ ), .A4(_06918_ ), .ZN(_06919_ ) );
OAI21_X1 _14219_ ( .A(_06884_ ), .B1(_06919_ ), .B2(_06106_ ), .ZN(_06920_ ) );
NAND2_X1 _14220_ ( .A1(_06920_ ), .A2(_06610_ ), .ZN(_06921_ ) );
OAI211_X1 _14221_ ( .A(_06109_ ), .B(_05290_ ), .C1(_06881_ ), .C2(_06883_ ), .ZN(_06922_ ) );
AOI21_X1 _14222_ ( .A(_06563_ ), .B1(_06921_ ), .B2(_06922_ ), .ZN(_06923_ ) );
BUF_X4 _14223_ ( .A(_04399_ ), .Z(_06924_ ) );
MUX2_X1 _14224_ ( .A(\EXU.xrd_o [8] ), .B(_06923_ ), .S(_06924_ ), .Z(_00257_ ) );
NAND3_X1 _14225_ ( .A1(_06203_ ), .A2(\EXU.mcause_i [7] ), .A3(_06204_ ), .ZN(_06925_ ) );
NAND3_X1 _14226_ ( .A1(_06206_ ), .A2(\EXU.mstatus_i [7] ), .A3(_05988_ ), .ZN(_06926_ ) );
NAND3_X1 _14227_ ( .A1(_06206_ ), .A2(\EXU.mtvec_i [7] ), .A3(_06208_ ), .ZN(_06927_ ) );
NAND4_X1 _14228_ ( .A1(_06202_ ), .A2(_06925_ ), .A3(_06926_ ), .A4(_06927_ ), .ZN(_06928_ ) );
OAI21_X1 _14229_ ( .A(_06928_ ), .B1(\EXU.mepc_i [7] ), .B2(_05993_ ), .ZN(_06929_ ) );
NAND4_X1 _14230_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_24_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_06930_ ) );
AOI22_X1 _14231_ ( .A1(_06929_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_24_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_05557_ ), .B2(_06930_ ), .ZN(_06931_ ) );
NAND3_X1 _14232_ ( .A1(_06123_ ), .A2(\EXU.pc_i [7] ), .A3(_04348_ ), .ZN(_06932_ ) );
OAI21_X1 _14233_ ( .A(_06932_ ), .B1(_04930_ ), .B2(_06002_ ), .ZN(_06933_ ) );
OR2_X1 _14234_ ( .A1(_06931_ ), .A2(_06933_ ), .ZN(_06934_ ) );
NOR2_X2 _14235_ ( .A1(_05601_ ), .A2(\EXU.r1_i [7] ), .ZN(_06935_ ) );
NOR3_X1 _14236_ ( .A1(_06160_ ), .A2(\EXU.r1_i [8] ), .A3(_06047_ ), .ZN(_06936_ ) );
NOR2_X1 _14237_ ( .A1(_06935_ ), .A2(_06936_ ), .ZN(_06937_ ) );
MUX2_X2 _14238_ ( .A(_06859_ ), .B(_06937_ ), .S(_05938_ ), .Z(_06938_ ) );
MUX2_X2 _14239_ ( .A(_06938_ ), .B(_06737_ ), .S(_06096_ ), .Z(_06939_ ) );
MUX2_X2 _14240_ ( .A(_06474_ ), .B(_06939_ ), .S(_05880_ ), .Z(_06940_ ) );
OR2_X2 _14241_ ( .A1(_06940_ ), .A2(_06063_ ), .ZN(_06941_ ) );
NAND3_X1 _14242_ ( .A1(_05605_ ), .A2(_06060_ ), .A3(_05881_ ), .ZN(_06942_ ) );
OAI21_X1 _14243_ ( .A(_06942_ ), .B1(_06466_ ), .B2(_06099_ ), .ZN(_06943_ ) );
OAI211_X1 _14244_ ( .A(_06941_ ), .B(_06538_ ), .C1(_06361_ ), .C2(_06943_ ), .ZN(_06944_ ) );
NAND2_X1 _14245_ ( .A1(_06854_ ), .A2(_06549_ ), .ZN(_06945_ ) );
AND2_X1 _14246_ ( .A1(_05652_ ), .A2(_04672_ ), .ZN(_06946_ ) );
OAI21_X1 _14247_ ( .A(_04668_ ), .B1(_06946_ ), .B2(_05656_ ), .ZN(_06947_ ) );
NAND2_X1 _14248_ ( .A1(_06947_ ), .A2(_05659_ ), .ZN(_06948_ ) );
XNOR2_X1 _14249_ ( .A(_06948_ ), .B(_05658_ ), .ZN(_06949_ ) );
NAND2_X1 _14250_ ( .A1(_06023_ ), .A2(_06949_ ), .ZN(_06950_ ) );
NAND2_X1 _14251_ ( .A1(_05764_ ), .A2(_05924_ ), .ZN(_06951_ ) );
NAND3_X1 _14252_ ( .A1(_05751_ ), .A2(_05753_ ), .A3(_05802_ ), .ZN(_06952_ ) );
NAND4_X1 _14253_ ( .A1(_06951_ ), .A2(_06356_ ), .A3(_06952_ ), .A4(_06495_ ), .ZN(_06953_ ) );
OAI21_X1 _14254_ ( .A(_05892_ ), .B1(_04933_ ), .B2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_24_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_06954_ ) );
OAI211_X1 _14255_ ( .A(_05887_ ), .B(_05888_ ), .C1(_04930_ ), .C2(_04933_ ), .ZN(_06955_ ) );
AOI22_X1 _14256_ ( .A1(_06955_ ), .A2(_05890_ ), .B1(_04930_ ), .B2(_04933_ ), .ZN(_06956_ ) );
OAI211_X1 _14257_ ( .A(_04427_ ), .B(_06954_ ), .C1(_06956_ ), .C2(_05892_ ), .ZN(_06957_ ) );
NAND4_X1 _14258_ ( .A1(_06945_ ), .A2(_06950_ ), .A3(_06953_ ), .A4(_06957_ ), .ZN(_06958_ ) );
AOI21_X1 _14259_ ( .A(_06958_ ), .B1(_05303_ ), .B2(_05585_ ), .ZN(_06959_ ) );
AOI21_X1 _14260_ ( .A(_05849_ ), .B1(_06944_ ), .B2(_06959_ ), .ZN(_06960_ ) );
NOR2_X1 _14261_ ( .A1(_06929_ ), .A2(_06011_ ), .ZN(_06961_ ) );
NAND2_X1 _14262_ ( .A1(_05300_ ), .A2(_06500_ ), .ZN(_06962_ ) );
AOI22_X1 _14263_ ( .A1(_06006_ ), .A2(\EXU.ls_rdata_i [7] ), .B1(_06009_ ), .B2(\EXU.imm_i [7] ), .ZN(_06963_ ) );
NAND2_X1 _14264_ ( .A1(_06962_ ), .A2(_06963_ ), .ZN(_06964_ ) );
OR3_X2 _14265_ ( .A1(_06960_ ), .A2(_06961_ ), .A3(_06964_ ), .ZN(_06965_ ) );
MUX2_X2 _14266_ ( .A(_06934_ ), .B(_06965_ ), .S(_05822_ ), .Z(_06966_ ) );
NAND2_X1 _14267_ ( .A1(_06966_ ), .A2(_06610_ ), .ZN(_06967_ ) );
NAND3_X1 _14268_ ( .A1(_04377_ ), .A2(_05977_ ), .A3(_06934_ ), .ZN(_06968_ ) );
AOI21_X1 _14269_ ( .A(_06563_ ), .B1(_06967_ ), .B2(_06968_ ), .ZN(_06969_ ) );
MUX2_X1 _14270_ ( .A(\EXU.xrd_o [7] ), .B(_06969_ ), .S(_06924_ ), .Z(_00258_ ) );
AND3_X1 _14271_ ( .A1(_06118_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_25_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05831_ ), .ZN(_06970_ ) );
OAI221_X1 _14272_ ( .A(_05830_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_25_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05981_ ), .C1(_05983_ ), .C2(_06970_ ), .ZN(_06971_ ) );
NAND4_X1 _14273_ ( .A1(_05987_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_25_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_05989_ ), .ZN(_06972_ ) );
NAND2_X1 _14274_ ( .A1(_06971_ ), .A2(_06972_ ), .ZN(_06973_ ) );
MUX2_X1 _14275_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_25_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ), .B(_06973_ ), .S(_05993_ ), .Z(_06974_ ) );
NAND4_X1 _14276_ ( .A1(_04940_ ), .A2(fanout_net_6 ), .A3(fanout_net_5 ), .A4(fanout_net_10 ), .ZN(_06975_ ) );
AOI22_X1 _14277_ ( .A1(_06974_ ), .A2(_04940_ ), .B1(_05996_ ), .B2(_06975_ ), .ZN(_06976_ ) );
NAND3_X1 _14278_ ( .A1(_06516_ ), .A2(\EXU.pc_i [6] ), .A3(_05999_ ), .ZN(_06977_ ) );
OAI21_X1 _14279_ ( .A(_06977_ ), .B1(_04940_ ), .B2(_06003_ ), .ZN(_06978_ ) );
OAI211_X1 _14280_ ( .A(_04371_ ), .B(_04374_ ), .C1(_06976_ ), .C2(_06978_ ), .ZN(_06979_ ) );
INV_X1 _14281_ ( .A(_06550_ ), .ZN(_06980_ ) );
OR3_X1 _14282_ ( .A1(_05864_ ), .A2(_05866_ ), .A3(_06980_ ), .ZN(_06981_ ) );
NOR3_X1 _14283_ ( .A1(_05876_ ), .A2(_06077_ ), .A3(_05878_ ), .ZN(_06982_ ) );
INV_X1 _14284_ ( .A(_06982_ ), .ZN(_06983_ ) );
MUX2_X1 _14285_ ( .A(_06983_ ), .B(_06536_ ), .S(_05804_ ), .Z(_06984_ ) );
OAI21_X1 _14286_ ( .A(_06981_ ), .B1(_06984_ ), .B2(_06361_ ), .ZN(_06985_ ) );
OR3_X1 _14287_ ( .A1(_06046_ ), .A2(\EXU.r1_i [7] ), .A3(_06050_ ), .ZN(_06986_ ) );
OAI21_X1 _14288_ ( .A(_04940_ ), .B1(_06046_ ), .B2(_06528_ ), .ZN(_06987_ ) );
NAND2_X1 _14289_ ( .A1(_06986_ ), .A2(_06987_ ), .ZN(_06988_ ) );
NAND2_X1 _14290_ ( .A1(_06988_ ), .A2(_06414_ ), .ZN(_06989_ ) );
NAND3_X1 _14291_ ( .A1(_06886_ ), .A2(_06383_ ), .A3(_06887_ ), .ZN(_06990_ ) );
NAND2_X1 _14292_ ( .A1(_06989_ ), .A2(_06990_ ), .ZN(_06991_ ) );
NAND2_X1 _14293_ ( .A1(_06991_ ), .A2(_06526_ ), .ZN(_06992_ ) );
OAI211_X1 _14294_ ( .A(_06992_ ), .B(_06532_ ), .C1(_06526_ ), .C2(_06794_ ), .ZN(_06993_ ) );
NAND3_X1 _14295_ ( .A1(_06521_ ), .A2(_06531_ ), .A3(_06100_ ), .ZN(_06994_ ) );
AOI21_X1 _14296_ ( .A(_06731_ ), .B1(_06993_ ), .B2(_06994_ ), .ZN(_06995_ ) );
OAI21_X1 _14297_ ( .A(_06538_ ), .B1(_06985_ ), .B2(_06995_ ), .ZN(_06996_ ) );
NAND3_X1 _14298_ ( .A1(_05925_ ), .A2(_06532_ ), .A3(_06495_ ), .ZN(_06997_ ) );
OR3_X1 _14299_ ( .A1(_06946_ ), .A2(_04668_ ), .A3(_05656_ ), .ZN(_06998_ ) );
NAND3_X1 _14300_ ( .A1(_06023_ ), .A2(_06947_ ), .A3(_06998_ ), .ZN(_06999_ ) );
OAI211_X1 _14301_ ( .A(_06313_ ), .B(_06314_ ), .C1(_04940_ ), .C2(_04939_ ), .ZN(_07000_ ) );
AOI21_X1 _14302_ ( .A(_04941_ ), .B1(_07000_ ), .B2(_06316_ ), .ZN(_07001_ ) );
NOR2_X1 _14303_ ( .A1(_07001_ ), .A2(_06186_ ), .ZN(_07002_ ) );
OAI21_X1 _14304_ ( .A(_04427_ ), .B1(_06071_ ), .B2(_04938_ ), .ZN(_07003_ ) );
OAI211_X1 _14305_ ( .A(_06997_ ), .B(_06999_ ), .C1(_07002_ ), .C2(_07003_ ), .ZN(_07004_ ) );
AOI21_X1 _14306_ ( .A(_07004_ ), .B1(_05306_ ), .B2(_06015_ ), .ZN(_07005_ ) );
AOI21_X1 _14307_ ( .A(_06014_ ), .B1(_06996_ ), .B2(_07005_ ), .ZN(_07006_ ) );
NOR2_X1 _14308_ ( .A1(_06974_ ), .A2(_06012_ ), .ZN(_07007_ ) );
AND2_X1 _14309_ ( .A1(_05309_ ), .A2(_05039_ ), .ZN(_07008_ ) );
NAND3_X1 _14310_ ( .A1(_05970_ ), .A2(\EXU.ls_rdata_i [6] ), .A3(_05971_ ), .ZN(_07009_ ) );
OAI21_X1 _14311_ ( .A(_07009_ ), .B1(_06763_ ), .B2(_04347_ ), .ZN(_07010_ ) );
NOR4_X1 _14312_ ( .A1(_07006_ ), .A2(_07007_ ), .A3(_07008_ ), .A4(_07010_ ), .ZN(_07011_ ) );
OAI21_X1 _14313_ ( .A(_06979_ ), .B1(_07011_ ), .B2(_06106_ ), .ZN(_07012_ ) );
NAND2_X1 _14314_ ( .A1(_07012_ ), .A2(_06610_ ), .ZN(_07013_ ) );
OAI211_X1 _14315_ ( .A(_06109_ ), .B(_05290_ ), .C1(_06976_ ), .C2(_06978_ ), .ZN(_07014_ ) );
AOI21_X1 _14316_ ( .A(_06563_ ), .B1(_07013_ ), .B2(_07014_ ), .ZN(_07015_ ) );
MUX2_X1 _14317_ ( .A(\EXU.xrd_o [6] ), .B(_07015_ ), .S(_06924_ ), .Z(_00259_ ) );
NAND4_X1 _14318_ ( .A1(_05831_ ), .A2(_05832_ ), .A3(\EXU.mtvec_i [5] ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_07016_ ) );
AOI22_X1 _14319_ ( .A1(_07016_ ), .A2(_05835_ ), .B1(_05836_ ), .B2(_05837_ ), .ZN(_07017_ ) );
AND3_X1 _14320_ ( .A1(_05837_ ), .A2(\EXU.mcause_i [5] ), .A3(_05839_ ), .ZN(_07018_ ) );
OAI21_X1 _14321_ ( .A(_05830_ ), .B1(_07017_ ), .B2(_07018_ ), .ZN(_07019_ ) );
NAND3_X1 _14322_ ( .A1(_06204_ ), .A2(_06208_ ), .A3(\EXU.mepc_i [5] ), .ZN(_07020_ ) );
NAND3_X1 _14323_ ( .A1(_06206_ ), .A2(\EXU.mstatus_i [5] ), .A3(_05989_ ), .ZN(_07021_ ) );
AND3_X1 _14324_ ( .A1(_07019_ ), .A2(_07020_ ), .A3(_07021_ ), .ZN(_07022_ ) );
NAND4_X1 _14325_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_26_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_07023_ ) );
AOI22_X1 _14326_ ( .A1(_07022_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_26_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_05557_ ), .B2(_07023_ ), .ZN(_07024_ ) );
NAND3_X1 _14327_ ( .A1(_06123_ ), .A2(\EXU.pc_i [5] ), .A3(_04348_ ), .ZN(_07025_ ) );
OAI21_X1 _14328_ ( .A(_07025_ ), .B1(_05006_ ), .B2(_06002_ ), .ZN(_07026_ ) );
OR2_X1 _14329_ ( .A1(_07024_ ), .A2(_07026_ ), .ZN(_07027_ ) );
NOR2_X1 _14330_ ( .A1(_06040_ ), .A2(\EXU.r1_i [5] ), .ZN(_07028_ ) );
NOR3_X1 _14331_ ( .A1(_06527_ ), .A2(\EXU.r1_i [6] ), .A3(_06050_ ), .ZN(_07029_ ) );
NOR2_X1 _14332_ ( .A1(_07028_ ), .A2(_07029_ ), .ZN(_07030_ ) );
MUX2_X1 _14333_ ( .A(_06937_ ), .B(_07030_ ), .S(_06144_ ), .Z(_07031_ ) );
MUX2_X1 _14334_ ( .A(_06860_ ), .B(_07031_ ), .S(_06526_ ), .Z(_07032_ ) );
NAND2_X1 _14335_ ( .A1(_07032_ ), .A2(_06532_ ), .ZN(_07033_ ) );
NAND2_X1 _14336_ ( .A1(_06580_ ), .A2(_06100_ ), .ZN(_07034_ ) );
AOI21_X1 _14337_ ( .A(_06731_ ), .B1(_07033_ ), .B2(_07034_ ), .ZN(_07035_ ) );
NAND3_X1 _14338_ ( .A1(_06025_ ), .A2(_06027_ ), .A3(_06550_ ), .ZN(_07036_ ) );
OAI21_X1 _14339_ ( .A(_07036_ ), .B1(_06062_ ), .B2(_06361_ ), .ZN(_07037_ ) );
OAI21_X1 _14340_ ( .A(_06538_ ), .B1(_07035_ ), .B2(_07037_ ), .ZN(_07038_ ) );
OR3_X1 _14341_ ( .A1(_06098_ ), .A2(_06081_ ), .A3(_06542_ ), .ZN(_07039_ ) );
AOI21_X1 _14342_ ( .A(_05654_ ), .B1(_05652_ ), .B2(_04671_ ), .ZN(_07040_ ) );
XNOR2_X1 _14343_ ( .A(_07040_ ), .B(_04670_ ), .ZN(_07041_ ) );
NAND3_X1 _14344_ ( .A1(_05638_ ), .A2(_05583_ ), .A3(_07041_ ), .ZN(_07042_ ) );
NAND3_X1 _14345_ ( .A1(_04943_ ), .A2(\EXU.r1_i [5] ), .A3(_04945_ ), .ZN(_07043_ ) );
AND3_X1 _14346_ ( .A1(_05572_ ), .A2(_05630_ ), .A3(_07043_ ), .ZN(_07044_ ) );
OAI22_X1 _14347_ ( .A1(_07044_ ), .A2(_05555_ ), .B1(\EXU.r1_i [5] ), .B2(_04948_ ), .ZN(_07045_ ) );
MUX2_X1 _14348_ ( .A(_04946_ ), .B(_07045_ ), .S(_06071_ ), .Z(_07046_ ) );
NAND3_X1 _14349_ ( .A1(_07039_ ), .A2(_07042_ ), .A3(_07046_ ), .ZN(_07047_ ) );
AOI21_X1 _14350_ ( .A(_07047_ ), .B1(_05313_ ), .B2(_05850_ ), .ZN(_07048_ ) );
AOI21_X1 _14351_ ( .A(_05849_ ), .B1(_07038_ ), .B2(_07048_ ), .ZN(_07049_ ) );
AOI22_X1 _14352_ ( .A1(_06006_ ), .A2(\EXU.ls_rdata_i [5] ), .B1(_06009_ ), .B2(\EXU.imm_i [5] ), .ZN(_07050_ ) );
OAI221_X1 _14353_ ( .A(_07050_ ), .B1(_05037_ ), .B2(_05318_ ), .C1(_07022_ ), .C2(_06011_ ), .ZN(_07051_ ) );
OR2_X1 _14354_ ( .A1(_07049_ ), .A2(_07051_ ), .ZN(_07052_ ) );
MUX2_X1 _14355_ ( .A(_07027_ ), .B(_07052_ ), .S(_05822_ ), .Z(_07053_ ) );
NAND2_X1 _14356_ ( .A1(_07053_ ), .A2(_06610_ ), .ZN(_07054_ ) );
BUF_X4 _14357_ ( .A(_04376_ ), .Z(_07055_ ) );
NAND3_X1 _14358_ ( .A1(_07055_ ), .A2(_05977_ ), .A3(_07027_ ), .ZN(_07056_ ) );
AOI21_X1 _14359_ ( .A(_06563_ ), .B1(_07054_ ), .B2(_07056_ ), .ZN(_07057_ ) );
MUX2_X1 _14360_ ( .A(\EXU.xrd_o [5] ), .B(_07057_ ), .S(_06924_ ), .Z(_00260_ ) );
BUF_X4 _14361_ ( .A(_04395_ ), .Z(_07058_ ) );
NAND4_X1 _14362_ ( .A1(_05831_ ), .A2(_05832_ ), .A3(\EXU.mtvec_i [4] ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_07059_ ) );
AOI22_X1 _14363_ ( .A1(_07059_ ), .A2(_05835_ ), .B1(_05836_ ), .B2(_05837_ ), .ZN(_07060_ ) );
AND3_X1 _14364_ ( .A1(_05837_ ), .A2(\EXU.mcause_i [4] ), .A3(_05839_ ), .ZN(_07061_ ) );
OAI21_X1 _14365_ ( .A(_05830_ ), .B1(_07060_ ), .B2(_07061_ ), .ZN(_07062_ ) );
NAND3_X1 _14366_ ( .A1(_06204_ ), .A2(_06208_ ), .A3(\EXU.mepc_i [4] ), .ZN(_07063_ ) );
NAND3_X1 _14367_ ( .A1(_06206_ ), .A2(\EXU.mstatus_i [4] ), .A3(_05989_ ), .ZN(_07064_ ) );
AND3_X1 _14368_ ( .A1(_07062_ ), .A2(_07063_ ), .A3(_07064_ ), .ZN(_07065_ ) );
NAND4_X1 _14369_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_27_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_07066_ ) );
AOI22_X1 _14370_ ( .A1(_07065_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_27_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .B1(_05557_ ), .B2(_07066_ ), .ZN(_07067_ ) );
NAND3_X1 _14371_ ( .A1(_06123_ ), .A2(\EXU.pc_i [4] ), .A3(_04348_ ), .ZN(_07068_ ) );
OAI21_X1 _14372_ ( .A(_07068_ ), .B1(_04955_ ), .B2(_06001_ ), .ZN(_07069_ ) );
OR2_X1 _14373_ ( .A1(_07067_ ), .A2(_07069_ ), .ZN(_07070_ ) );
OAI211_X1 _14374_ ( .A(_06027_ ), .B(_06549_ ), .C1(_06236_ ), .C2(_06152_ ), .ZN(_07071_ ) );
OAI21_X1 _14375_ ( .A(_07071_ ), .B1(_06180_ ), .B2(_06091_ ), .ZN(_07072_ ) );
NAND2_X1 _14376_ ( .A1(_06635_ ), .A2(_06100_ ), .ZN(_07073_ ) );
OR3_X1 _14377_ ( .A1(_06046_ ), .A2(\EXU.r1_i [5] ), .A3(_06050_ ), .ZN(_07074_ ) );
OAI21_X1 _14378_ ( .A(_04955_ ), .B1(_06046_ ), .B2(_06050_ ), .ZN(_07075_ ) );
NAND2_X1 _14379_ ( .A1(_07074_ ), .A2(_07075_ ), .ZN(_07076_ ) );
MUX2_X2 _14380_ ( .A(_07076_ ), .B(_06988_ ), .S(_05878_ ), .Z(_07077_ ) );
NOR2_X1 _14381_ ( .A1(_07077_ ), .A2(_06289_ ), .ZN(_07078_ ) );
AND3_X1 _14382_ ( .A1(_06888_ ), .A2(_06889_ ), .A3(_06289_ ), .ZN(_07079_ ) );
OAI21_X1 _14383_ ( .A(_06532_ ), .B1(_07078_ ), .B2(_07079_ ), .ZN(_07080_ ) );
AOI21_X1 _14384_ ( .A(_06731_ ), .B1(_07073_ ), .B2(_07080_ ), .ZN(_07081_ ) );
OAI21_X1 _14385_ ( .A(_06538_ ), .B1(_07072_ ), .B2(_07081_ ), .ZN(_07082_ ) );
XNOR2_X1 _14386_ ( .A(_05651_ ), .B(_04671_ ), .ZN(_07083_ ) );
AND3_X1 _14387_ ( .A1(_05638_ ), .A2(_05583_ ), .A3(_07083_ ), .ZN(_07084_ ) );
NAND3_X1 _14388_ ( .A1(_04950_ ), .A2(\EXU.r1_i [4] ), .A3(_04952_ ), .ZN(_07085_ ) );
NAND3_X1 _14389_ ( .A1(_05572_ ), .A2(_05630_ ), .A3(_07085_ ), .ZN(_07086_ ) );
AOI21_X1 _14390_ ( .A(_04956_ ), .B1(_07086_ ), .B2(_05556_ ), .ZN(_07087_ ) );
MUX2_X1 _14391_ ( .A(_04953_ ), .B(_07087_ ), .S(_05635_ ), .Z(_07088_ ) );
NOR3_X1 _14392_ ( .A1(_06133_ ), .A2(_06099_ ), .A3(_06542_ ), .ZN(_07089_ ) );
OR3_X1 _14393_ ( .A1(_07084_ ), .A2(_07088_ ), .A3(_07089_ ), .ZN(_07090_ ) );
AOI21_X1 _14394_ ( .A(_07090_ ), .B1(_05329_ ), .B2(_05585_ ), .ZN(_07091_ ) );
AOI21_X1 _14395_ ( .A(_05535_ ), .B1(_07082_ ), .B2(_07091_ ), .ZN(_07092_ ) );
NOR2_X1 _14396_ ( .A1(_07065_ ), .A2(_06011_ ), .ZN(_07093_ ) );
NAND3_X1 _14397_ ( .A1(_05817_ ), .A2(_05531_ ), .A3(\EXU.imm_i [4] ), .ZN(_07094_ ) );
INV_X1 _14398_ ( .A(\EXU.ls_rdata_i [4] ), .ZN(_07095_ ) );
OAI221_X1 _14399_ ( .A(_07094_ ), .B1(_04414_ ), .B2(_07095_ ), .C1(_05037_ ), .C2(_05324_ ), .ZN(_07096_ ) );
OR3_X1 _14400_ ( .A1(_07092_ ), .A2(_07093_ ), .A3(_07096_ ), .ZN(_07097_ ) );
BUF_X4 _14401_ ( .A(_05821_ ), .Z(_07098_ ) );
MUX2_X1 _14402_ ( .A(_07070_ ), .B(_07097_ ), .S(_07098_ ), .Z(_07099_ ) );
NAND2_X1 _14403_ ( .A1(_07099_ ), .A2(_06610_ ), .ZN(_07100_ ) );
NAND3_X1 _14404_ ( .A1(_07055_ ), .A2(_05977_ ), .A3(_07070_ ), .ZN(_07101_ ) );
AOI21_X1 _14405_ ( .A(_07058_ ), .B1(_07100_ ), .B2(_07101_ ), .ZN(_07102_ ) );
MUX2_X1 _14406_ ( .A(\EXU.xrd_o [4] ), .B(_07102_ ), .S(_06924_ ), .Z(_00261_ ) );
NAND4_X1 _14407_ ( .A1(_06208_ ), .A2(_05987_ ), .A3(\EXU.mtvec_i [3] ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_07103_ ) );
AOI22_X1 _14408_ ( .A1(_07103_ ), .A2(_05835_ ), .B1(_06204_ ), .B2(_06203_ ), .ZN(_07104_ ) );
AND3_X1 _14409_ ( .A1(_06203_ ), .A2(\EXU.mcause_i [3] ), .A3(_06204_ ), .ZN(_07105_ ) );
OAI21_X1 _14410_ ( .A(_05830_ ), .B1(_07104_ ), .B2(_07105_ ), .ZN(_07106_ ) );
AOI22_X1 _14411_ ( .A1(_05516_ ), .A2(\EXU.mstatus_i [3] ), .B1(_05518_ ), .B2(\EXU.mepc_i [3] ), .ZN(_07107_ ) );
NAND2_X1 _14412_ ( .A1(_07106_ ), .A2(_07107_ ), .ZN(_07108_ ) );
AND4_X1 _14413_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_07109_ ) );
OAI22_X1 _14414_ ( .A1(_07108_ ), .A2(_04882_ ), .B1(_05525_ ), .B2(_07109_ ), .ZN(_07110_ ) );
NAND3_X1 _14415_ ( .A1(_05045_ ), .A2(\EXU.pc_i [3] ), .A3(_05999_ ), .ZN(_07111_ ) );
NAND3_X1 _14416_ ( .A1(_04715_ ), .A2(_04710_ ), .A3(\EXU.r1_i [3] ), .ZN(_07112_ ) );
NAND3_X1 _14417_ ( .A1(_07110_ ), .A2(_07111_ ), .A3(_07112_ ), .ZN(_07113_ ) );
NOR2_X1 _14418_ ( .A1(_06738_ ), .A2(_06356_ ), .ZN(_07114_ ) );
NAND2_X1 _14419_ ( .A1(_06938_ ), .A2(_06289_ ), .ZN(_07115_ ) );
OAI21_X1 _14420_ ( .A(_06383_ ), .B1(_07028_ ), .B2(_07029_ ), .ZN(_07116_ ) );
OR3_X1 _14421_ ( .A1(_06527_ ), .A2(_04955_ ), .A3(_06528_ ), .ZN(_07117_ ) );
OAI21_X1 _14422_ ( .A(\EXU.r1_i [3] ), .B1(_06527_ ), .B2(_06528_ ), .ZN(_07118_ ) );
NAND2_X1 _14423_ ( .A1(_07117_ ), .A2(_07118_ ), .ZN(_07119_ ) );
OAI211_X1 _14424_ ( .A(_07116_ ), .B(_05881_ ), .C1(_06383_ ), .C2(_07119_ ), .ZN(_07120_ ) );
AOI21_X1 _14425_ ( .A(_06081_ ), .B1(_07115_ ), .B2(_07120_ ), .ZN(_07121_ ) );
OAI21_X1 _14426_ ( .A(_06091_ ), .B1(_07114_ ), .B2(_07121_ ), .ZN(_07122_ ) );
NAND3_X1 _14427_ ( .A1(_06236_ ), .A2(_06550_ ), .A3(_06027_ ), .ZN(_07123_ ) );
OAI211_X1 _14428_ ( .A(_07122_ ), .B(_07123_ ), .C1(_06234_ ), .C2(_06091_ ), .ZN(_07124_ ) );
NAND2_X1 _14429_ ( .A1(_07124_ ), .A2(_06538_ ), .ZN(_07125_ ) );
AOI21_X1 _14430_ ( .A(_05574_ ), .B1(\EXU.r1_i [3] ), .B2(_05757_ ), .ZN(_07126_ ) );
OAI22_X1 _14431_ ( .A1(_07126_ ), .A2(_05555_ ), .B1(\EXU.r1_i [3] ), .B2(_05757_ ), .ZN(_07127_ ) );
MUX2_X1 _14432_ ( .A(_04884_ ), .B(_07127_ ), .S(_05635_ ), .Z(_07128_ ) );
NAND2_X1 _14433_ ( .A1(_06251_ ), .A2(_06495_ ), .ZN(_07129_ ) );
NAND2_X1 _14434_ ( .A1(_07128_ ), .A2(_07129_ ), .ZN(_07130_ ) );
AOI21_X1 _14435_ ( .A(_05643_ ), .B1(_05644_ ), .B2(_05645_ ), .ZN(_07131_ ) );
OR3_X1 _14436_ ( .A1(_07131_ ), .A2(_05642_ ), .A3(_05647_ ), .ZN(_07132_ ) );
OAI21_X1 _14437_ ( .A(_05642_ ), .B1(_07131_ ), .B2(_05647_ ), .ZN(_07133_ ) );
AOI21_X1 _14438_ ( .A(_05640_ ), .B1(_07132_ ), .B2(_07133_ ), .ZN(_07134_ ) );
OR2_X1 _14439_ ( .A1(_07130_ ), .A2(_07134_ ), .ZN(_07135_ ) );
AOI21_X1 _14440_ ( .A(_07135_ ), .B1(_05338_ ), .B2(_05585_ ), .ZN(_07136_ ) );
AOI21_X1 _14441_ ( .A(_05535_ ), .B1(_07125_ ), .B2(_07136_ ), .ZN(_07137_ ) );
AOI21_X1 _14442_ ( .A(_06011_ ), .B1(_07106_ ), .B2(_07107_ ), .ZN(_07138_ ) );
NAND3_X1 _14443_ ( .A1(_05817_ ), .A2(_05531_ ), .A3(\EXU.imm_i [3] ), .ZN(_07139_ ) );
INV_X1 _14444_ ( .A(\EXU.ls_rdata_i [3] ), .ZN(_07140_ ) );
OAI221_X1 _14445_ ( .A(_07139_ ), .B1(_04414_ ), .B2(_07140_ ), .C1(_05037_ ), .C2(_05334_ ), .ZN(_07141_ ) );
OR3_X1 _14446_ ( .A1(_07137_ ), .A2(_07138_ ), .A3(_07141_ ), .ZN(_07142_ ) );
MUX2_X1 _14447_ ( .A(_07113_ ), .B(_07142_ ), .S(_07098_ ), .Z(_07143_ ) );
NAND2_X1 _14448_ ( .A1(_07143_ ), .A2(_06610_ ), .ZN(_07144_ ) );
OAI21_X1 _14449_ ( .A(_07055_ ), .B1(_05103_ ), .B2(_07113_ ), .ZN(_07145_ ) );
AOI21_X1 _14450_ ( .A(_07058_ ), .B1(_07144_ ), .B2(_07145_ ), .ZN(_07146_ ) );
MUX2_X1 _14451_ ( .A(\EXU.xrd_o [3] ), .B(_07146_ ), .S(_06924_ ), .Z(_00262_ ) );
AOI22_X1 _14452_ ( .A1(_05516_ ), .A2(\EXU.mstatus_i [2] ), .B1(_04336_ ), .B2(\EXU.mcause_i [2] ), .ZN(_07147_ ) );
AOI22_X1 _14453_ ( .A1(_04353_ ), .A2(\EXU.mtvec_i [2] ), .B1(_05518_ ), .B2(\EXU.mepc_i [2] ), .ZN(_07148_ ) );
NAND2_X1 _14454_ ( .A1(_07147_ ), .A2(_07148_ ), .ZN(_07149_ ) );
AND4_X1 _14455_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_B_$_MUX__Y_A ), .A4(fanout_net_10 ), .ZN(_07150_ ) );
OAI22_X1 _14456_ ( .A1(_07149_ ), .A2(_04458_ ), .B1(_05525_ ), .B2(_07150_ ), .ZN(_07151_ ) );
AOI22_X1 _14457_ ( .A1(_04359_ ), .A2(\EXU.pc_i [2] ), .B1(\EXU.r1_i [2] ), .B2(_05528_ ), .ZN(_07152_ ) );
NAND2_X1 _14458_ ( .A1(_07151_ ), .A2(_07152_ ), .ZN(_07153_ ) );
NAND3_X1 _14459_ ( .A1(_06292_ ), .A2(_06027_ ), .A3(_06550_ ), .ZN(_07154_ ) );
OAI21_X1 _14460_ ( .A(_07154_ ), .B1(_06310_ ), .B2(_06361_ ), .ZN(_07155_ ) );
NAND2_X1 _14461_ ( .A1(_06795_ ), .A2(_06081_ ), .ZN(_07156_ ) );
NAND2_X1 _14462_ ( .A1(_07076_ ), .A2(_06383_ ), .ZN(_07157_ ) );
OR3_X1 _14463_ ( .A1(_06527_ ), .A2(_05649_ ), .A3(_06528_ ), .ZN(_07158_ ) );
OAI21_X1 _14464_ ( .A(\EXU.r1_i [2] ), .B1(_06527_ ), .B2(_06528_ ), .ZN(_07159_ ) );
NAND2_X1 _14465_ ( .A1(_07158_ ), .A2(_07159_ ), .ZN(_07160_ ) );
OAI211_X1 _14466_ ( .A(_07157_ ), .B(_06526_ ), .C1(_06383_ ), .C2(_07160_ ), .ZN(_07161_ ) );
OAI211_X1 _14467_ ( .A(_07161_ ), .B(_06356_ ), .C1(_06526_ ), .C2(_06991_ ), .ZN(_07162_ ) );
AND3_X1 _14468_ ( .A1(_07156_ ), .A2(_06091_ ), .A3(_07162_ ), .ZN(_07163_ ) );
OAI21_X1 _14469_ ( .A(_06538_ ), .B1(_07155_ ), .B2(_07163_ ), .ZN(_07164_ ) );
AND3_X1 _14470_ ( .A1(_05644_ ), .A2(_05645_ ), .A3(_05643_ ), .ZN(_07165_ ) );
NOR3_X1 _14471_ ( .A1(_05640_ ), .A2(_07131_ ), .A3(_07165_ ), .ZN(_07166_ ) );
NAND3_X1 _14472_ ( .A1(_04889_ ), .A2(\EXU.r1_i [2] ), .A3(_04890_ ), .ZN(_07167_ ) );
NAND3_X1 _14473_ ( .A1(_05572_ ), .A2(_05630_ ), .A3(_07167_ ), .ZN(_07168_ ) );
AOI21_X1 _14474_ ( .A(_04894_ ), .B1(_07168_ ), .B2(_05556_ ), .ZN(_07169_ ) );
MUX2_X1 _14475_ ( .A(_04891_ ), .B(_07169_ ), .S(_05635_ ), .Z(_07170_ ) );
NOR4_X1 _14476_ ( .A1(_05923_ ), .A2(_06099_ ), .A3(_06289_ ), .A4(_06542_ ), .ZN(_07171_ ) );
OR3_X1 _14477_ ( .A1(_07166_ ), .A2(_07170_ ), .A3(_07171_ ), .ZN(_07172_ ) );
AOI21_X1 _14478_ ( .A(_07172_ ), .B1(_05343_ ), .B2(_05850_ ), .ZN(_07173_ ) );
AOI21_X1 _14479_ ( .A(_05849_ ), .B1(_07164_ ), .B2(_07173_ ), .ZN(_07174_ ) );
NAND2_X1 _14480_ ( .A1(_07149_ ), .A2(_06516_ ), .ZN(_07175_ ) );
OAI211_X1 _14481_ ( .A(_04415_ ), .B(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_B_$_MUX__Y_B ), .C1(_05968_ ), .C2(_05035_ ), .ZN(_07176_ ) );
NAND3_X1 _14482_ ( .A1(_05967_ ), .A2(_05968_ ), .A3(\EXU.imm_i [2] ), .ZN(_07177_ ) );
NAND3_X1 _14483_ ( .A1(_05970_ ), .A2(\EXU.ls_rdata_i [2] ), .A3(_05971_ ), .ZN(_07178_ ) );
NAND4_X1 _14484_ ( .A1(_07175_ ), .A2(_07176_ ), .A3(_07177_ ), .A4(_07178_ ), .ZN(_07179_ ) );
OR2_X1 _14485_ ( .A1(_07174_ ), .A2(_07179_ ), .ZN(_07180_ ) );
MUX2_X1 _14486_ ( .A(_07153_ ), .B(_07180_ ), .S(_07098_ ), .Z(_07181_ ) );
BUF_X4 _14487_ ( .A(_05824_ ), .Z(_07182_ ) );
NAND2_X1 _14488_ ( .A1(_07181_ ), .A2(_07182_ ), .ZN(_07183_ ) );
NAND3_X1 _14489_ ( .A1(_07055_ ), .A2(_05264_ ), .A3(_07153_ ), .ZN(_07184_ ) );
AOI21_X1 _14490_ ( .A(_07058_ ), .B1(_07183_ ), .B2(_07184_ ), .ZN(_07185_ ) );
MUX2_X1 _14491_ ( .A(\EXU.xrd_o [2] ), .B(_07185_ ), .S(_06924_ ), .Z(_00263_ ) );
NAND4_X1 _14492_ ( .A1(_05984_ ), .A2(_05832_ ), .A3(\EXU.mtvec_i [28] ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_07186_ ) );
AOI22_X1 _14493_ ( .A1(_07186_ ), .A2(_05835_ ), .B1(_05836_ ), .B2(_05837_ ), .ZN(_07187_ ) );
AND3_X1 _14494_ ( .A1(_04334_ ), .A2(\EXU.mcause_i [28] ), .A3(_05839_ ), .ZN(_07188_ ) );
OAI21_X1 _14495_ ( .A(_05830_ ), .B1(_07187_ ), .B2(_07188_ ), .ZN(_07189_ ) );
AOI22_X1 _14496_ ( .A1(_05516_ ), .A2(\EXU.mstatus_i [28] ), .B1(_05518_ ), .B2(\EXU.mepc_i [28] ), .ZN(_07190_ ) );
NAND2_X1 _14497_ ( .A1(_07189_ ), .A2(_07190_ ), .ZN(_07191_ ) );
AND4_X1 _14498_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_3_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_07192_ ) );
OAI22_X1 _14499_ ( .A1(_07191_ ), .A2(_06723_ ), .B1(_05525_ ), .B2(_07192_ ), .ZN(_07193_ ) );
AOI22_X1 _14500_ ( .A1(_04359_ ), .A2(\EXU.pc_i [28] ), .B1(\EXU.r1_i [28] ), .B2(_04716_ ), .ZN(_07194_ ) );
NAND2_X1 _14501_ ( .A1(_07193_ ), .A2(_07194_ ), .ZN(_07195_ ) );
NAND2_X1 _14502_ ( .A1(_05345_ ), .A2(_05850_ ), .ZN(_07196_ ) );
NOR2_X1 _14503_ ( .A1(_06699_ ), .A2(_05641_ ), .ZN(_07197_ ) );
NAND3_X1 _14504_ ( .A1(_06697_ ), .A2(_06696_ ), .A3(_06698_ ), .ZN(_07198_ ) );
NAND2_X1 _14505_ ( .A1(_07197_ ), .A2(_07198_ ), .ZN(_07199_ ) );
AOI21_X1 _14506_ ( .A(_05855_ ), .B1(_06642_ ), .B2(_05868_ ), .ZN(_07200_ ) );
NOR4_X1 _14507_ ( .A1(_07200_ ), .A2(_05591_ ), .A3(_05626_ ), .A4(_05870_ ), .ZN(_07201_ ) );
NOR3_X1 _14508_ ( .A1(_06639_ ), .A2(_06060_ ), .A3(_06357_ ), .ZN(_07202_ ) );
AND2_X1 _14509_ ( .A1(_07202_ ), .A2(_05807_ ), .ZN(_07203_ ) );
OAI21_X1 _14510_ ( .A(_06066_ ), .B1(_07201_ ), .B2(_07203_ ), .ZN(_07204_ ) );
OAI211_X1 _14511_ ( .A(_05887_ ), .B(_05888_ ), .C1(_04778_ ), .C2(_04776_ ), .ZN(_07205_ ) );
AOI21_X1 _14512_ ( .A(_04779_ ), .B1(_07205_ ), .B2(_05890_ ), .ZN(_07206_ ) );
AOI21_X1 _14513_ ( .A(_07206_ ), .B1(_04777_ ), .B2(_06186_ ), .ZN(_07207_ ) );
AOI21_X1 _14514_ ( .A(_05767_ ), .B1(_06652_ ), .B2(_06181_ ), .ZN(_07208_ ) );
NAND3_X1 _14515_ ( .A1(_06145_ ), .A2(_06099_ ), .A3(_06147_ ), .ZN(_07209_ ) );
NAND3_X1 _14516_ ( .A1(_05929_ ), .A2(_06144_ ), .A3(_05930_ ), .ZN(_07210_ ) );
OAI211_X1 _14517_ ( .A(_07210_ ), .B(_06030_ ), .C1(_05937_ ), .C2(_06414_ ), .ZN(_07211_ ) );
NAND2_X1 _14518_ ( .A1(_05928_ ), .A2(_04825_ ), .ZN(_07212_ ) );
OAI211_X1 _14519_ ( .A(_07212_ ), .B(_05877_ ), .C1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ), .C2(_05928_ ), .ZN(_07213_ ) );
OAI211_X1 _14520_ ( .A(_05940_ ), .B(_06049_ ), .C1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ), .C2(_05928_ ), .ZN(_07214_ ) );
AND2_X1 _14521_ ( .A1(_07213_ ), .A2(_07214_ ), .ZN(_07215_ ) );
OAI211_X1 _14522_ ( .A(_05880_ ), .B(_07211_ ), .C1(_07215_ ), .C2(_05881_ ), .ZN(_07216_ ) );
NAND3_X1 _14523_ ( .A1(_07209_ ), .A2(_07216_ ), .A3(_05807_ ), .ZN(_07217_ ) );
NAND2_X1 _14524_ ( .A1(_07208_ ), .A2(_07217_ ), .ZN(_07218_ ) );
AND4_X1 _14525_ ( .A1(_07199_ ), .A2(_07204_ ), .A3(_07207_ ), .A4(_07218_ ), .ZN(_07219_ ) );
AOI21_X1 _14526_ ( .A(_05535_ ), .B1(_07196_ ), .B2(_07219_ ), .ZN(_07220_ ) );
AND2_X1 _14527_ ( .A1(_05347_ ), .A2(_06500_ ), .ZN(_07221_ ) );
NAND2_X1 _14528_ ( .A1(_07191_ ), .A2(_05044_ ), .ZN(_07222_ ) );
NAND3_X1 _14529_ ( .A1(_05967_ ), .A2(_05968_ ), .A3(\EXU.imm_i [28] ), .ZN(_07223_ ) );
NAND3_X1 _14530_ ( .A1(_05970_ ), .A2(\EXU.ls_rdata_i [28] ), .A3(_05971_ ), .ZN(_07224_ ) );
NAND3_X1 _14531_ ( .A1(_07222_ ), .A2(_07223_ ), .A3(_07224_ ), .ZN(_07225_ ) );
OR3_X1 _14532_ ( .A1(_07220_ ), .A2(_07221_ ), .A3(_07225_ ), .ZN(_07226_ ) );
MUX2_X1 _14533_ ( .A(_07195_ ), .B(_07226_ ), .S(_07098_ ), .Z(_07227_ ) );
NAND2_X1 _14534_ ( .A1(_07227_ ), .A2(_07182_ ), .ZN(_07228_ ) );
NAND3_X1 _14535_ ( .A1(_07055_ ), .A2(_05264_ ), .A3(_07195_ ), .ZN(_07229_ ) );
AOI21_X1 _14536_ ( .A(_07058_ ), .B1(_07228_ ), .B2(_07229_ ), .ZN(_07230_ ) );
MUX2_X1 _14537_ ( .A(\EXU.xrd_o [28] ), .B(_07230_ ), .S(_06924_ ), .Z(_00264_ ) );
AOI22_X1 _14538_ ( .A1(_05516_ ), .A2(\EXU.mstatus_i [1] ), .B1(_04336_ ), .B2(\EXU.mcause_i [1] ), .ZN(_07231_ ) );
AOI22_X1 _14539_ ( .A1(_04353_ ), .A2(\EXU.mtvec_i [1] ), .B1(_05518_ ), .B2(\EXU.mepc_i [1] ), .ZN(_07232_ ) );
NAND2_X1 _14540_ ( .A1(_07231_ ), .A2(_07232_ ), .ZN(_07233_ ) );
AND4_X1 _14541_ ( .A1(fanout_net_6 ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_07234_ ) );
OAI22_X1 _14542_ ( .A1(_07233_ ), .A2(_04898_ ), .B1(_05525_ ), .B2(_07234_ ), .ZN(_07235_ ) );
AOI22_X1 _14543_ ( .A1(_05103_ ), .A2(\EXU.add_pc_4 [1] ), .B1(\EXU.r1_i [1] ), .B2(_05528_ ), .ZN(_07236_ ) );
NAND2_X1 _14544_ ( .A1(_07235_ ), .A2(_07236_ ), .ZN(_07237_ ) );
AND3_X1 _14545_ ( .A1(_06363_ ), .A2(_06027_ ), .A3(_06550_ ), .ZN(_07238_ ) );
AOI21_X1 _14546_ ( .A(_07238_ ), .B1(_06360_ ), .B2(_06731_ ), .ZN(_07239_ ) );
AND2_X1 _14547_ ( .A1(_06861_ ), .A2(_06100_ ), .ZN(_07240_ ) );
NAND2_X1 _14548_ ( .A1(_07031_ ), .A2(_06289_ ), .ZN(_07241_ ) );
OR3_X1 _14549_ ( .A1(_06527_ ), .A2(_04893_ ), .A3(_06528_ ), .ZN(_07242_ ) );
OAI211_X1 _14550_ ( .A(_07242_ ), .B(_06414_ ), .C1(_05000_ ), .C2(_06040_ ), .ZN(_07243_ ) );
OAI211_X1 _14551_ ( .A(_07243_ ), .B(_06526_ ), .C1(_06414_ ), .C2(_07119_ ), .ZN(_07244_ ) );
AOI21_X1 _14552_ ( .A(_06100_ ), .B1(_07241_ ), .B2(_07244_ ), .ZN(_07245_ ) );
OAI21_X1 _14553_ ( .A(_06361_ ), .B1(_07240_ ), .B2(_07245_ ), .ZN(_07246_ ) );
AOI21_X1 _14554_ ( .A(_05852_ ), .B1(_07239_ ), .B2(_07246_ ), .ZN(_07247_ ) );
NAND3_X1 _14555_ ( .A1(_04655_ ), .A2(_04911_ ), .A3(\EXU.r2_i [0] ), .ZN(_07248_ ) );
AND3_X1 _14556_ ( .A1(_06023_ ), .A2(_05644_ ), .A3(_07248_ ), .ZN(_07249_ ) );
AND3_X1 _14557_ ( .A1(_04900_ ), .A2(_05539_ ), .A3(_05537_ ), .ZN(_07250_ ) );
NAND3_X1 _14558_ ( .A1(_04897_ ), .A2(\EXU.r1_i [1] ), .A3(_04899_ ), .ZN(_07251_ ) );
AND3_X1 _14559_ ( .A1(_05887_ ), .A2(_05888_ ), .A3(_07251_ ), .ZN(_07252_ ) );
OAI22_X1 _14560_ ( .A1(_07252_ ), .A2(_05555_ ), .B1(\EXU.r1_i [1] ), .B2(_06383_ ), .ZN(_07253_ ) );
AOI21_X1 _14561_ ( .A(_07250_ ), .B1(_07253_ ), .B2(_06071_ ), .ZN(_07254_ ) );
AND4_X1 _14562_ ( .A1(_06532_ ), .A2(_06097_ ), .A3(_06526_ ), .A4(_06495_ ), .ZN(_07255_ ) );
NOR3_X1 _14563_ ( .A1(_07249_ ), .A2(_07254_ ), .A3(_07255_ ), .ZN(_07256_ ) );
OAI21_X1 _14564_ ( .A(_07256_ ), .B1(_05354_ ), .B2(_06787_ ), .ZN(_07257_ ) );
OAI21_X1 _14565_ ( .A(_06626_ ), .B1(_07247_ ), .B2(_07257_ ), .ZN(_07258_ ) );
NAND2_X1 _14566_ ( .A1(_07233_ ), .A2(_05045_ ), .ZN(_07259_ ) );
OAI211_X1 _14567_ ( .A(_04415_ ), .B(\EXU.add_pc_4 [1] ), .C1(_05968_ ), .C2(_05035_ ), .ZN(_07260_ ) );
AOI22_X1 _14568_ ( .A1(_06007_ ), .A2(\EXU.ls_rdata_i [1] ), .B1(_06009_ ), .B2(\EXU.imm_i [1] ), .ZN(_07261_ ) );
NAND4_X1 _14569_ ( .A1(_07258_ ), .A2(_07259_ ), .A3(_07260_ ), .A4(_07261_ ), .ZN(_07262_ ) );
MUX2_X1 _14570_ ( .A(_07237_ ), .B(_07262_ ), .S(_07098_ ), .Z(_07263_ ) );
NAND2_X1 _14571_ ( .A1(_07263_ ), .A2(_07182_ ), .ZN(_07264_ ) );
OAI21_X1 _14572_ ( .A(_07055_ ), .B1(_05103_ ), .B2(_07237_ ), .ZN(_07265_ ) );
AOI21_X1 _14573_ ( .A(_07058_ ), .B1(_07264_ ), .B2(_07265_ ), .ZN(_07266_ ) );
MUX2_X1 _14574_ ( .A(\EXU.xrd_o [1] ), .B(_07266_ ), .S(_06924_ ), .Z(_00265_ ) );
NAND4_X1 _14575_ ( .A1(_05832_ ), .A2(\EXU.dnpc_$_MUX__Y_31_B_$_MUX__B_Y_$_MUX__B_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_04345_ ), .ZN(_07267_ ) );
NOR2_X1 _14576_ ( .A1(_05980_ ), .A2(\EXU.dnpc_$_MUX__Y_31_B_$_MUX__B_Y_$_MUX__B_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07268_ ) );
AND3_X1 _14577_ ( .A1(_04352_ ), .A2(_05363_ ), .A3(_04349_ ), .ZN(_07269_ ) );
OR3_X1 _14578_ ( .A1(_07268_ ), .A2(_06201_ ), .A3(_07269_ ), .ZN(_07270_ ) );
OAI21_X1 _14579_ ( .A(_07267_ ), .B1(_07270_ ), .B2(_04355_ ), .ZN(_07271_ ) );
MUX2_X1 _14580_ ( .A(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_B_$_MUX__A_B ), .B(_07271_ ), .S(_05992_ ), .Z(_07272_ ) );
NAND4_X1 _14581_ ( .A1(_04911_ ), .A2(fanout_net_6 ), .A3(fanout_net_5 ), .A4(fanout_net_10 ), .ZN(_07273_ ) );
AOI22_X1 _14582_ ( .A1(_07272_ ), .A2(_04911_ ), .B1(_05995_ ), .B2(_07273_ ), .ZN(_07274_ ) );
NAND3_X1 _14583_ ( .A1(_06123_ ), .A2(\EXU.add_pc_4 [0] ), .A3(_05046_ ), .ZN(_07275_ ) );
OAI21_X1 _14584_ ( .A(_07275_ ), .B1(_04911_ ), .B2(_06002_ ), .ZN(_07276_ ) );
OR2_X1 _14585_ ( .A1(_07274_ ), .A2(_07276_ ), .ZN(_07277_ ) );
AOI21_X1 _14586_ ( .A(_05852_ ), .B1(_06425_ ), .B2(_06731_ ), .ZN(_07278_ ) );
MUX2_X1 _14587_ ( .A(\EXU.r1_i [0] ), .B(\EXU.r1_i [1] ), .S(_06040_ ), .Z(_07279_ ) );
OAI21_X1 _14588_ ( .A(_05881_ ), .B1(_07279_ ), .B2(_06383_ ), .ZN(_07280_ ) );
AND3_X1 _14589_ ( .A1(_07158_ ), .A2(_06383_ ), .A3(_07159_ ), .ZN(_07281_ ) );
OAI22_X1 _14590_ ( .A1(_07280_ ), .A2(_07281_ ), .B1(_07077_ ), .B2(_06526_ ), .ZN(_07282_ ) );
MUX2_X1 _14591_ ( .A(_07282_ ), .B(_06891_ ), .S(_06081_ ), .Z(_07283_ ) );
OAI21_X1 _14592_ ( .A(_07278_ ), .B1(_07283_ ), .B2(_06731_ ), .ZN(_07284_ ) );
NAND3_X1 _14593_ ( .A1(_05638_ ), .A2(_04658_ ), .A3(_05583_ ), .ZN(_07285_ ) );
OAI211_X1 _14594_ ( .A(_05572_ ), .B(_05630_ ), .C1(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_A ), .C2(_04909_ ), .ZN(_07286_ ) );
AOI21_X1 _14595_ ( .A(_04910_ ), .B1(_07286_ ), .B2(_05890_ ), .ZN(_07287_ ) );
AND4_X1 _14596_ ( .A1(_05747_ ), .A2(_06128_ ), .A3(_06495_ ), .A4(_05934_ ), .ZN(_07288_ ) );
AND2_X1 _14597_ ( .A1(_05634_ ), .A2(_04912_ ), .ZN(_07289_ ) );
NOR3_X1 _14598_ ( .A1(_07287_ ), .A2(_07288_ ), .A3(_07289_ ), .ZN(_07290_ ) );
OAI211_X1 _14599_ ( .A(_07285_ ), .B(_07290_ ), .C1(_06787_ ), .C2(_05361_ ), .ZN(_07291_ ) );
AND4_X1 _14600_ ( .A1(_06027_ ), .A2(_06549_ ), .A3(_06153_ ), .A4(_06152_ ), .ZN(_07292_ ) );
AOI211_X1 _14601_ ( .A(_07291_ ), .B(_07292_ ), .C1(_05031_ ), .C2(_05577_ ), .ZN(_07293_ ) );
AOI21_X1 _14602_ ( .A(_05534_ ), .B1(_07284_ ), .B2(_07293_ ), .ZN(_07294_ ) );
NOR2_X1 _14603_ ( .A1(_07272_ ), .A2(_05814_ ), .ZN(_07295_ ) );
AND2_X1 _14604_ ( .A1(_06500_ ), .A2(\EXU.add_pc_4 [0] ), .ZN(_07296_ ) );
NAND3_X1 _14605_ ( .A1(_04387_ ), .A2(\EXU.ls_rdata_i [0] ), .A3(_04388_ ), .ZN(_07297_ ) );
OAI21_X1 _14606_ ( .A(_07297_ ), .B1(_06763_ ), .B2(_04333_ ), .ZN(_07298_ ) );
OR4_X2 _14607_ ( .A1(_07294_ ), .A2(_07295_ ), .A3(_07296_ ), .A4(_07298_ ), .ZN(_07299_ ) );
MUX2_X2 _14608_ ( .A(_07277_ ), .B(_07299_ ), .S(_07098_ ), .Z(_07300_ ) );
NAND2_X1 _14609_ ( .A1(_07300_ ), .A2(_07182_ ), .ZN(_07301_ ) );
OAI21_X1 _14610_ ( .A(_06109_ ), .B1(_07277_ ), .B2(_05103_ ), .ZN(_07302_ ) );
AOI21_X1 _14611_ ( .A(_07058_ ), .B1(_07301_ ), .B2(_07302_ ), .ZN(_07303_ ) );
MUX2_X1 _14612_ ( .A(\EXU.xrd_o [0] ), .B(_07303_ ), .S(_06924_ ), .Z(_00266_ ) );
NAND4_X1 _14613_ ( .A1(_05984_ ), .A2(_05832_ ), .A3(\EXU.mtvec_i [27] ), .A4(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_07304_ ) );
AOI22_X1 _14614_ ( .A1(_07304_ ), .A2(_05835_ ), .B1(_05839_ ), .B2(_05837_ ), .ZN(_07305_ ) );
AND3_X1 _14615_ ( .A1(_04334_ ), .A2(\EXU.mcause_i [27] ), .A3(_05839_ ), .ZN(_07306_ ) );
OAI21_X1 _14616_ ( .A(_05829_ ), .B1(_07305_ ), .B2(_07306_ ), .ZN(_07307_ ) );
AOI22_X1 _14617_ ( .A1(_05516_ ), .A2(\EXU.mstatus_i [27] ), .B1(_05518_ ), .B2(\EXU.mepc_i [27] ), .ZN(_07308_ ) );
NAND2_X1 _14618_ ( .A1(_07307_ ), .A2(_07308_ ), .ZN(_07309_ ) );
INV_X1 _14619_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_4_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_07310_ ) );
AND4_X1 _14620_ ( .A1(\EXU.funct3_i [1] ), .A2(fanout_net_5 ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_4_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A4(fanout_net_10 ), .ZN(_07311_ ) );
OAI22_X1 _14621_ ( .A1(_07309_ ), .A2(_07310_ ), .B1(_05525_ ), .B2(_07311_ ), .ZN(_07312_ ) );
AOI22_X1 _14622_ ( .A1(_04359_ ), .A2(\EXU.pc_i [27] ), .B1(\EXU.r1_i [27] ), .B2(_04716_ ), .ZN(_07313_ ) );
NAND2_X1 _14623_ ( .A1(_07312_ ), .A2(_07313_ ), .ZN(_07314_ ) );
NAND2_X1 _14624_ ( .A1(_05370_ ), .A2(_05585_ ), .ZN(_07315_ ) );
INV_X1 _14625_ ( .A(_04677_ ), .ZN(_07316_ ) );
NAND2_X1 _14626_ ( .A1(_05706_ ), .A2(_04675_ ), .ZN(_07317_ ) );
AOI21_X1 _14627_ ( .A(_07316_ ), .B1(_07317_ ), .B2(_05710_ ), .ZN(_07318_ ) );
AOI21_X1 _14628_ ( .A(_07318_ ), .B1(\EXU.r1_i [26] ), .B2(_05714_ ), .ZN(_07319_ ) );
XNOR2_X1 _14629_ ( .A(_07319_ ), .B(_04676_ ), .ZN(_07320_ ) );
NAND2_X1 _14630_ ( .A1(_07320_ ), .A2(_06023_ ), .ZN(_07321_ ) );
NOR2_X1 _14631_ ( .A1(_06729_ ), .A2(_06181_ ), .ZN(_07322_ ) );
NOR3_X1 _14632_ ( .A1(_05855_ ), .A2(_06854_ ), .A3(_06236_ ), .ZN(_07323_ ) );
NOR4_X1 _14633_ ( .A1(_07323_ ), .A2(_05591_ ), .A3(_05626_ ), .A4(_05870_ ), .ZN(_07324_ ) );
OAI21_X1 _14634_ ( .A(_06066_ ), .B1(_07322_ ), .B2(_07324_ ), .ZN(_07325_ ) );
OAI21_X1 _14635_ ( .A(_05914_ ), .B1(_06743_ ), .B2(_06744_ ), .ZN(_07326_ ) );
AND2_X1 _14636_ ( .A1(_05775_ ), .A2(_05778_ ), .ZN(_07327_ ) );
MUX2_X1 _14637_ ( .A(_05796_ ), .B(_07327_ ), .S(_05755_ ), .Z(_07328_ ) );
MUX2_X1 _14638_ ( .A(_06257_ ), .B(_07328_ ), .S(_05747_ ), .Z(_07329_ ) );
OAI21_X1 _14639_ ( .A(_07326_ ), .B1(_07329_ ), .B2(_06181_ ), .ZN(_07330_ ) );
NAND2_X1 _14640_ ( .A1(_07330_ ), .A2(_05565_ ), .ZN(_07331_ ) );
AND4_X1 _14641_ ( .A1(_07310_ ), .A2(_05892_ ), .A3(_04798_ ), .A4(_04799_ ), .ZN(_07332_ ) );
OAI211_X1 _14642_ ( .A(_06313_ ), .B(_06314_ ), .C1(_04801_ ), .C2(_04800_ ), .ZN(_07333_ ) );
NAND2_X1 _14643_ ( .A1(_07333_ ), .A2(_06316_ ), .ZN(_07334_ ) );
AOI21_X1 _14644_ ( .A(_07332_ ), .B1(_07334_ ), .B2(_04802_ ), .ZN(_07335_ ) );
AND4_X1 _14645_ ( .A1(_07321_ ), .A2(_07325_ ), .A3(_07331_ ), .A4(_07335_ ), .ZN(_07336_ ) );
AOI21_X1 _14646_ ( .A(_05535_ ), .B1(_07315_ ), .B2(_07336_ ), .ZN(_07337_ ) );
AND2_X1 _14647_ ( .A1(_05373_ ), .A2(_06500_ ), .ZN(_07338_ ) );
NAND2_X1 _14648_ ( .A1(_07309_ ), .A2(_05044_ ), .ZN(_07339_ ) );
NAND3_X1 _14649_ ( .A1(_05967_ ), .A2(_05531_ ), .A3(\EXU.imm_i [27] ), .ZN(_07340_ ) );
NAND3_X1 _14650_ ( .A1(_05970_ ), .A2(\EXU.ls_rdata_i [27] ), .A3(_05971_ ), .ZN(_07341_ ) );
NAND3_X1 _14651_ ( .A1(_07339_ ), .A2(_07340_ ), .A3(_07341_ ), .ZN(_07342_ ) );
OR3_X1 _14652_ ( .A1(_07337_ ), .A2(_07338_ ), .A3(_07342_ ), .ZN(_07343_ ) );
MUX2_X1 _14653_ ( .A(_07314_ ), .B(_07343_ ), .S(_07098_ ), .Z(_07344_ ) );
NAND2_X1 _14654_ ( .A1(_07344_ ), .A2(_07182_ ), .ZN(_07345_ ) );
NAND3_X1 _14655_ ( .A1(_07055_ ), .A2(_05264_ ), .A3(_07314_ ), .ZN(_07346_ ) );
AOI21_X1 _14656_ ( .A(_07058_ ), .B1(_07345_ ), .B2(_07346_ ), .ZN(_07347_ ) );
MUX2_X1 _14657_ ( .A(\EXU.xrd_o [27] ), .B(_07347_ ), .S(_04399_ ), .Z(_00267_ ) );
AOI22_X1 _14658_ ( .A1(_04355_ ), .A2(\EXU.mstatus_i [26] ), .B1(_04336_ ), .B2(\EXU.mcause_i [26] ), .ZN(_07348_ ) );
AOI22_X1 _14659_ ( .A1(_04353_ ), .A2(\EXU.mtvec_i [26] ), .B1(_05518_ ), .B2(\EXU.mepc_i [26] ), .ZN(_07349_ ) );
NAND2_X1 _14660_ ( .A1(_07348_ ), .A2(_07349_ ), .ZN(_07350_ ) );
NAND3_X1 _14661_ ( .A1(_07350_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_5_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A3(_05559_ ), .ZN(_07351_ ) );
AND3_X1 _14662_ ( .A1(_07348_ ), .A2(_07349_ ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_5_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_07352_ ) );
OAI221_X1 _14663_ ( .A(_07351_ ), .B1(_04808_ ), .B2(_06001_ ), .C1(_07352_ ), .C2(_05995_ ), .ZN(_07353_ ) );
AND3_X1 _14664_ ( .A1(_06516_ ), .A2(\EXU.pc_i [26] ), .A3(_05046_ ), .ZN(_07354_ ) );
OR2_X1 _14665_ ( .A1(_07353_ ), .A2(_07354_ ), .ZN(_07355_ ) );
NAND2_X1 _14666_ ( .A1(_05382_ ), .A2(_05585_ ), .ZN(_07356_ ) );
NOR2_X1 _14667_ ( .A1(_07318_ ), .A2(_05641_ ), .ZN(_07357_ ) );
NAND3_X1 _14668_ ( .A1(_07317_ ), .A2(_07316_ ), .A3(_05710_ ), .ZN(_07358_ ) );
NAND2_X1 _14669_ ( .A1(_07357_ ), .A2(_07358_ ), .ZN(_07359_ ) );
AND2_X1 _14670_ ( .A1(_06806_ ), .A2(_05807_ ), .ZN(_07360_ ) );
AOI21_X1 _14671_ ( .A(_05855_ ), .B1(_06798_ ), .B2(_05868_ ), .ZN(_07361_ ) );
NOR4_X1 _14672_ ( .A1(_07361_ ), .A2(_05591_ ), .A3(_05626_ ), .A4(_05870_ ), .ZN(_07362_ ) );
OAI21_X1 _14673_ ( .A(_06065_ ), .B1(_07360_ ), .B2(_07362_ ), .ZN(_07363_ ) );
AOI21_X1 _14674_ ( .A(_05767_ ), .B1(_06780_ ), .B2(_06181_ ), .ZN(_07364_ ) );
NAND2_X1 _14675_ ( .A1(_06286_ ), .A2(_06099_ ), .ZN(_07365_ ) );
NAND3_X1 _14676_ ( .A1(_05946_ ), .A2(_06357_ ), .A3(_05948_ ), .ZN(_07366_ ) );
OAI211_X1 _14677_ ( .A(_05880_ ), .B(_07366_ ), .C1(_05942_ ), .C2(_06357_ ), .ZN(_07367_ ) );
NAND3_X1 _14678_ ( .A1(_07365_ ), .A2(_05769_ ), .A3(_07367_ ), .ZN(_07368_ ) );
NAND2_X1 _14679_ ( .A1(_07364_ ), .A2(_07368_ ), .ZN(_07369_ ) );
OAI211_X1 _14680_ ( .A(_05887_ ), .B(_05888_ ), .C1(_04808_ ), .C2(_04806_ ), .ZN(_07370_ ) );
AOI21_X1 _14681_ ( .A(_04809_ ), .B1(_07370_ ), .B2(_05890_ ), .ZN(_07371_ ) );
AOI21_X1 _14682_ ( .A(_07371_ ), .B1(_04807_ ), .B2(_06186_ ), .ZN(_07372_ ) );
AND4_X1 _14683_ ( .A1(_07359_ ), .A2(_07363_ ), .A3(_07369_ ), .A4(_07372_ ), .ZN(_07373_ ) );
AOI21_X1 _14684_ ( .A(_05535_ ), .B1(_07356_ ), .B2(_07373_ ), .ZN(_07374_ ) );
AND2_X1 _14685_ ( .A1(_05379_ ), .A2(_06500_ ), .ZN(_07375_ ) );
NAND2_X1 _14686_ ( .A1(_07350_ ), .A2(_05044_ ), .ZN(_07376_ ) );
NAND3_X1 _14687_ ( .A1(_05967_ ), .A2(_05531_ ), .A3(\EXU.imm_i [26] ), .ZN(_07377_ ) );
NAND3_X1 _14688_ ( .A1(_05970_ ), .A2(\EXU.ls_rdata_i [26] ), .A3(_05971_ ), .ZN(_07378_ ) );
NAND3_X1 _14689_ ( .A1(_07376_ ), .A2(_07377_ ), .A3(_07378_ ), .ZN(_07379_ ) );
OR3_X1 _14690_ ( .A1(_07374_ ), .A2(_07375_ ), .A3(_07379_ ), .ZN(_07380_ ) );
MUX2_X1 _14691_ ( .A(_07355_ ), .B(_07380_ ), .S(_07098_ ), .Z(_07381_ ) );
NAND2_X1 _14692_ ( .A1(_07381_ ), .A2(_07182_ ), .ZN(_07382_ ) );
NAND3_X1 _14693_ ( .A1(_07055_ ), .A2(_05264_ ), .A3(_07355_ ), .ZN(_07383_ ) );
AOI21_X1 _14694_ ( .A(_07058_ ), .B1(_07382_ ), .B2(_07383_ ), .ZN(_07384_ ) );
MUX2_X1 _14695_ ( .A(\EXU.xrd_o [26] ), .B(_07384_ ), .S(_04399_ ), .Z(_00268_ ) );
AOI22_X1 _14696_ ( .A1(_04355_ ), .A2(\EXU.mstatus_i [25] ), .B1(_04336_ ), .B2(\EXU.mcause_i [25] ), .ZN(_07385_ ) );
AOI22_X1 _14697_ ( .A1(_04353_ ), .A2(\EXU.mtvec_i [25] ), .B1(_04350_ ), .B2(\EXU.mepc_i [25] ), .ZN(_07386_ ) );
NAND2_X1 _14698_ ( .A1(_07385_ ), .A2(_07386_ ), .ZN(_07387_ ) );
NAND3_X1 _14699_ ( .A1(_07387_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_6_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A3(_05559_ ), .ZN(_07388_ ) );
AND3_X1 _14700_ ( .A1(_07385_ ), .A2(_07386_ ), .A3(\EXU.xrd_o_$_SDFFCE_PP0P__Q_6_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .ZN(_07389_ ) );
OAI221_X1 _14701_ ( .A(_07388_ ), .B1(_04814_ ), .B2(_06001_ ), .C1(_07389_ ), .C2(_05995_ ), .ZN(_07390_ ) );
AND3_X1 _14702_ ( .A1(_06516_ ), .A2(\EXU.pc_i [25] ), .A3(_05046_ ), .ZN(_07391_ ) );
OR2_X1 _14703_ ( .A1(_07390_ ), .A2(_07391_ ), .ZN(_07392_ ) );
OR2_X1 _14704_ ( .A1(_05394_ ), .A2(_06787_ ), .ZN(_07393_ ) );
NOR2_X1 _14705_ ( .A1(_06844_ ), .A2(_06845_ ), .ZN(_07394_ ) );
AOI21_X1 _14706_ ( .A(_05767_ ), .B1(_07394_ ), .B2(_05914_ ), .ZN(_07395_ ) );
NAND3_X1 _14707_ ( .A1(_06379_ ), .A2(_06380_ ), .A3(_05757_ ), .ZN(_07396_ ) );
AND2_X1 _14708_ ( .A1(_06073_ ), .A2(_06074_ ), .ZN(_07397_ ) );
MUX2_X1 _14709_ ( .A(_06684_ ), .B(_07397_ ), .S(_05755_ ), .Z(_07398_ ) );
OAI21_X1 _14710_ ( .A(_07396_ ), .B1(_07398_ ), .B2(_05960_ ), .ZN(_07399_ ) );
OAI21_X1 _14711_ ( .A(_07395_ ), .B1(_07399_ ), .B2(_05914_ ), .ZN(_07400_ ) );
OAI211_X1 _14712_ ( .A(_05572_ ), .B(_05630_ ), .C1(_04814_ ), .C2(_04813_ ), .ZN(_07401_ ) );
NAND2_X1 _14713_ ( .A1(_07401_ ), .A2(_05556_ ), .ZN(_07402_ ) );
NAND2_X1 _14714_ ( .A1(_07402_ ), .A2(_04815_ ), .ZN(_07403_ ) );
OR3_X1 _14715_ ( .A1(_05635_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_6_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A3(_04813_ ), .ZN(_07404_ ) );
NAND3_X1 _14716_ ( .A1(_07400_ ), .A2(_07403_ ), .A3(_07404_ ), .ZN(_07405_ ) );
AOI21_X1 _14717_ ( .A(_05709_ ), .B1(_05706_ ), .B2(_04674_ ), .ZN(_07406_ ) );
XNOR2_X1 _14718_ ( .A(_07406_ ), .B(_04673_ ), .ZN(_07407_ ) );
OR3_X1 _14719_ ( .A1(_05855_ ), .A2(_06854_ ), .A3(_06363_ ), .ZN(_07408_ ) );
NAND2_X1 _14720_ ( .A1(_05873_ ), .A2(_07408_ ), .ZN(_07409_ ) );
OAI21_X1 _14721_ ( .A(_05880_ ), .B1(_06851_ ), .B2(_06852_ ), .ZN(_07410_ ) );
OAI21_X1 _14722_ ( .A(_07409_ ), .B1(_07410_ ), .B2(_06181_ ), .ZN(_07411_ ) );
AOI221_X2 _14723_ ( .A(_07405_ ), .B1(_05639_ ), .B2(_07407_ ), .C1(_07411_ ), .C2(_06065_ ), .ZN(_07412_ ) );
AOI21_X1 _14724_ ( .A(_05535_ ), .B1(_07393_ ), .B2(_07412_ ), .ZN(_07413_ ) );
AND2_X1 _14725_ ( .A1(_05389_ ), .A2(_06500_ ), .ZN(_07414_ ) );
NAND2_X1 _14726_ ( .A1(_07387_ ), .A2(_05044_ ), .ZN(_07415_ ) );
NAND3_X1 _14727_ ( .A1(_05817_ ), .A2(_05531_ ), .A3(\EXU.imm_i [25] ), .ZN(_07416_ ) );
NAND3_X1 _14728_ ( .A1(_05970_ ), .A2(\EXU.ls_rdata_i [25] ), .A3(_05971_ ), .ZN(_07417_ ) );
NAND3_X1 _14729_ ( .A1(_07415_ ), .A2(_07416_ ), .A3(_07417_ ), .ZN(_07418_ ) );
OR3_X1 _14730_ ( .A1(_07413_ ), .A2(_07414_ ), .A3(_07418_ ), .ZN(_07419_ ) );
MUX2_X1 _14731_ ( .A(_07392_ ), .B(_07419_ ), .S(_07098_ ), .Z(_07420_ ) );
NAND2_X1 _14732_ ( .A1(_07420_ ), .A2(_07182_ ), .ZN(_07421_ ) );
NAND3_X1 _14733_ ( .A1(_07055_ ), .A2(_05264_ ), .A3(_07392_ ), .ZN(_07422_ ) );
AOI21_X1 _14734_ ( .A(_07058_ ), .B1(_07421_ ), .B2(_07422_ ), .ZN(_07423_ ) );
MUX2_X1 _14735_ ( .A(\EXU.xrd_o [25] ), .B(_07423_ ), .S(_04399_ ), .Z(_00269_ ) );
AND3_X1 _14736_ ( .A1(_04352_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05984_ ), .ZN(_07424_ ) );
OAI221_X1 _14737_ ( .A(_05829_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05981_ ), .C1(_05983_ ), .C2(_07424_ ), .ZN(_07425_ ) );
NAND4_X1 _14738_ ( .A1(_05987_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_05988_ ), .ZN(_07426_ ) );
NAND2_X1 _14739_ ( .A1(_07425_ ), .A2(_07426_ ), .ZN(_07427_ ) );
MUX2_X1 _14740_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ), .B(_07427_ ), .S(_05993_ ), .Z(_07428_ ) );
NAND4_X1 _14741_ ( .A1(_04821_ ), .A2(\EXU.funct3_i [1] ), .A3(\EXU.funct3_i [0] ), .A4(fanout_net_10 ), .ZN(_07429_ ) );
AOI22_X1 _14742_ ( .A1(_07428_ ), .A2(_04821_ ), .B1(_05996_ ), .B2(_07429_ ), .ZN(_07430_ ) );
NAND3_X1 _14743_ ( .A1(_06516_ ), .A2(\EXU.pc_i [24] ), .A3(_05999_ ), .ZN(_07431_ ) );
OAI21_X1 _14744_ ( .A(_07431_ ), .B1(_04821_ ), .B2(_06003_ ), .ZN(_07432_ ) );
OAI211_X1 _14745_ ( .A(_04370_ ), .B(_04373_ ), .C1(_07430_ ), .C2(_07432_ ), .ZN(_07433_ ) );
AOI22_X1 _14746_ ( .A1(_06007_ ), .A2(\EXU.ls_rdata_i [24] ), .B1(_06009_ ), .B2(\EXU.imm_i [24] ), .ZN(_07434_ ) );
OAI21_X1 _14747_ ( .A(_07434_ ), .B1(_07428_ ), .B2(_06012_ ), .ZN(_07435_ ) );
NAND2_X1 _14748_ ( .A1(_05396_ ), .A2(_06015_ ), .ZN(_07436_ ) );
NAND3_X1 _14749_ ( .A1(_05954_ ), .A2(_06039_ ), .A3(_05955_ ), .ZN(_07437_ ) );
AOI21_X1 _14750_ ( .A(_05607_ ), .B1(_06143_ ), .B2(_07437_ ), .ZN(_07438_ ) );
AOI211_X1 _14751_ ( .A(_05960_ ), .B(_07438_ ), .C1(_05881_ ), .C2(_07215_ ), .ZN(_07439_ ) );
AOI21_X1 _14752_ ( .A(_05804_ ), .B1(_06437_ ), .B2(_06438_ ), .ZN(_07440_ ) );
OAI21_X1 _14753_ ( .A(_05807_ ), .B1(_07439_ ), .B2(_07440_ ), .ZN(_07441_ ) );
OAI211_X1 _14754_ ( .A(_07441_ ), .B(_04427_ ), .C1(_05769_ ), .C2(_06905_ ), .ZN(_07442_ ) );
OR2_X1 _14755_ ( .A1(_07442_ ), .A2(_05767_ ), .ZN(_07443_ ) );
AND2_X1 _14756_ ( .A1(_06894_ ), .A2(_05868_ ), .ZN(_07444_ ) );
OAI211_X1 _14757_ ( .A(_05872_ ), .B(_05871_ ), .C1(_07444_ ), .C2(_05856_ ), .ZN(_07445_ ) );
OAI21_X1 _14758_ ( .A(_07445_ ), .B1(_06899_ ), .B2(_06063_ ), .ZN(_07446_ ) );
NAND2_X1 _14759_ ( .A1(_07446_ ), .A2(_06066_ ), .ZN(_07447_ ) );
OAI211_X1 _14760_ ( .A(_06313_ ), .B(_06314_ ), .C1(_04821_ ), .C2(_04819_ ), .ZN(_07448_ ) );
AOI21_X1 _14761_ ( .A(_04822_ ), .B1(_07448_ ), .B2(_06316_ ), .ZN(_07449_ ) );
AOI21_X1 _14762_ ( .A(_07449_ ), .B1(_04820_ ), .B2(_06186_ ), .ZN(_07450_ ) );
AOI21_X1 _14763_ ( .A(_05641_ ), .B1(_05706_ ), .B2(_04674_ ), .ZN(_07451_ ) );
OAI21_X1 _14764_ ( .A(_07451_ ), .B1(_04674_ ), .B2(_05706_ ), .ZN(_07452_ ) );
AND4_X1 _14765_ ( .A1(_07443_ ), .A2(_07447_ ), .A3(_07450_ ), .A4(_07452_ ), .ZN(_07453_ ) );
AOI21_X1 _14766_ ( .A(_06014_ ), .B1(_07436_ ), .B2(_07453_ ), .ZN(_07454_ ) );
AOI211_X1 _14767_ ( .A(_07435_ ), .B(_07454_ ), .C1(_05211_ ), .C2(_05401_ ), .ZN(_07455_ ) );
OAI21_X1 _14768_ ( .A(_07433_ ), .B1(_07455_ ), .B2(_04394_ ), .ZN(_07456_ ) );
NAND2_X1 _14769_ ( .A1(_07456_ ), .A2(_07182_ ), .ZN(_07457_ ) );
OAI211_X1 _14770_ ( .A(_06109_ ), .B(_05050_ ), .C1(_07430_ ), .C2(_07432_ ), .ZN(_07458_ ) );
AOI21_X1 _14771_ ( .A(_07058_ ), .B1(_07457_ ), .B2(_07458_ ), .ZN(_07459_ ) );
MUX2_X1 _14772_ ( .A(\EXU.xrd_o [24] ), .B(_07459_ ), .S(_04399_ ), .Z(_00270_ ) );
AOI22_X1 _14773_ ( .A1(_04355_ ), .A2(\EXU.mstatus_i [23] ), .B1(_04336_ ), .B2(\EXU.mcause_i [23] ), .ZN(_07460_ ) );
AOI22_X1 _14774_ ( .A1(_04353_ ), .A2(\EXU.mtvec_i [23] ), .B1(_04350_ ), .B2(\EXU.mepc_i [23] ), .ZN(_07461_ ) );
NAND2_X1 _14775_ ( .A1(_07460_ ), .A2(_07461_ ), .ZN(_07462_ ) );
OAI21_X1 _14776_ ( .A(_05525_ ), .B1(_07462_ ), .B2(_04794_ ), .ZN(_07463_ ) );
NAND3_X1 _14777_ ( .A1(_07462_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_8_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ), .A3(_05559_ ), .ZN(_07464_ ) );
OAI211_X1 _14778_ ( .A(_07463_ ), .B(_07464_ ), .C1(_04792_ ), .C2(_06001_ ), .ZN(_07465_ ) );
AND3_X1 _14779_ ( .A1(_06123_ ), .A2(\EXU.pc_i [23] ), .A3(_05046_ ), .ZN(_07466_ ) );
OR2_X1 _14780_ ( .A1(_07465_ ), .A2(_07466_ ), .ZN(_07467_ ) );
NAND2_X1 _14781_ ( .A1(_05409_ ), .A2(_05585_ ), .ZN(_07468_ ) );
NAND2_X1 _14782_ ( .A1(_06943_ ), .A2(_05769_ ), .ZN(_07469_ ) );
OAI211_X1 _14783_ ( .A(_05871_ ), .B(_05872_ ), .C1(_05856_ ), .C2(_06854_ ), .ZN(_07470_ ) );
AOI21_X1 _14784_ ( .A(_05852_ ), .B1(_07469_ ), .B2(_07470_ ), .ZN(_07471_ ) );
INV_X1 _14785_ ( .A(_04692_ ), .ZN(_07472_ ) );
OAI21_X1 _14786_ ( .A(_04690_ ), .B1(_06018_ ), .B2(_05703_ ), .ZN(_07473_ ) );
AOI21_X1 _14787_ ( .A(_07472_ ), .B1(_07473_ ), .B2(_05689_ ), .ZN(_07474_ ) );
AOI21_X1 _14788_ ( .A(_07474_ ), .B1(\EXU.r1_i [22] ), .B2(_05684_ ), .ZN(_07475_ ) );
XNOR2_X1 _14789_ ( .A(_07475_ ), .B(_04691_ ), .ZN(_07476_ ) );
AND2_X1 _14790_ ( .A1(_07476_ ), .A2(_05639_ ), .ZN(_07477_ ) );
OAI211_X1 _14791_ ( .A(_05887_ ), .B(_05888_ ), .C1(_04792_ ), .C2(_04791_ ), .ZN(_07478_ ) );
AOI21_X1 _14792_ ( .A(_04793_ ), .B1(_07478_ ), .B2(_05890_ ), .ZN(_07479_ ) );
MUX2_X1 _14793_ ( .A(_04795_ ), .B(_07479_ ), .S(_06071_ ), .Z(_07480_ ) );
NAND2_X1 _14794_ ( .A1(_05789_ ), .A2(_06254_ ), .ZN(_07481_ ) );
NAND2_X1 _14795_ ( .A1(_07481_ ), .A2(_05565_ ), .ZN(_07482_ ) );
NAND3_X1 _14796_ ( .A1(_06951_ ), .A2(_05747_ ), .A3(_06952_ ), .ZN(_07483_ ) );
AOI221_X4 _14797_ ( .A(_07482_ ), .B1(_05914_ ), .B2(_07483_ ), .C1(_06060_ ), .C2(_05746_ ), .ZN(_07484_ ) );
NOR4_X1 _14798_ ( .A1(_07471_ ), .A2(_07477_ ), .A3(_07480_ ), .A4(_07484_ ), .ZN(_07485_ ) );
AOI21_X1 _14799_ ( .A(_05535_ ), .B1(_07468_ ), .B2(_07485_ ), .ZN(_07486_ ) );
AND2_X1 _14800_ ( .A1(_05412_ ), .A2(_06500_ ), .ZN(_07487_ ) );
NAND2_X1 _14801_ ( .A1(_07462_ ), .A2(_05044_ ), .ZN(_07488_ ) );
NAND3_X1 _14802_ ( .A1(_05817_ ), .A2(_05531_ ), .A3(\EXU.imm_i [23] ), .ZN(_07489_ ) );
NAND3_X1 _14803_ ( .A1(_04387_ ), .A2(\EXU.ls_rdata_i [23] ), .A3(_04388_ ), .ZN(_07490_ ) );
NAND3_X1 _14804_ ( .A1(_07488_ ), .A2(_07489_ ), .A3(_07490_ ), .ZN(_07491_ ) );
OR3_X1 _14805_ ( .A1(_07486_ ), .A2(_07487_ ), .A3(_07491_ ), .ZN(_07492_ ) );
MUX2_X1 _14806_ ( .A(_07467_ ), .B(_07492_ ), .S(_07098_ ), .Z(_07493_ ) );
NAND2_X1 _14807_ ( .A1(_07493_ ), .A2(_07182_ ), .ZN(_07494_ ) );
NAND3_X1 _14808_ ( .A1(_07055_ ), .A2(_05264_ ), .A3(_07467_ ), .ZN(_07495_ ) );
AOI21_X1 _14809_ ( .A(_04395_ ), .B1(_07494_ ), .B2(_07495_ ), .ZN(_07496_ ) );
MUX2_X1 _14810_ ( .A(\EXU.xrd_o [23] ), .B(_07496_ ), .S(_04399_ ), .Z(_00271_ ) );
AND3_X1 _14811_ ( .A1(_04352_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05984_ ), .ZN(_07497_ ) );
OAI221_X1 _14812_ ( .A(_05829_ ), .B1(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .B2(_05981_ ), .C1(_05983_ ), .C2(_07497_ ), .ZN(_07498_ ) );
NAND4_X1 _14813_ ( .A1(_05987_ ), .A2(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A4(_05988_ ), .ZN(_07499_ ) );
NAND2_X1 _14814_ ( .A1(_07498_ ), .A2(_07499_ ), .ZN(_07500_ ) );
MUX2_X1 _14815_ ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ), .B(_07500_ ), .S(_05993_ ), .Z(_07501_ ) );
NAND4_X1 _14816_ ( .A1(_04785_ ), .A2(\EXU.funct3_i [1] ), .A3(\EXU.funct3_i [0] ), .A4(io_master_arsize_$_ANDNOT__Y_1_B_$_OR__Y_A_$_OR__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_AND__Y_B_$_OR__Y_B ), .ZN(_07502_ ) );
AOI22_X1 _14817_ ( .A1(_07501_ ), .A2(_04785_ ), .B1(_05995_ ), .B2(_07502_ ), .ZN(_07503_ ) );
NAND3_X1 _14818_ ( .A1(_06516_ ), .A2(\EXU.pc_i [22] ), .A3(_05046_ ), .ZN(_07504_ ) );
OAI21_X1 _14819_ ( .A(_07504_ ), .B1(_04785_ ), .B2(_06002_ ), .ZN(_07505_ ) );
OAI211_X1 _14820_ ( .A(_04370_ ), .B(_04373_ ), .C1(_07503_ ), .C2(_07505_ ), .ZN(_07506_ ) );
AOI22_X1 _14821_ ( .A1(_06007_ ), .A2(\EXU.ls_rdata_i [22] ), .B1(_06009_ ), .B2(\EXU.imm_i [22] ), .ZN(_07507_ ) );
OAI21_X1 _14822_ ( .A(_07507_ ), .B1(_07501_ ), .B2(_06012_ ), .ZN(_07508_ ) );
NAND2_X1 _14823_ ( .A1(_05416_ ), .A2(_06015_ ), .ZN(_07509_ ) );
OR2_X1 _14824_ ( .A1(_06984_ ), .A2(_06063_ ), .ZN(_07510_ ) );
NOR2_X1 _14825_ ( .A1(_05864_ ), .A2(_05866_ ), .ZN(_07511_ ) );
OAI211_X1 _14826_ ( .A(_05872_ ), .B(_05871_ ), .C1(_07511_ ), .C2(_05856_ ), .ZN(_07512_ ) );
AOI21_X1 _14827_ ( .A(_05852_ ), .B1(_07510_ ), .B2(_07512_ ), .ZN(_07513_ ) );
AND3_X1 _14828_ ( .A1(_07473_ ), .A2(_07472_ ), .A3(_05689_ ), .ZN(_07514_ ) );
NOR3_X1 _14829_ ( .A1(_07514_ ), .A2(_07474_ ), .A3(_05641_ ), .ZN(_07515_ ) );
NAND3_X1 _14830_ ( .A1(_04782_ ), .A2(\EXU.r1_i [22] ), .A3(_04783_ ), .ZN(_07516_ ) );
NAND3_X1 _14831_ ( .A1(_06313_ ), .A2(_06314_ ), .A3(_07516_ ), .ZN(_07517_ ) );
AOI21_X1 _14832_ ( .A(_04786_ ), .B1(_07517_ ), .B2(_06316_ ), .ZN(_07518_ ) );
MUX2_X1 _14833_ ( .A(_04787_ ), .B(_07518_ ), .S(_06071_ ), .Z(_07519_ ) );
OAI21_X1 _14834_ ( .A(_06254_ ), .B1(_05949_ ), .B2(_05958_ ), .ZN(_07520_ ) );
NAND2_X1 _14835_ ( .A1(_07520_ ), .A2(_05565_ ), .ZN(_07521_ ) );
AOI21_X1 _14836_ ( .A(_05807_ ), .B1(_05925_ ), .B2(_06356_ ), .ZN(_07522_ ) );
AOI211_X1 _14837_ ( .A(_07521_ ), .B(_07522_ ), .C1(_06100_ ), .C2(_05912_ ), .ZN(_07523_ ) );
NOR4_X1 _14838_ ( .A1(_07513_ ), .A2(_07515_ ), .A3(_07519_ ), .A4(_07523_ ), .ZN(_07524_ ) );
AOI21_X1 _14839_ ( .A(_06014_ ), .B1(_07509_ ), .B2(_07524_ ), .ZN(_07525_ ) );
AOI211_X1 _14840_ ( .A(_07508_ ), .B(_07525_ ), .C1(_05211_ ), .C2(_05421_ ), .ZN(_07526_ ) );
OAI21_X1 _14841_ ( .A(_07506_ ), .B1(_07526_ ), .B2(_04394_ ), .ZN(_07527_ ) );
NAND2_X1 _14842_ ( .A1(_07527_ ), .A2(_07182_ ), .ZN(_07528_ ) );
OAI211_X1 _14843_ ( .A(_04376_ ), .B(_05050_ ), .C1(_07503_ ), .C2(_07505_ ), .ZN(_07529_ ) );
AOI21_X1 _14844_ ( .A(_04395_ ), .B1(_07528_ ), .B2(_07529_ ), .ZN(_07530_ ) );
MUX2_X1 _14845_ ( .A(\EXU.xrd_o [22] ), .B(_07530_ ), .S(_04399_ ), .Z(_00272_ ) );
INV_X1 _14846_ ( .A(\ICACHE.burst_counter [0] ), .ZN(_07531_ ) );
AND2_X1 _14847_ ( .A1(_07531_ ), .A2(\ICACHE.burst_counter [1] ), .ZN(_07532_ ) );
NOR2_X1 _14848_ ( .A1(_07531_ ), .A2(\ICACHE.burst_counter [1] ), .ZN(_07533_ ) );
INV_X2 _14849_ ( .A(\ICACHE.s_axi_rready ), .ZN(_07534_ ) );
BUF_X2 _14850_ ( .A(_07534_ ), .Z(_07535_ ) );
NOR3_X1 _14851_ ( .A1(_07532_ ), .A2(_07533_ ), .A3(_07535_ ), .ZN(_07536_ ) );
AND2_X1 _14852_ ( .A1(_07534_ ), .A2(\ICACHE.state_$_MUX__S_A ), .ZN(_07537_ ) );
NOR2_X1 _14853_ ( .A1(_07536_ ), .A2(_07537_ ), .ZN(_07538_ ) );
OAI211_X1 _14854_ ( .A(\CLINT.c_axi_rvalid_$_NOT__A_Y ), .B(_04089_ ), .C1(_04073_ ), .C2(_04097_ ), .ZN(_07539_ ) );
NOR2_X1 _14855_ ( .A1(_04110_ ), .A2(_04113_ ), .ZN(_07540_ ) );
INV_X1 _14856_ ( .A(_07540_ ), .ZN(_07541_ ) );
OAI21_X1 _14857_ ( .A(_07539_ ), .B1(_07541_ ), .B2(io_master_rvalid ), .ZN(_07542_ ) );
INV_X2 _14858_ ( .A(_04058_ ), .ZN(_07543_ ) );
NOR2_X1 _14859_ ( .A1(_07542_ ), .A2(_07543_ ), .ZN(_07544_ ) );
INV_X1 _14860_ ( .A(_07544_ ), .ZN(_07545_ ) );
MUX2_X1 _14861_ ( .A(\ICACHE.burst_counter_$_DFFE_PP__Q_E_$_ANDNOT__Y_B_$_MUX__Y_A ), .B(_07545_ ), .S(\ICACHE.s_axi_rready ), .Z(_07546_ ) );
INV_X1 _14862_ ( .A(\BTB.btag [1] ), .ZN(_07547_ ) );
NAND2_X2 _14863_ ( .A1(_07547_ ), .A2(_07534_ ), .ZN(_07548_ ) );
INV_X1 _14864_ ( .A(\ICACHE.s_axi_araddr [4] ), .ZN(_07549_ ) );
NAND2_X2 _14865_ ( .A1(_07549_ ), .A2(\ICACHE.s_axi_rready ), .ZN(_07550_ ) );
AND2_X2 _14866_ ( .A1(_07548_ ), .A2(_07550_ ), .ZN(_07551_ ) );
MUX2_X1 _14867_ ( .A(\ICACHE.tag_reg[0][1] ), .B(\ICACHE.tag_reg[1][1] ), .S(_07551_ ), .Z(_07552_ ) );
INV_X1 _14868_ ( .A(\BTB.btag [3] ), .ZN(_07553_ ) );
NAND2_X1 _14869_ ( .A1(_07553_ ), .A2(_07534_ ), .ZN(_07554_ ) );
INV_X1 _14870_ ( .A(\ICACHE.s_axi_araddr [6] ), .ZN(_07555_ ) );
NAND2_X1 _14871_ ( .A1(_07555_ ), .A2(\ICACHE.s_axi_rready ), .ZN(_07556_ ) );
AND2_X1 _14872_ ( .A1(_07554_ ), .A2(_07556_ ), .ZN(_07557_ ) );
INV_X1 _14873_ ( .A(_07557_ ), .ZN(_07558_ ) );
MUX2_X1 _14874_ ( .A(\ICACHE.tag_reg[0][3] ), .B(\ICACHE.tag_reg[1][3] ), .S(_07551_ ), .Z(_07559_ ) );
INV_X1 _14875_ ( .A(\BTB.btag [5] ), .ZN(_07560_ ) );
NAND2_X1 _14876_ ( .A1(_07560_ ), .A2(_07534_ ), .ZN(_07561_ ) );
INV_X1 _14877_ ( .A(\ICACHE.s_axi_araddr [8] ), .ZN(_07562_ ) );
NAND2_X1 _14878_ ( .A1(_07562_ ), .A2(\ICACHE.s_axi_rready ), .ZN(_07563_ ) );
AND2_X1 _14879_ ( .A1(_07561_ ), .A2(_07563_ ), .ZN(_07564_ ) );
INV_X1 _14880_ ( .A(_07564_ ), .ZN(_07565_ ) );
OAI22_X1 _14881_ ( .A1(_07552_ ), .A2(_07558_ ), .B1(_07559_ ), .B2(_07565_ ), .ZN(_07566_ ) );
MUX2_X1 _14882_ ( .A(\ICACHE.tag_reg[0][2] ), .B(\ICACHE.tag_reg[1][2] ), .S(_07551_ ), .Z(_07567_ ) );
INV_X1 _14883_ ( .A(_07567_ ), .ZN(_07568_ ) );
NAND2_X1 _14884_ ( .A1(_07534_ ), .A2(\BTB.btag [4] ), .ZN(_07569_ ) );
NAND2_X1 _14885_ ( .A1(\ICACHE.s_axi_araddr [7] ), .A2(\ICACHE.s_axi_rready ), .ZN(_07570_ ) );
NAND2_X1 _14886_ ( .A1(_07569_ ), .A2(_07570_ ), .ZN(_07571_ ) );
AOI221_X4 _14887_ ( .A(_07566_ ), .B1(_07568_ ), .B2(_07571_ ), .C1(_07559_ ), .C2(_07565_ ), .ZN(_07572_ ) );
BUF_X4 _14888_ ( .A(_07551_ ), .Z(_07573_ ) );
MUX2_X1 _14889_ ( .A(\ICACHE.tag_reg[0][5] ), .B(\ICACHE.tag_reg[1][5] ), .S(_07573_ ), .Z(_07574_ ) );
INV_X1 _14890_ ( .A(\BTB.btag [7] ), .ZN(_07575_ ) );
NAND2_X1 _14891_ ( .A1(_07575_ ), .A2(_07534_ ), .ZN(_07576_ ) );
INV_X1 _14892_ ( .A(\ICACHE.s_axi_araddr [10] ), .ZN(_07577_ ) );
NAND2_X1 _14893_ ( .A1(_07577_ ), .A2(\ICACHE.s_axi_rready ), .ZN(_07578_ ) );
AND2_X1 _14894_ ( .A1(_07576_ ), .A2(_07578_ ), .ZN(_07579_ ) );
INV_X1 _14895_ ( .A(_07579_ ), .ZN(_07580_ ) );
MUX2_X1 _14896_ ( .A(\ICACHE.tag_reg[0][9] ), .B(\ICACHE.tag_reg[1][9] ), .S(_07573_ ), .Z(_07581_ ) );
INV_X1 _14897_ ( .A(\BTB.btag [11] ), .ZN(_07582_ ) );
NAND2_X1 _14898_ ( .A1(_07582_ ), .A2(_07535_ ), .ZN(_07583_ ) );
INV_X1 _14899_ ( .A(\ICACHE.s_axi_araddr [14] ), .ZN(_07584_ ) );
NAND2_X1 _14900_ ( .A1(_07584_ ), .A2(\ICACHE.s_axi_rready ), .ZN(_07585_ ) );
AND2_X1 _14901_ ( .A1(_07583_ ), .A2(_07585_ ), .ZN(_07586_ ) );
INV_X1 _14902_ ( .A(_07586_ ), .ZN(_07587_ ) );
AOI22_X1 _14903_ ( .A1(_07574_ ), .A2(_07580_ ), .B1(_07581_ ), .B2(_07587_ ), .ZN(_07588_ ) );
OR2_X1 _14904_ ( .A1(_07581_ ), .A2(_07587_ ), .ZN(_07589_ ) );
MUX2_X1 _14905_ ( .A(\ICACHE.tag_reg[0][8] ), .B(\ICACHE.tag_reg[1][8] ), .S(_07573_ ), .Z(_07590_ ) );
INV_X1 _14906_ ( .A(\BTB.btag [10] ), .ZN(_07591_ ) );
NAND2_X1 _14907_ ( .A1(_07591_ ), .A2(_07535_ ), .ZN(_07592_ ) );
INV_X1 _14908_ ( .A(\ICACHE.s_axi_araddr [13] ), .ZN(_07593_ ) );
NAND2_X1 _14909_ ( .A1(_07593_ ), .A2(\ICACHE.s_axi_rready ), .ZN(_07594_ ) );
AND2_X1 _14910_ ( .A1(_07592_ ), .A2(_07594_ ), .ZN(_07595_ ) );
INV_X1 _14911_ ( .A(_07595_ ), .ZN(_07596_ ) );
NAND2_X1 _14912_ ( .A1(_07590_ ), .A2(_07596_ ), .ZN(_07597_ ) );
AND4_X1 _14913_ ( .A1(_07572_ ), .A2(_07588_ ), .A3(_07589_ ), .A4(_07597_ ), .ZN(_07598_ ) );
INV_X1 _14914_ ( .A(\ICACHE.tag_reg[0][0] ), .ZN(_07599_ ) );
INV_X1 _14915_ ( .A(\ICACHE.tag_reg[1][0] ), .ZN(_07600_ ) );
BUF_X4 _14916_ ( .A(_07573_ ), .Z(_07601_ ) );
MUX2_X1 _14917_ ( .A(_07599_ ), .B(_07600_ ), .S(_07601_ ), .Z(_07602_ ) );
INV_X1 _14918_ ( .A(\BTB.btag [2] ), .ZN(_07603_ ) );
NAND2_X1 _14919_ ( .A1(_07603_ ), .A2(_07535_ ), .ZN(_07604_ ) );
INV_X1 _14920_ ( .A(\ICACHE.s_axi_araddr [5] ), .ZN(_07605_ ) );
NAND2_X1 _14921_ ( .A1(_07605_ ), .A2(\ICACHE.s_axi_rready ), .ZN(_07606_ ) );
NAND2_X1 _14922_ ( .A1(_07604_ ), .A2(_07606_ ), .ZN(_07607_ ) );
XNOR2_X1 _14923_ ( .A(_07602_ ), .B(_07607_ ), .ZN(_07608_ ) );
MUX2_X1 _14924_ ( .A(\ICACHE.tag_reg[0][7] ), .B(\ICACHE.tag_reg[1][7] ), .S(_07601_ ), .Z(_07609_ ) );
INV_X1 _14925_ ( .A(\BTB.btag [9] ), .ZN(_07610_ ) );
NOR2_X1 _14926_ ( .A1(_07610_ ), .A2(\ICACHE.s_axi_rready ), .ZN(_07611_ ) );
AND2_X1 _14927_ ( .A1(\ICACHE.s_axi_araddr [12] ), .A2(\ICACHE.s_axi_rready ), .ZN(_07612_ ) );
NOR2_X1 _14928_ ( .A1(_07611_ ), .A2(_07612_ ), .ZN(_07613_ ) );
XOR2_X1 _14929_ ( .A(_07609_ ), .B(_07613_ ), .Z(_07614_ ) );
MUX2_X1 _14930_ ( .A(\ICACHE.tag_reg[0][6] ), .B(\ICACHE.tag_reg[1][6] ), .S(_07601_ ), .Z(_07615_ ) );
INV_X1 _14931_ ( .A(\BTB.btag [8] ), .ZN(_07616_ ) );
NAND2_X1 _14932_ ( .A1(_07616_ ), .A2(_07535_ ), .ZN(_07617_ ) );
INV_X1 _14933_ ( .A(\ICACHE.s_axi_araddr [11] ), .ZN(_07618_ ) );
NAND2_X1 _14934_ ( .A1(_07618_ ), .A2(\ICACHE.s_axi_rready ), .ZN(_07619_ ) );
NAND2_X1 _14935_ ( .A1(_07617_ ), .A2(_07619_ ), .ZN(_07620_ ) );
XOR2_X1 _14936_ ( .A(_07615_ ), .B(_07620_ ), .Z(_07621_ ) );
NAND4_X1 _14937_ ( .A1(_07598_ ), .A2(_07608_ ), .A3(_07614_ ), .A4(_07621_ ), .ZN(_07622_ ) );
MUX2_X1 _14938_ ( .A(\ICACHE.tag_reg[0][4] ), .B(\ICACHE.tag_reg[1][4] ), .S(_07573_ ), .Z(_07623_ ) );
INV_X1 _14939_ ( .A(\BTB.btag [6] ), .ZN(_07624_ ) );
NAND2_X1 _14940_ ( .A1(_07624_ ), .A2(_07534_ ), .ZN(_07625_ ) );
INV_X1 _14941_ ( .A(\ICACHE.s_axi_araddr [9] ), .ZN(_07626_ ) );
NAND2_X1 _14942_ ( .A1(_07626_ ), .A2(\ICACHE.s_axi_rready ), .ZN(_07627_ ) );
AND2_X1 _14943_ ( .A1(_07625_ ), .A2(_07627_ ), .ZN(_07628_ ) );
INV_X1 _14944_ ( .A(_07628_ ), .ZN(_07629_ ) );
NOR2_X1 _14945_ ( .A1(_07623_ ), .A2(_07629_ ), .ZN(_07630_ ) );
MUX2_X1 _14946_ ( .A(\ICACHE.tag_reg[0][10] ), .B(\ICACHE.tag_reg[1][10] ), .S(_07573_ ), .Z(_07631_ ) );
INV_X1 _14947_ ( .A(\BTB.btag [12] ), .ZN(_07632_ ) );
NAND2_X1 _14948_ ( .A1(_07632_ ), .A2(_07535_ ), .ZN(_07633_ ) );
INV_X1 _14949_ ( .A(\ICACHE.s_axi_araddr [15] ), .ZN(_07634_ ) );
NAND2_X1 _14950_ ( .A1(_07634_ ), .A2(\ICACHE.s_axi_rready ), .ZN(_07635_ ) );
AND2_X1 _14951_ ( .A1(_07633_ ), .A2(_07635_ ), .ZN(_07636_ ) );
INV_X1 _14952_ ( .A(_07636_ ), .ZN(_07637_ ) );
AOI21_X1 _14953_ ( .A(_07630_ ), .B1(_07631_ ), .B2(_07637_ ), .ZN(_07638_ ) );
OAI221_X1 _14954_ ( .A(_07638_ ), .B1(_07631_ ), .B2(_07637_ ), .C1(_07568_ ), .C2(_07571_ ), .ZN(_07639_ ) );
MUX2_X1 _14955_ ( .A(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_07573_ ), .Z(_07640_ ) );
MUX2_X1 _14956_ ( .A(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(_07573_ ), .Z(_07641_ ) );
NAND2_X1 _14957_ ( .A1(_07534_ ), .A2(\BTB.bindex ), .ZN(_07642_ ) );
NAND2_X1 _14958_ ( .A1(\ICACHE.s_axi_araddr [2] ), .A2(\ICACHE.s_axi_rready ), .ZN(_07643_ ) );
AND2_X1 _14959_ ( .A1(_07642_ ), .A2(_07643_ ), .ZN(_07644_ ) );
BUF_X4 _14960_ ( .A(_07644_ ), .Z(_07645_ ) );
INV_X2 _14961_ ( .A(_07645_ ), .ZN(_07646_ ) );
MUX2_X1 _14962_ ( .A(_07640_ ), .B(_07641_ ), .S(_07646_ ), .Z(_07647_ ) );
MUX2_X1 _14963_ ( .A(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(_07573_ ), .Z(_07648_ ) );
MUX2_X1 _14964_ ( .A(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(_07573_ ), .Z(_07649_ ) );
MUX2_X1 _14965_ ( .A(_07648_ ), .B(_07649_ ), .S(_07646_ ), .Z(_07650_ ) );
AND2_X1 _14966_ ( .A1(\ICACHE.s_axi_rready ), .A2(\ICACHE.state_$_MUX__S_B ), .ZN(_07651_ ) );
NOR2_X2 _14967_ ( .A1(_07537_ ), .A2(_07651_ ), .ZN(_07652_ ) );
MUX2_X1 _14968_ ( .A(_07647_ ), .B(_07650_ ), .S(_07652_ ), .Z(_07653_ ) );
NOR2_X1 _14969_ ( .A1(_07574_ ), .A2(_07580_ ), .ZN(_07654_ ) );
AOI21_X1 _14970_ ( .A(_07654_ ), .B1(_07623_ ), .B2(_07629_ ), .ZN(_07655_ ) );
NAND2_X1 _14971_ ( .A1(_07552_ ), .A2(_07558_ ), .ZN(_07656_ ) );
OAI211_X1 _14972_ ( .A(_07655_ ), .B(_07656_ ), .C1(_07590_ ), .C2(_07596_ ), .ZN(_07657_ ) );
OR3_X1 _14973_ ( .A1(_07639_ ), .A2(_07653_ ), .A3(_07657_ ), .ZN(_07658_ ) );
NOR2_X1 _14974_ ( .A1(_07622_ ), .A2(_07658_ ), .ZN(_07659_ ) );
AND2_X2 _14975_ ( .A1(_07535_ ), .A2(\ICACHE.m_axi_arvalid ), .ZN(_07660_ ) );
XNOR2_X1 _14976_ ( .A(\BTB.pc_i [23] ), .B(\ICACHE.tag_check [7] ), .ZN(_07661_ ) );
XNOR2_X1 _14977_ ( .A(\BTB.pc_i [22] ), .B(\ICACHE.tag_check [6] ), .ZN(_07662_ ) );
XNOR2_X1 _14978_ ( .A(\BTB.pc_i [25] ), .B(\ICACHE.tag_check [9] ), .ZN(_07663_ ) );
XNOR2_X1 _14979_ ( .A(\BTB.pc_i [26] ), .B(\ICACHE.tag_check [10] ), .ZN(_07664_ ) );
AND4_X1 _14980_ ( .A1(_07661_ ), .A2(_07662_ ), .A3(_07663_ ), .A4(_07664_ ), .ZN(_07665_ ) );
XOR2_X1 _14981_ ( .A(\BTB.pc_i [27] ), .B(\ICACHE.tag_check [11] ), .Z(_07666_ ) );
XOR2_X1 _14982_ ( .A(\BTB.pc_i [20] ), .B(\ICACHE.tag_check [4] ), .Z(_07667_ ) );
XOR2_X1 _14983_ ( .A(\BTB.pc_i [30] ), .B(\ICACHE.tag_check [14] ), .Z(_07668_ ) );
XOR2_X1 _14984_ ( .A(\BTB.pc_i [24] ), .B(\ICACHE.tag_check [8] ), .Z(_07669_ ) );
NOR4_X1 _14985_ ( .A1(_07666_ ), .A2(_07667_ ), .A3(_07668_ ), .A4(_07669_ ), .ZN(_07670_ ) );
XOR2_X1 _14986_ ( .A(\BTB.pc_i [18] ), .B(\ICACHE.tag_check [2] ), .Z(_07671_ ) );
XOR2_X1 _14987_ ( .A(\BTB.pc_i [21] ), .B(\ICACHE.tag_check [5] ), .Z(_07672_ ) );
XOR2_X1 _14988_ ( .A(\BTB.pc_i [19] ), .B(\ICACHE.tag_check [3] ), .Z(_07673_ ) );
XOR2_X1 _14989_ ( .A(\BTB.pc_i [17] ), .B(\ICACHE.tag_check [1] ), .Z(_07674_ ) );
NOR4_X1 _14990_ ( .A1(_07671_ ), .A2(_07672_ ), .A3(_07673_ ), .A4(_07674_ ), .ZN(_07675_ ) );
XNOR2_X1 _14991_ ( .A(\BTB.pc_i [29] ), .B(\ICACHE.tag_check [13] ), .ZN(_07676_ ) );
XNOR2_X1 _14992_ ( .A(\BTB.pc_i [16] ), .B(\ICACHE.tag_check [0] ), .ZN(_07677_ ) );
XNOR2_X1 _14993_ ( .A(\BTB.pc_i [28] ), .B(\ICACHE.tag_check [12] ), .ZN(_07678_ ) );
XNOR2_X1 _14994_ ( .A(\BTB.pc_i [31] ), .B(\ICACHE.tag_check [15] ), .ZN(_07679_ ) );
AND4_X1 _14995_ ( .A1(_07676_ ), .A2(_07677_ ), .A3(_07678_ ), .A4(_07679_ ), .ZN(_07680_ ) );
AND4_X1 _14996_ ( .A1(_07665_ ), .A2(_07670_ ), .A3(_07675_ ), .A4(_07680_ ), .ZN(_07681_ ) );
NAND4_X1 _14997_ ( .A1(_07659_ ), .A2(\ICACHE.m_axi_arready ), .A3(_07660_ ), .A4(_07681_ ), .ZN(_07682_ ) );
AND2_X1 _14998_ ( .A1(_07682_ ), .A2(_03805_ ), .ZN(_07683_ ) );
INV_X1 _14999_ ( .A(_07683_ ), .ZN(_07684_ ) );
OR2_X1 _15000_ ( .A1(_07546_ ), .A2(_07684_ ), .ZN(_07685_ ) );
MUX2_X1 _15001_ ( .A(_07538_ ), .B(\ICACHE.burst_counter [1] ), .S(_07685_ ), .Z(_00273_ ) );
MUX2_X1 _15002_ ( .A(\BTB.bindex ), .B(\ICACHE.burst_counter_$_DFFE_PP__Q_1_D_$_MUX__Y_B ), .S(\ICACHE.s_axi_rready ), .Z(_07686_ ) );
MUX2_X1 _15003_ ( .A(_07686_ ), .B(\ICACHE.burst_counter [0] ), .S(_07685_ ), .Z(_00274_ ) );
OAI211_X1 _15004_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_B_$_MUX__Y_A ), .B(_04089_ ), .C1(_04074_ ), .C2(_04098_ ), .ZN(_07687_ ) );
OAI21_X1 _15005_ ( .A(_07687_ ), .B1(_07541_ ), .B2(\io_master_rdata [31] ), .ZN(_07688_ ) );
BUF_X2 _15006_ ( .A(_07543_ ), .Z(\io_master_awburst [0] ) );
NOR2_X1 _15007_ ( .A1(_07688_ ), .A2(\io_master_awburst [0] ), .ZN(_07689_ ) );
INV_X1 _15008_ ( .A(\ICACHE.m_axi_arready ), .ZN(_07690_ ) );
AND2_X1 _15009_ ( .A1(_07544_ ), .A2(_07690_ ), .ZN(_07691_ ) );
AND2_X1 _15010_ ( .A1(_07691_ ), .A2(_03798_ ), .ZN(_07692_ ) );
INV_X2 _15011_ ( .A(_07601_ ), .ZN(_07693_ ) );
AND2_X1 _15012_ ( .A1(_07692_ ), .A2(_07693_ ), .ZN(_07694_ ) );
NOR2_X1 _15013_ ( .A1(\ICACHE.burst_counter [1] ), .A2(\ICACHE.burst_counter [0] ), .ZN(_07695_ ) );
NAND2_X1 _15014_ ( .A1(_07694_ ), .A2(_07695_ ), .ZN(_07696_ ) );
BUF_X4 _15015_ ( .A(_07696_ ), .Z(_07697_ ) );
MUX2_X1 _15016_ ( .A(_07689_ ), .B(\ICACHE.cache_reg[0][31] ), .S(_07697_ ), .Z(_00275_ ) );
BUF_X4 _15017_ ( .A(_04089_ ), .Z(_07698_ ) );
OAI211_X1 _15018_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_1_B_$_MUX__Y_A ), .B(_07698_ ), .C1(_04075_ ), .C2(_04099_ ), .ZN(_07699_ ) );
BUF_X4 _15019_ ( .A(_07541_ ), .Z(_07700_ ) );
OAI21_X1 _15020_ ( .A(_07699_ ), .B1(_07700_ ), .B2(\io_master_rdata [30] ), .ZN(_07701_ ) );
NOR2_X1 _15021_ ( .A1(_07701_ ), .A2(\io_master_awburst [0] ), .ZN(_07702_ ) );
MUX2_X1 _15022_ ( .A(_07702_ ), .B(\ICACHE.cache_reg[0][30] ), .S(_07697_ ), .Z(_00276_ ) );
BUF_X4 _15023_ ( .A(_04075_ ), .Z(_07703_ ) );
BUF_X4 _15024_ ( .A(_04099_ ), .Z(_07704_ ) );
OAI211_X1 _15025_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_10_B_$_MUX__Y_A ), .B(_04091_ ), .C1(_07703_ ), .C2(_07704_ ), .ZN(_07705_ ) );
BUF_X4 _15026_ ( .A(_07700_ ), .Z(_07706_ ) );
OAI21_X1 _15027_ ( .A(_07705_ ), .B1(_07706_ ), .B2(\io_master_rdata [21] ), .ZN(_07707_ ) );
NOR2_X1 _15028_ ( .A1(_07707_ ), .A2(\io_master_awburst [0] ), .ZN(_07708_ ) );
MUX2_X1 _15029_ ( .A(_07708_ ), .B(\ICACHE.cache_reg[0][21] ), .S(_07697_ ), .Z(_00277_ ) );
OAI211_X1 _15030_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_11_B_$_MUX__Y_A ), .B(_04091_ ), .C1(_04076_ ), .C2(_04100_ ), .ZN(_07709_ ) );
OAI21_X1 _15031_ ( .A(_07709_ ), .B1(_07706_ ), .B2(\io_master_rdata [20] ), .ZN(_07710_ ) );
NOR2_X1 _15032_ ( .A1(_07710_ ), .A2(\io_master_awburst [0] ), .ZN(_07711_ ) );
MUX2_X1 _15033_ ( .A(_07711_ ), .B(\ICACHE.cache_reg[0][20] ), .S(_07697_ ), .Z(_00278_ ) );
OAI211_X1 _15034_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_12_B_$_MUX__Y_A ), .B(_04091_ ), .C1(_04076_ ), .C2(_04100_ ), .ZN(_07712_ ) );
OAI21_X1 _15035_ ( .A(_07712_ ), .B1(_07706_ ), .B2(\io_master_rdata [19] ), .ZN(_07713_ ) );
NOR2_X1 _15036_ ( .A1(_07713_ ), .A2(\io_master_awburst [0] ), .ZN(_07714_ ) );
MUX2_X1 _15037_ ( .A(_07714_ ), .B(\ICACHE.cache_reg[0][19] ), .S(_07697_ ), .Z(_00279_ ) );
OAI211_X1 _15038_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_13_B_$_MUX__Y_A ), .B(_04091_ ), .C1(_07703_ ), .C2(_07704_ ), .ZN(_07715_ ) );
OAI21_X1 _15039_ ( .A(_07715_ ), .B1(_07706_ ), .B2(\io_master_rdata [18] ), .ZN(_07716_ ) );
NOR2_X1 _15040_ ( .A1(_07716_ ), .A2(\io_master_awburst [0] ), .ZN(_07717_ ) );
MUX2_X1 _15041_ ( .A(_07717_ ), .B(\ICACHE.cache_reg[0][18] ), .S(_07697_ ), .Z(_00280_ ) );
OAI211_X1 _15042_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_14_B_$_MUX__Y_A ), .B(_07698_ ), .C1(_07703_ ), .C2(_07704_ ), .ZN(_07718_ ) );
OAI21_X1 _15043_ ( .A(_07718_ ), .B1(_07700_ ), .B2(\io_master_rdata [17] ), .ZN(_07719_ ) );
BUF_X4 _15044_ ( .A(_07543_ ), .Z(_07720_ ) );
NOR2_X1 _15045_ ( .A1(_07719_ ), .A2(_07720_ ), .ZN(_07721_ ) );
MUX2_X1 _15046_ ( .A(_07721_ ), .B(\ICACHE.cache_reg[0][17] ), .S(_07697_ ), .Z(_00281_ ) );
OAI211_X1 _15047_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_15_B_$_MUX__Y_A ), .B(_07698_ ), .C1(_07703_ ), .C2(_07704_ ), .ZN(_07722_ ) );
OAI21_X1 _15048_ ( .A(_07722_ ), .B1(_07700_ ), .B2(\io_master_rdata [16] ), .ZN(_07723_ ) );
NOR2_X1 _15049_ ( .A1(_07723_ ), .A2(_07720_ ), .ZN(_07724_ ) );
MUX2_X1 _15050_ ( .A(_07724_ ), .B(\ICACHE.cache_reg[0][16] ), .S(_07697_ ), .Z(_00282_ ) );
OAI211_X1 _15051_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_16_B_$_MUX__Y_A ), .B(_04089_ ), .C1(_04074_ ), .C2(_04098_ ), .ZN(_07725_ ) );
OAI21_X1 _15052_ ( .A(_07725_ ), .B1(_07541_ ), .B2(\io_master_rdata [15] ), .ZN(_07726_ ) );
NOR2_X1 _15053_ ( .A1(_07726_ ), .A2(_07720_ ), .ZN(_07727_ ) );
MUX2_X1 _15054_ ( .A(_07727_ ), .B(\ICACHE.cache_reg[0][15] ), .S(_07697_ ), .Z(_00283_ ) );
OAI211_X1 _15055_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_17_B_$_MUX__Y_A ), .B(_04089_ ), .C1(_04074_ ), .C2(_04098_ ), .ZN(_07728_ ) );
BUF_X4 _15056_ ( .A(_07541_ ), .Z(_07729_ ) );
OAI21_X1 _15057_ ( .A(_07728_ ), .B1(_07729_ ), .B2(\io_master_rdata [14] ), .ZN(_07730_ ) );
NOR2_X1 _15058_ ( .A1(_07730_ ), .A2(_07720_ ), .ZN(_07731_ ) );
MUX2_X1 _15059_ ( .A(_07731_ ), .B(\ICACHE.cache_reg[0][14] ), .S(_07697_ ), .Z(_00284_ ) );
OAI211_X1 _15060_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_18_B_$_MUX__Y_A ), .B(_04090_ ), .C1(_04074_ ), .C2(_04098_ ), .ZN(_07732_ ) );
OAI21_X1 _15061_ ( .A(_07732_ ), .B1(_07729_ ), .B2(\io_master_rdata [13] ), .ZN(_07733_ ) );
NOR2_X1 _15062_ ( .A1(_07733_ ), .A2(_07720_ ), .ZN(_07734_ ) );
BUF_X4 _15063_ ( .A(_07696_ ), .Z(_07735_ ) );
MUX2_X1 _15064_ ( .A(_07734_ ), .B(\ICACHE.cache_reg[0][13] ), .S(_07735_ ), .Z(_00285_ ) );
OAI211_X1 _15065_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_19_B_$_MUX__Y_A ), .B(_04090_ ), .C1(_04074_ ), .C2(_04098_ ), .ZN(_07736_ ) );
OAI21_X1 _15066_ ( .A(_07736_ ), .B1(_07729_ ), .B2(\io_master_rdata [12] ), .ZN(_07737_ ) );
NOR2_X1 _15067_ ( .A1(_07737_ ), .A2(_07720_ ), .ZN(_07738_ ) );
MUX2_X1 _15068_ ( .A(_07738_ ), .B(\ICACHE.cache_reg[0][12] ), .S(_07735_ ), .Z(_00286_ ) );
OAI211_X1 _15069_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_2_B_$_MUX__Y_A ), .B(_04090_ ), .C1(_04075_ ), .C2(_04099_ ), .ZN(_07739_ ) );
OAI21_X1 _15070_ ( .A(_07739_ ), .B1(_07729_ ), .B2(\io_master_rdata [29] ), .ZN(_07740_ ) );
NOR2_X1 _15071_ ( .A1(_07740_ ), .A2(_07720_ ), .ZN(_07741_ ) );
MUX2_X1 _15072_ ( .A(_07741_ ), .B(\ICACHE.cache_reg[0][29] ), .S(_07735_ ), .Z(_00287_ ) );
OAI211_X1 _15073_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_20_B_$_MUX__Y_A ), .B(_07698_ ), .C1(_04075_ ), .C2(_04099_ ), .ZN(_07742_ ) );
OAI21_X1 _15074_ ( .A(_07742_ ), .B1(_07700_ ), .B2(\io_master_rdata [11] ), .ZN(_07743_ ) );
NOR2_X1 _15075_ ( .A1(_07743_ ), .A2(_07720_ ), .ZN(_07744_ ) );
MUX2_X1 _15076_ ( .A(_07744_ ), .B(\ICACHE.cache_reg[0][11] ), .S(_07735_ ), .Z(_00288_ ) );
OAI211_X1 _15077_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_21_B_$_MUX__Y_A ), .B(_04090_ ), .C1(_04074_ ), .C2(_04098_ ), .ZN(_07745_ ) );
OAI21_X1 _15078_ ( .A(_07745_ ), .B1(_07729_ ), .B2(\io_master_rdata [10] ), .ZN(_07746_ ) );
NOR2_X1 _15079_ ( .A1(_07746_ ), .A2(_07720_ ), .ZN(_07747_ ) );
MUX2_X1 _15080_ ( .A(_07747_ ), .B(\ICACHE.cache_reg[0][10] ), .S(_07735_ ), .Z(_00289_ ) );
OAI211_X1 _15081_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_22_B_$_MUX__Y_A ), .B(_07698_ ), .C1(_04075_ ), .C2(_04099_ ), .ZN(_07748_ ) );
OAI21_X1 _15082_ ( .A(_07748_ ), .B1(_07700_ ), .B2(\io_master_rdata [9] ), .ZN(_07749_ ) );
NOR2_X1 _15083_ ( .A1(_07749_ ), .A2(_07720_ ), .ZN(_07750_ ) );
MUX2_X1 _15084_ ( .A(_07750_ ), .B(\ICACHE.cache_reg[0][9] ), .S(_07735_ ), .Z(_00290_ ) );
OAI211_X1 _15085_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_23_B_$_MUX__Y_A ), .B(_04090_ ), .C1(_04074_ ), .C2(_04098_ ), .ZN(_07751_ ) );
OAI21_X1 _15086_ ( .A(_07751_ ), .B1(_07729_ ), .B2(\io_master_rdata [8] ), .ZN(_07752_ ) );
BUF_X4 _15087_ ( .A(_07543_ ), .Z(_07753_ ) );
NOR2_X1 _15088_ ( .A1(_07752_ ), .A2(_07753_ ), .ZN(_07754_ ) );
MUX2_X1 _15089_ ( .A(_07754_ ), .B(\ICACHE.cache_reg[0][8] ), .S(_07735_ ), .Z(_00291_ ) );
OAI211_X1 _15090_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_24_B_$_MUX__Y_A ), .B(_07698_ ), .C1(_04075_ ), .C2(_04099_ ), .ZN(_07755_ ) );
OAI21_X1 _15091_ ( .A(_07755_ ), .B1(_07700_ ), .B2(\io_master_rdata [7] ), .ZN(_07756_ ) );
NOR2_X1 _15092_ ( .A1(_07756_ ), .A2(_07753_ ), .ZN(_07757_ ) );
MUX2_X1 _15093_ ( .A(_07757_ ), .B(\ICACHE.cache_reg[0][7] ), .S(_07735_ ), .Z(_00292_ ) );
OAI211_X1 _15094_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_25_B_$_MUX__Y_A ), .B(_04091_ ), .C1(_07703_ ), .C2(_07704_ ), .ZN(_07758_ ) );
OAI21_X1 _15095_ ( .A(_07758_ ), .B1(_07706_ ), .B2(\io_master_rdata [6] ), .ZN(_07759_ ) );
NOR2_X1 _15096_ ( .A1(_07759_ ), .A2(_07753_ ), .ZN(_07760_ ) );
MUX2_X1 _15097_ ( .A(_07760_ ), .B(\ICACHE.cache_reg[0][6] ), .S(_07735_ ), .Z(_00293_ ) );
OAI211_X1 _15098_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_26_B_$_MUX__Y_A ), .B(_07698_ ), .C1(_07703_ ), .C2(_07704_ ), .ZN(_07761_ ) );
OAI21_X1 _15099_ ( .A(_07761_ ), .B1(_07706_ ), .B2(\io_master_rdata [5] ), .ZN(_07762_ ) );
NOR2_X1 _15100_ ( .A1(_07762_ ), .A2(_07753_ ), .ZN(_07763_ ) );
MUX2_X1 _15101_ ( .A(_07763_ ), .B(\ICACHE.cache_reg[0][5] ), .S(_07735_ ), .Z(_00294_ ) );
OAI211_X1 _15102_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_27_B_$_MUX__Y_A ), .B(_04091_ ), .C1(_04076_ ), .C2(_04100_ ), .ZN(_07764_ ) );
OAI21_X1 _15103_ ( .A(_07764_ ), .B1(_07706_ ), .B2(\io_master_rdata [4] ), .ZN(_07765_ ) );
NOR2_X1 _15104_ ( .A1(_07765_ ), .A2(_07753_ ), .ZN(_07766_ ) );
BUF_X4 _15105_ ( .A(_07696_ ), .Z(_07767_ ) );
MUX2_X1 _15106_ ( .A(_07766_ ), .B(\ICACHE.cache_reg[0][4] ), .S(_07767_ ), .Z(_00295_ ) );
OAI211_X1 _15107_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_28_B_$_MUX__Y_A ), .B(_04091_ ), .C1(_04076_ ), .C2(_04100_ ), .ZN(_07768_ ) );
OAI21_X1 _15108_ ( .A(_07768_ ), .B1(_07706_ ), .B2(\io_master_rdata [3] ), .ZN(_07769_ ) );
NOR2_X1 _15109_ ( .A1(_07769_ ), .A2(_07753_ ), .ZN(_07770_ ) );
MUX2_X1 _15110_ ( .A(_07770_ ), .B(\ICACHE.cache_reg[0][3] ), .S(_07767_ ), .Z(_00296_ ) );
OAI211_X1 _15111_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_29_B_$_MUX__Y_A ), .B(_07698_ ), .C1(_07703_ ), .C2(_07704_ ), .ZN(_07771_ ) );
OAI21_X1 _15112_ ( .A(_07771_ ), .B1(_07700_ ), .B2(\io_master_rdata [2] ), .ZN(_07772_ ) );
NOR2_X1 _15113_ ( .A1(_07772_ ), .A2(_07753_ ), .ZN(_07773_ ) );
MUX2_X1 _15114_ ( .A(_07773_ ), .B(\ICACHE.cache_reg[0][2] ), .S(_07767_ ), .Z(_00297_ ) );
OAI211_X1 _15115_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_3_B_$_MUX__Y_A ), .B(_07698_ ), .C1(_07703_ ), .C2(_07704_ ), .ZN(_07774_ ) );
OAI21_X1 _15116_ ( .A(_07774_ ), .B1(_07700_ ), .B2(\io_master_rdata [28] ), .ZN(_07775_ ) );
NOR2_X1 _15117_ ( .A1(_07775_ ), .A2(_07753_ ), .ZN(_07776_ ) );
MUX2_X1 _15118_ ( .A(_07776_ ), .B(\ICACHE.cache_reg[0][28] ), .S(_07767_ ), .Z(_00298_ ) );
OAI211_X1 _15119_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_4_B_$_MUX__Y_A ), .B(_04090_ ), .C1(_04075_ ), .C2(_04099_ ), .ZN(_07777_ ) );
OAI21_X1 _15120_ ( .A(_07777_ ), .B1(_07729_ ), .B2(\io_master_rdata [27] ), .ZN(_07778_ ) );
NOR2_X1 _15121_ ( .A1(_07778_ ), .A2(_07753_ ), .ZN(_07779_ ) );
MUX2_X1 _15122_ ( .A(_07779_ ), .B(\ICACHE.cache_reg[0][27] ), .S(_07767_ ), .Z(_00299_ ) );
OAI211_X1 _15123_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_5_B_$_MUX__Y_A ), .B(_04090_ ), .C1(_04075_ ), .C2(_04099_ ), .ZN(_07780_ ) );
OAI21_X1 _15124_ ( .A(_07780_ ), .B1(_07729_ ), .B2(\io_master_rdata [26] ), .ZN(_07781_ ) );
NOR2_X1 _15125_ ( .A1(_07781_ ), .A2(_07753_ ), .ZN(_07782_ ) );
MUX2_X1 _15126_ ( .A(_07782_ ), .B(\ICACHE.cache_reg[0][26] ), .S(_07767_ ), .Z(_00300_ ) );
OAI211_X1 _15127_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_6_B_$_MUX__Y_A ), .B(_04090_ ), .C1(_04074_ ), .C2(_04098_ ), .ZN(_07783_ ) );
OAI21_X1 _15128_ ( .A(_07783_ ), .B1(_07729_ ), .B2(\io_master_rdata [25] ), .ZN(_07784_ ) );
NOR2_X1 _15129_ ( .A1(_07784_ ), .A2(_07543_ ), .ZN(_07785_ ) );
MUX2_X1 _15130_ ( .A(_07785_ ), .B(\ICACHE.cache_reg[0][25] ), .S(_07767_ ), .Z(_00301_ ) );
OAI211_X1 _15131_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_7_B_$_MUX__Y_A ), .B(_04090_ ), .C1(_04075_ ), .C2(_04099_ ), .ZN(_07786_ ) );
OAI21_X1 _15132_ ( .A(_07786_ ), .B1(_07729_ ), .B2(\io_master_rdata [24] ), .ZN(_07787_ ) );
NOR2_X1 _15133_ ( .A1(_07787_ ), .A2(_07543_ ), .ZN(_07788_ ) );
MUX2_X1 _15134_ ( .A(_07788_ ), .B(\ICACHE.cache_reg[0][24] ), .S(_07767_ ), .Z(_00302_ ) );
OAI211_X1 _15135_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_8_B_$_MUX__Y_A ), .B(_07698_ ), .C1(_07703_ ), .C2(_07704_ ), .ZN(_07789_ ) );
OAI21_X1 _15136_ ( .A(_07789_ ), .B1(_07700_ ), .B2(\io_master_rdata [23] ), .ZN(_07790_ ) );
NOR2_X1 _15137_ ( .A1(_07790_ ), .A2(_07543_ ), .ZN(_07791_ ) );
MUX2_X1 _15138_ ( .A(_07791_ ), .B(\ICACHE.cache_reg[0][23] ), .S(_07767_ ), .Z(_00303_ ) );
OAI211_X1 _15139_ ( .A(\ICACHE.s_axi_rdata_$_ANDNOT__Y_9_B_$_MUX__Y_A ), .B(_04091_ ), .C1(_07703_ ), .C2(_07704_ ), .ZN(_07792_ ) );
OAI21_X1 _15140_ ( .A(_07792_ ), .B1(_07706_ ), .B2(\io_master_rdata [22] ), .ZN(_07793_ ) );
NOR2_X1 _15141_ ( .A1(_07793_ ), .A2(_07543_ ), .ZN(_07794_ ) );
MUX2_X1 _15142_ ( .A(_07794_ ), .B(\ICACHE.cache_reg[0][22] ), .S(_07767_ ), .Z(_00304_ ) );
NAND3_X1 _15143_ ( .A1(_07544_ ), .A2(_07690_ ), .A3(_07695_ ), .ZN(_07795_ ) );
NAND2_X1 _15144_ ( .A1(_07601_ ), .A2(_03805_ ), .ZN(_07796_ ) );
NOR2_X1 _15145_ ( .A1(_07795_ ), .A2(_07796_ ), .ZN(_07797_ ) );
BUF_X4 _15146_ ( .A(_07797_ ), .Z(_07798_ ) );
MUX2_X1 _15147_ ( .A(\ICACHE.cache_reg[1][31] ), .B(_07689_ ), .S(_07798_ ), .Z(_00305_ ) );
MUX2_X1 _15148_ ( .A(\ICACHE.cache_reg[1][30] ), .B(_07702_ ), .S(_07798_ ), .Z(_00306_ ) );
MUX2_X1 _15149_ ( .A(\ICACHE.cache_reg[1][21] ), .B(_07708_ ), .S(_07798_ ), .Z(_00307_ ) );
MUX2_X1 _15150_ ( .A(\ICACHE.cache_reg[1][20] ), .B(_07711_ ), .S(_07798_ ), .Z(_00308_ ) );
MUX2_X1 _15151_ ( .A(\ICACHE.cache_reg[1][19] ), .B(_07714_ ), .S(_07798_ ), .Z(_00309_ ) );
MUX2_X1 _15152_ ( .A(\ICACHE.cache_reg[1][18] ), .B(_07717_ ), .S(_07798_ ), .Z(_00310_ ) );
MUX2_X1 _15153_ ( .A(\ICACHE.cache_reg[1][17] ), .B(_07721_ ), .S(_07798_ ), .Z(_00311_ ) );
MUX2_X1 _15154_ ( .A(\ICACHE.cache_reg[1][16] ), .B(_07724_ ), .S(_07798_ ), .Z(_00312_ ) );
MUX2_X1 _15155_ ( .A(\ICACHE.cache_reg[1][15] ), .B(_07727_ ), .S(_07798_ ), .Z(_00313_ ) );
MUX2_X1 _15156_ ( .A(\ICACHE.cache_reg[1][14] ), .B(_07731_ ), .S(_07798_ ), .Z(_00314_ ) );
BUF_X4 _15157_ ( .A(_07797_ ), .Z(_07799_ ) );
MUX2_X1 _15158_ ( .A(\ICACHE.cache_reg[1][13] ), .B(_07734_ ), .S(_07799_ ), .Z(_00315_ ) );
MUX2_X1 _15159_ ( .A(\ICACHE.cache_reg[1][12] ), .B(_07738_ ), .S(_07799_ ), .Z(_00316_ ) );
MUX2_X1 _15160_ ( .A(\ICACHE.cache_reg[1][29] ), .B(_07741_ ), .S(_07799_ ), .Z(_00317_ ) );
MUX2_X1 _15161_ ( .A(\ICACHE.cache_reg[1][11] ), .B(_07744_ ), .S(_07799_ ), .Z(_00318_ ) );
MUX2_X1 _15162_ ( .A(\ICACHE.cache_reg[1][10] ), .B(_07747_ ), .S(_07799_ ), .Z(_00319_ ) );
MUX2_X1 _15163_ ( .A(\ICACHE.cache_reg[1][9] ), .B(_07750_ ), .S(_07799_ ), .Z(_00320_ ) );
MUX2_X1 _15164_ ( .A(\ICACHE.cache_reg[1][8] ), .B(_07754_ ), .S(_07799_ ), .Z(_00321_ ) );
MUX2_X1 _15165_ ( .A(\ICACHE.cache_reg[1][7] ), .B(_07757_ ), .S(_07799_ ), .Z(_00322_ ) );
MUX2_X1 _15166_ ( .A(\ICACHE.cache_reg[1][6] ), .B(_07760_ ), .S(_07799_ ), .Z(_00323_ ) );
MUX2_X1 _15167_ ( .A(\ICACHE.cache_reg[1][5] ), .B(_07763_ ), .S(_07799_ ), .Z(_00324_ ) );
BUF_X4 _15168_ ( .A(_07797_ ), .Z(_07800_ ) );
MUX2_X1 _15169_ ( .A(\ICACHE.cache_reg[1][4] ), .B(_07766_ ), .S(_07800_ ), .Z(_00325_ ) );
MUX2_X1 _15170_ ( .A(\ICACHE.cache_reg[1][3] ), .B(_07770_ ), .S(_07800_ ), .Z(_00326_ ) );
MUX2_X1 _15171_ ( .A(\ICACHE.cache_reg[1][2] ), .B(_07773_ ), .S(_07800_ ), .Z(_00327_ ) );
MUX2_X1 _15172_ ( .A(\ICACHE.cache_reg[1][28] ), .B(_07776_ ), .S(_07800_ ), .Z(_00328_ ) );
MUX2_X1 _15173_ ( .A(\ICACHE.cache_reg[1][27] ), .B(_07779_ ), .S(_07800_ ), .Z(_00329_ ) );
MUX2_X1 _15174_ ( .A(\ICACHE.cache_reg[1][26] ), .B(_07782_ ), .S(_07800_ ), .Z(_00330_ ) );
MUX2_X1 _15175_ ( .A(\ICACHE.cache_reg[1][25] ), .B(_07785_ ), .S(_07800_ ), .Z(_00331_ ) );
MUX2_X1 _15176_ ( .A(\ICACHE.cache_reg[1][24] ), .B(_07788_ ), .S(_07800_ ), .Z(_00332_ ) );
MUX2_X1 _15177_ ( .A(\ICACHE.cache_reg[1][23] ), .B(_07791_ ), .S(_07800_ ), .Z(_00333_ ) );
MUX2_X1 _15178_ ( .A(\ICACHE.cache_reg[1][22] ), .B(_07794_ ), .S(_07800_ ), .Z(_00334_ ) );
NAND2_X1 _15179_ ( .A1(_07694_ ), .A2(_07533_ ), .ZN(_07801_ ) );
BUF_X4 _15180_ ( .A(_07801_ ), .Z(_07802_ ) );
MUX2_X1 _15181_ ( .A(_07689_ ), .B(\ICACHE.cache_reg[2][31] ), .S(_07802_ ), .Z(_00335_ ) );
MUX2_X1 _15182_ ( .A(_07702_ ), .B(\ICACHE.cache_reg[2][30] ), .S(_07802_ ), .Z(_00336_ ) );
MUX2_X1 _15183_ ( .A(_07708_ ), .B(\ICACHE.cache_reg[2][21] ), .S(_07802_ ), .Z(_00337_ ) );
MUX2_X1 _15184_ ( .A(_07711_ ), .B(\ICACHE.cache_reg[2][20] ), .S(_07802_ ), .Z(_00338_ ) );
MUX2_X1 _15185_ ( .A(_07714_ ), .B(\ICACHE.cache_reg[2][19] ), .S(_07802_ ), .Z(_00339_ ) );
MUX2_X1 _15186_ ( .A(_07717_ ), .B(\ICACHE.cache_reg[2][18] ), .S(_07802_ ), .Z(_00340_ ) );
MUX2_X1 _15187_ ( .A(_07721_ ), .B(\ICACHE.cache_reg[2][17] ), .S(_07802_ ), .Z(_00341_ ) );
MUX2_X1 _15188_ ( .A(_07724_ ), .B(\ICACHE.cache_reg[2][16] ), .S(_07802_ ), .Z(_00342_ ) );
MUX2_X1 _15189_ ( .A(_07727_ ), .B(\ICACHE.cache_reg[2][15] ), .S(_07802_ ), .Z(_00343_ ) );
MUX2_X1 _15190_ ( .A(_07731_ ), .B(\ICACHE.cache_reg[2][14] ), .S(_07802_ ), .Z(_00344_ ) );
BUF_X4 _15191_ ( .A(_07801_ ), .Z(_07803_ ) );
MUX2_X1 _15192_ ( .A(_07734_ ), .B(\ICACHE.cache_reg[2][13] ), .S(_07803_ ), .Z(_00345_ ) );
MUX2_X1 _15193_ ( .A(_07738_ ), .B(\ICACHE.cache_reg[2][12] ), .S(_07803_ ), .Z(_00346_ ) );
MUX2_X1 _15194_ ( .A(_07741_ ), .B(\ICACHE.cache_reg[2][29] ), .S(_07803_ ), .Z(_00347_ ) );
MUX2_X1 _15195_ ( .A(_07744_ ), .B(\ICACHE.cache_reg[2][11] ), .S(_07803_ ), .Z(_00348_ ) );
MUX2_X1 _15196_ ( .A(_07747_ ), .B(\ICACHE.cache_reg[2][10] ), .S(_07803_ ), .Z(_00349_ ) );
MUX2_X1 _15197_ ( .A(_07750_ ), .B(\ICACHE.cache_reg[2][9] ), .S(_07803_ ), .Z(_00350_ ) );
MUX2_X1 _15198_ ( .A(_07754_ ), .B(\ICACHE.cache_reg[2][8] ), .S(_07803_ ), .Z(_00351_ ) );
MUX2_X1 _15199_ ( .A(_07757_ ), .B(\ICACHE.cache_reg[2][7] ), .S(_07803_ ), .Z(_00352_ ) );
MUX2_X1 _15200_ ( .A(_07760_ ), .B(\ICACHE.cache_reg[2][6] ), .S(_07803_ ), .Z(_00353_ ) );
MUX2_X1 _15201_ ( .A(_07763_ ), .B(\ICACHE.cache_reg[2][5] ), .S(_07803_ ), .Z(_00354_ ) );
BUF_X4 _15202_ ( .A(_07801_ ), .Z(_07804_ ) );
MUX2_X1 _15203_ ( .A(_07766_ ), .B(\ICACHE.cache_reg[2][4] ), .S(_07804_ ), .Z(_00355_ ) );
MUX2_X1 _15204_ ( .A(_07770_ ), .B(\ICACHE.cache_reg[2][3] ), .S(_07804_ ), .Z(_00356_ ) );
MUX2_X1 _15205_ ( .A(_07773_ ), .B(\ICACHE.cache_reg[2][2] ), .S(_07804_ ), .Z(_00357_ ) );
MUX2_X1 _15206_ ( .A(_07776_ ), .B(\ICACHE.cache_reg[2][28] ), .S(_07804_ ), .Z(_00358_ ) );
MUX2_X1 _15207_ ( .A(_07779_ ), .B(\ICACHE.cache_reg[2][27] ), .S(_07804_ ), .Z(_00359_ ) );
MUX2_X1 _15208_ ( .A(_07782_ ), .B(\ICACHE.cache_reg[2][26] ), .S(_07804_ ), .Z(_00360_ ) );
MUX2_X1 _15209_ ( .A(_07785_ ), .B(\ICACHE.cache_reg[2][25] ), .S(_07804_ ), .Z(_00361_ ) );
MUX2_X1 _15210_ ( .A(_07788_ ), .B(\ICACHE.cache_reg[2][24] ), .S(_07804_ ), .Z(_00362_ ) );
MUX2_X1 _15211_ ( .A(_07791_ ), .B(\ICACHE.cache_reg[2][23] ), .S(_07804_ ), .Z(_00363_ ) );
MUX2_X1 _15212_ ( .A(_07794_ ), .B(\ICACHE.cache_reg[2][22] ), .S(_07804_ ), .Z(_00364_ ) );
NAND3_X1 _15213_ ( .A1(_07544_ ), .A2(_07690_ ), .A3(_07533_ ), .ZN(_07805_ ) );
NOR2_X1 _15214_ ( .A1(_07805_ ), .A2(_07796_ ), .ZN(_07806_ ) );
BUF_X4 _15215_ ( .A(_07806_ ), .Z(_07807_ ) );
MUX2_X1 _15216_ ( .A(\ICACHE.cache_reg[3][31] ), .B(_07689_ ), .S(_07807_ ), .Z(_00365_ ) );
MUX2_X1 _15217_ ( .A(\ICACHE.cache_reg[3][30] ), .B(_07702_ ), .S(_07807_ ), .Z(_00366_ ) );
MUX2_X1 _15218_ ( .A(\ICACHE.cache_reg[3][21] ), .B(_07708_ ), .S(_07807_ ), .Z(_00367_ ) );
MUX2_X1 _15219_ ( .A(\ICACHE.cache_reg[3][20] ), .B(_07711_ ), .S(_07807_ ), .Z(_00368_ ) );
MUX2_X1 _15220_ ( .A(\ICACHE.cache_reg[3][19] ), .B(_07714_ ), .S(_07807_ ), .Z(_00369_ ) );
MUX2_X1 _15221_ ( .A(\ICACHE.cache_reg[3][18] ), .B(_07717_ ), .S(_07807_ ), .Z(_00370_ ) );
MUX2_X1 _15222_ ( .A(\ICACHE.cache_reg[3][17] ), .B(_07721_ ), .S(_07807_ ), .Z(_00371_ ) );
MUX2_X1 _15223_ ( .A(\ICACHE.cache_reg[3][16] ), .B(_07724_ ), .S(_07807_ ), .Z(_00372_ ) );
MUX2_X1 _15224_ ( .A(\ICACHE.cache_reg[3][15] ), .B(_07727_ ), .S(_07807_ ), .Z(_00373_ ) );
MUX2_X1 _15225_ ( .A(\ICACHE.cache_reg[3][14] ), .B(_07731_ ), .S(_07807_ ), .Z(_00374_ ) );
BUF_X4 _15226_ ( .A(_07806_ ), .Z(_07808_ ) );
MUX2_X1 _15227_ ( .A(\ICACHE.cache_reg[3][13] ), .B(_07734_ ), .S(_07808_ ), .Z(_00375_ ) );
MUX2_X1 _15228_ ( .A(\ICACHE.cache_reg[3][12] ), .B(_07738_ ), .S(_07808_ ), .Z(_00376_ ) );
MUX2_X1 _15229_ ( .A(\ICACHE.cache_reg[3][29] ), .B(_07741_ ), .S(_07808_ ), .Z(_00377_ ) );
MUX2_X1 _15230_ ( .A(\ICACHE.cache_reg[3][11] ), .B(_07744_ ), .S(_07808_ ), .Z(_00378_ ) );
MUX2_X1 _15231_ ( .A(\ICACHE.cache_reg[3][10] ), .B(_07747_ ), .S(_07808_ ), .Z(_00379_ ) );
MUX2_X1 _15232_ ( .A(\ICACHE.cache_reg[3][9] ), .B(_07750_ ), .S(_07808_ ), .Z(_00380_ ) );
MUX2_X1 _15233_ ( .A(\ICACHE.cache_reg[3][8] ), .B(_07754_ ), .S(_07808_ ), .Z(_00381_ ) );
MUX2_X1 _15234_ ( .A(\ICACHE.cache_reg[3][7] ), .B(_07757_ ), .S(_07808_ ), .Z(_00382_ ) );
MUX2_X1 _15235_ ( .A(\ICACHE.cache_reg[3][6] ), .B(_07760_ ), .S(_07808_ ), .Z(_00383_ ) );
MUX2_X1 _15236_ ( .A(\ICACHE.cache_reg[3][5] ), .B(_07763_ ), .S(_07808_ ), .Z(_00384_ ) );
BUF_X4 _15237_ ( .A(_07806_ ), .Z(_07809_ ) );
MUX2_X1 _15238_ ( .A(\ICACHE.cache_reg[3][4] ), .B(_07766_ ), .S(_07809_ ), .Z(_00385_ ) );
MUX2_X1 _15239_ ( .A(\ICACHE.cache_reg[3][3] ), .B(_07770_ ), .S(_07809_ ), .Z(_00386_ ) );
MUX2_X1 _15240_ ( .A(\ICACHE.cache_reg[3][2] ), .B(_07773_ ), .S(_07809_ ), .Z(_00387_ ) );
MUX2_X1 _15241_ ( .A(\ICACHE.cache_reg[3][28] ), .B(_07776_ ), .S(_07809_ ), .Z(_00388_ ) );
MUX2_X1 _15242_ ( .A(\ICACHE.cache_reg[3][27] ), .B(_07779_ ), .S(_07809_ ), .Z(_00389_ ) );
MUX2_X1 _15243_ ( .A(\ICACHE.cache_reg[3][26] ), .B(_07782_ ), .S(_07809_ ), .Z(_00390_ ) );
MUX2_X1 _15244_ ( .A(\ICACHE.cache_reg[3][25] ), .B(_07785_ ), .S(_07809_ ), .Z(_00391_ ) );
MUX2_X1 _15245_ ( .A(\ICACHE.cache_reg[3][24] ), .B(_07788_ ), .S(_07809_ ), .Z(_00392_ ) );
MUX2_X1 _15246_ ( .A(\ICACHE.cache_reg[3][23] ), .B(_07791_ ), .S(_07809_ ), .Z(_00393_ ) );
MUX2_X1 _15247_ ( .A(\ICACHE.cache_reg[3][22] ), .B(_07794_ ), .S(_07809_ ), .Z(_00394_ ) );
AND2_X2 _15248_ ( .A1(_07694_ ), .A2(_07532_ ), .ZN(_07810_ ) );
BUF_X4 _15249_ ( .A(_07810_ ), .Z(_07811_ ) );
MUX2_X1 _15250_ ( .A(\ICACHE.cache_reg[4][31] ), .B(_07689_ ), .S(_07811_ ), .Z(_00395_ ) );
MUX2_X1 _15251_ ( .A(\ICACHE.cache_reg[4][30] ), .B(_07702_ ), .S(_07811_ ), .Z(_00396_ ) );
MUX2_X1 _15252_ ( .A(\ICACHE.cache_reg[4][21] ), .B(_07708_ ), .S(_07811_ ), .Z(_00397_ ) );
MUX2_X1 _15253_ ( .A(\ICACHE.cache_reg[4][20] ), .B(_07711_ ), .S(_07811_ ), .Z(_00398_ ) );
MUX2_X1 _15254_ ( .A(\ICACHE.cache_reg[4][19] ), .B(_07714_ ), .S(_07811_ ), .Z(_00399_ ) );
MUX2_X1 _15255_ ( .A(\ICACHE.cache_reg[4][18] ), .B(_07717_ ), .S(_07811_ ), .Z(_00400_ ) );
MUX2_X1 _15256_ ( .A(\ICACHE.cache_reg[4][17] ), .B(_07721_ ), .S(_07811_ ), .Z(_00401_ ) );
MUX2_X1 _15257_ ( .A(\ICACHE.cache_reg[4][16] ), .B(_07724_ ), .S(_07811_ ), .Z(_00402_ ) );
MUX2_X1 _15258_ ( .A(\ICACHE.cache_reg[4][15] ), .B(_07727_ ), .S(_07811_ ), .Z(_00403_ ) );
MUX2_X1 _15259_ ( .A(\ICACHE.cache_reg[4][14] ), .B(_07731_ ), .S(_07811_ ), .Z(_00404_ ) );
BUF_X4 _15260_ ( .A(_07810_ ), .Z(_07812_ ) );
MUX2_X1 _15261_ ( .A(\ICACHE.cache_reg[4][13] ), .B(_07734_ ), .S(_07812_ ), .Z(_00405_ ) );
MUX2_X1 _15262_ ( .A(\ICACHE.cache_reg[4][12] ), .B(_07738_ ), .S(_07812_ ), .Z(_00406_ ) );
MUX2_X1 _15263_ ( .A(\ICACHE.cache_reg[4][29] ), .B(_07741_ ), .S(_07812_ ), .Z(_00407_ ) );
MUX2_X1 _15264_ ( .A(\ICACHE.cache_reg[4][11] ), .B(_07744_ ), .S(_07812_ ), .Z(_00408_ ) );
MUX2_X1 _15265_ ( .A(\ICACHE.cache_reg[4][10] ), .B(_07747_ ), .S(_07812_ ), .Z(_00409_ ) );
MUX2_X1 _15266_ ( .A(\ICACHE.cache_reg[4][9] ), .B(_07750_ ), .S(_07812_ ), .Z(_00410_ ) );
MUX2_X1 _15267_ ( .A(\ICACHE.cache_reg[4][8] ), .B(_07754_ ), .S(_07812_ ), .Z(_00411_ ) );
MUX2_X1 _15268_ ( .A(\ICACHE.cache_reg[4][7] ), .B(_07757_ ), .S(_07812_ ), .Z(_00412_ ) );
MUX2_X1 _15269_ ( .A(\ICACHE.cache_reg[4][6] ), .B(_07760_ ), .S(_07812_ ), .Z(_00413_ ) );
MUX2_X1 _15270_ ( .A(\ICACHE.cache_reg[4][5] ), .B(_07763_ ), .S(_07812_ ), .Z(_00414_ ) );
BUF_X4 _15271_ ( .A(_07810_ ), .Z(_07813_ ) );
MUX2_X1 _15272_ ( .A(\ICACHE.cache_reg[4][4] ), .B(_07766_ ), .S(_07813_ ), .Z(_00415_ ) );
MUX2_X1 _15273_ ( .A(\ICACHE.cache_reg[4][3] ), .B(_07770_ ), .S(_07813_ ), .Z(_00416_ ) );
MUX2_X1 _15274_ ( .A(\ICACHE.cache_reg[4][2] ), .B(_07773_ ), .S(_07813_ ), .Z(_00417_ ) );
MUX2_X1 _15275_ ( .A(\ICACHE.cache_reg[4][28] ), .B(_07776_ ), .S(_07813_ ), .Z(_00418_ ) );
MUX2_X1 _15276_ ( .A(\ICACHE.cache_reg[4][27] ), .B(_07779_ ), .S(_07813_ ), .Z(_00419_ ) );
MUX2_X1 _15277_ ( .A(\ICACHE.cache_reg[4][26] ), .B(_07782_ ), .S(_07813_ ), .Z(_00420_ ) );
MUX2_X1 _15278_ ( .A(\ICACHE.cache_reg[4][25] ), .B(_07785_ ), .S(_07813_ ), .Z(_00421_ ) );
MUX2_X1 _15279_ ( .A(\ICACHE.cache_reg[4][24] ), .B(_07788_ ), .S(_07813_ ), .Z(_00422_ ) );
MUX2_X1 _15280_ ( .A(\ICACHE.cache_reg[4][23] ), .B(_07791_ ), .S(_07813_ ), .Z(_00423_ ) );
MUX2_X1 _15281_ ( .A(\ICACHE.cache_reg[4][22] ), .B(_07794_ ), .S(_07813_ ), .Z(_00424_ ) );
NAND3_X1 _15282_ ( .A1(_07544_ ), .A2(_07690_ ), .A3(_07532_ ), .ZN(_07814_ ) );
OR2_X2 _15283_ ( .A1(_07814_ ), .A2(_07796_ ), .ZN(_07815_ ) );
BUF_X4 _15284_ ( .A(_07815_ ), .Z(_07816_ ) );
MUX2_X1 _15285_ ( .A(_07689_ ), .B(\ICACHE.cache_reg[5][31] ), .S(_07816_ ), .Z(_00425_ ) );
MUX2_X1 _15286_ ( .A(_07702_ ), .B(\ICACHE.cache_reg[5][30] ), .S(_07816_ ), .Z(_00426_ ) );
MUX2_X1 _15287_ ( .A(_07708_ ), .B(\ICACHE.cache_reg[5][21] ), .S(_07816_ ), .Z(_00427_ ) );
MUX2_X1 _15288_ ( .A(_07711_ ), .B(\ICACHE.cache_reg[5][20] ), .S(_07816_ ), .Z(_00428_ ) );
MUX2_X1 _15289_ ( .A(_07714_ ), .B(\ICACHE.cache_reg[5][19] ), .S(_07816_ ), .Z(_00429_ ) );
MUX2_X1 _15290_ ( .A(_07717_ ), .B(\ICACHE.cache_reg[5][18] ), .S(_07816_ ), .Z(_00430_ ) );
MUX2_X1 _15291_ ( .A(_07721_ ), .B(\ICACHE.cache_reg[5][17] ), .S(_07816_ ), .Z(_00431_ ) );
MUX2_X1 _15292_ ( .A(_07724_ ), .B(\ICACHE.cache_reg[5][16] ), .S(_07816_ ), .Z(_00432_ ) );
MUX2_X1 _15293_ ( .A(_07727_ ), .B(\ICACHE.cache_reg[5][15] ), .S(_07816_ ), .Z(_00433_ ) );
MUX2_X1 _15294_ ( .A(_07731_ ), .B(\ICACHE.cache_reg[5][14] ), .S(_07816_ ), .Z(_00434_ ) );
BUF_X4 _15295_ ( .A(_07815_ ), .Z(_07817_ ) );
MUX2_X1 _15296_ ( .A(_07734_ ), .B(\ICACHE.cache_reg[5][13] ), .S(_07817_ ), .Z(_00435_ ) );
MUX2_X1 _15297_ ( .A(_07738_ ), .B(\ICACHE.cache_reg[5][12] ), .S(_07817_ ), .Z(_00436_ ) );
MUX2_X1 _15298_ ( .A(_07741_ ), .B(\ICACHE.cache_reg[5][29] ), .S(_07817_ ), .Z(_00437_ ) );
MUX2_X1 _15299_ ( .A(_07744_ ), .B(\ICACHE.cache_reg[5][11] ), .S(_07817_ ), .Z(_00438_ ) );
MUX2_X1 _15300_ ( .A(_07747_ ), .B(\ICACHE.cache_reg[5][10] ), .S(_07817_ ), .Z(_00439_ ) );
MUX2_X1 _15301_ ( .A(_07750_ ), .B(\ICACHE.cache_reg[5][9] ), .S(_07817_ ), .Z(_00440_ ) );
MUX2_X1 _15302_ ( .A(_07754_ ), .B(\ICACHE.cache_reg[5][8] ), .S(_07817_ ), .Z(_00441_ ) );
MUX2_X1 _15303_ ( .A(_07757_ ), .B(\ICACHE.cache_reg[5][7] ), .S(_07817_ ), .Z(_00442_ ) );
MUX2_X1 _15304_ ( .A(_07760_ ), .B(\ICACHE.cache_reg[5][6] ), .S(_07817_ ), .Z(_00443_ ) );
MUX2_X1 _15305_ ( .A(_07763_ ), .B(\ICACHE.cache_reg[5][5] ), .S(_07817_ ), .Z(_00444_ ) );
BUF_X4 _15306_ ( .A(_07815_ ), .Z(_07818_ ) );
MUX2_X1 _15307_ ( .A(_07766_ ), .B(\ICACHE.cache_reg[5][4] ), .S(_07818_ ), .Z(_00445_ ) );
MUX2_X1 _15308_ ( .A(_07770_ ), .B(\ICACHE.cache_reg[5][3] ), .S(_07818_ ), .Z(_00446_ ) );
MUX2_X1 _15309_ ( .A(_07773_ ), .B(\ICACHE.cache_reg[5][2] ), .S(_07818_ ), .Z(_00447_ ) );
MUX2_X1 _15310_ ( .A(_07776_ ), .B(\ICACHE.cache_reg[5][28] ), .S(_07818_ ), .Z(_00448_ ) );
MUX2_X1 _15311_ ( .A(_07779_ ), .B(\ICACHE.cache_reg[5][27] ), .S(_07818_ ), .Z(_00449_ ) );
MUX2_X1 _15312_ ( .A(_07782_ ), .B(\ICACHE.cache_reg[5][26] ), .S(_07818_ ), .Z(_00450_ ) );
MUX2_X1 _15313_ ( .A(_07785_ ), .B(\ICACHE.cache_reg[5][25] ), .S(_07818_ ), .Z(_00451_ ) );
MUX2_X1 _15314_ ( .A(_07788_ ), .B(\ICACHE.cache_reg[5][24] ), .S(_07818_ ), .Z(_00452_ ) );
MUX2_X1 _15315_ ( .A(_07791_ ), .B(\ICACHE.cache_reg[5][23] ), .S(_07818_ ), .Z(_00453_ ) );
MUX2_X1 _15316_ ( .A(_07794_ ), .B(\ICACHE.cache_reg[5][22] ), .S(_07818_ ), .Z(_00454_ ) );
AND2_X1 _15317_ ( .A1(\ICACHE.burst_counter [1] ), .A2(\ICACHE.burst_counter [0] ), .ZN(_07819_ ) );
NAND2_X1 _15318_ ( .A1(_07694_ ), .A2(_07819_ ), .ZN(_07820_ ) );
BUF_X4 _15319_ ( .A(_07820_ ), .Z(_07821_ ) );
MUX2_X1 _15320_ ( .A(_07689_ ), .B(\ICACHE.cache_reg[6][31] ), .S(_07821_ ), .Z(_00455_ ) );
MUX2_X1 _15321_ ( .A(_07702_ ), .B(\ICACHE.cache_reg[6][30] ), .S(_07821_ ), .Z(_00456_ ) );
MUX2_X1 _15322_ ( .A(_07708_ ), .B(\ICACHE.cache_reg[6][21] ), .S(_07821_ ), .Z(_00457_ ) );
MUX2_X1 _15323_ ( .A(_07711_ ), .B(\ICACHE.cache_reg[6][20] ), .S(_07821_ ), .Z(_00458_ ) );
MUX2_X1 _15324_ ( .A(_07714_ ), .B(\ICACHE.cache_reg[6][19] ), .S(_07821_ ), .Z(_00459_ ) );
MUX2_X1 _15325_ ( .A(_07717_ ), .B(\ICACHE.cache_reg[6][18] ), .S(_07821_ ), .Z(_00460_ ) );
MUX2_X1 _15326_ ( .A(_07721_ ), .B(\ICACHE.cache_reg[6][17] ), .S(_07821_ ), .Z(_00461_ ) );
MUX2_X1 _15327_ ( .A(_07724_ ), .B(\ICACHE.cache_reg[6][16] ), .S(_07821_ ), .Z(_00462_ ) );
MUX2_X1 _15328_ ( .A(_07727_ ), .B(\ICACHE.cache_reg[6][15] ), .S(_07821_ ), .Z(_00463_ ) );
MUX2_X1 _15329_ ( .A(_07731_ ), .B(\ICACHE.cache_reg[6][14] ), .S(_07821_ ), .Z(_00464_ ) );
BUF_X4 _15330_ ( .A(_07820_ ), .Z(_07822_ ) );
MUX2_X1 _15331_ ( .A(_07734_ ), .B(\ICACHE.cache_reg[6][13] ), .S(_07822_ ), .Z(_00465_ ) );
MUX2_X1 _15332_ ( .A(_07738_ ), .B(\ICACHE.cache_reg[6][12] ), .S(_07822_ ), .Z(_00466_ ) );
MUX2_X1 _15333_ ( .A(_07741_ ), .B(\ICACHE.cache_reg[6][29] ), .S(_07822_ ), .Z(_00467_ ) );
MUX2_X1 _15334_ ( .A(_07744_ ), .B(\ICACHE.cache_reg[6][11] ), .S(_07822_ ), .Z(_00468_ ) );
MUX2_X1 _15335_ ( .A(_07747_ ), .B(\ICACHE.cache_reg[6][10] ), .S(_07822_ ), .Z(_00469_ ) );
MUX2_X1 _15336_ ( .A(_07750_ ), .B(\ICACHE.cache_reg[6][9] ), .S(_07822_ ), .Z(_00470_ ) );
MUX2_X1 _15337_ ( .A(_07754_ ), .B(\ICACHE.cache_reg[6][8] ), .S(_07822_ ), .Z(_00471_ ) );
MUX2_X1 _15338_ ( .A(_07757_ ), .B(\ICACHE.cache_reg[6][7] ), .S(_07822_ ), .Z(_00472_ ) );
MUX2_X1 _15339_ ( .A(_07760_ ), .B(\ICACHE.cache_reg[6][6] ), .S(_07822_ ), .Z(_00473_ ) );
MUX2_X1 _15340_ ( .A(_07763_ ), .B(\ICACHE.cache_reg[6][5] ), .S(_07822_ ), .Z(_00474_ ) );
BUF_X4 _15341_ ( .A(_07820_ ), .Z(_07823_ ) );
MUX2_X1 _15342_ ( .A(_07766_ ), .B(\ICACHE.cache_reg[6][4] ), .S(_07823_ ), .Z(_00475_ ) );
MUX2_X1 _15343_ ( .A(_07770_ ), .B(\ICACHE.cache_reg[6][3] ), .S(_07823_ ), .Z(_00476_ ) );
MUX2_X1 _15344_ ( .A(_07773_ ), .B(\ICACHE.cache_reg[6][2] ), .S(_07823_ ), .Z(_00477_ ) );
MUX2_X1 _15345_ ( .A(_07776_ ), .B(\ICACHE.cache_reg[6][28] ), .S(_07823_ ), .Z(_00478_ ) );
MUX2_X1 _15346_ ( .A(_07779_ ), .B(\ICACHE.cache_reg[6][27] ), .S(_07823_ ), .Z(_00479_ ) );
MUX2_X1 _15347_ ( .A(_07782_ ), .B(\ICACHE.cache_reg[6][26] ), .S(_07823_ ), .Z(_00480_ ) );
MUX2_X1 _15348_ ( .A(_07785_ ), .B(\ICACHE.cache_reg[6][25] ), .S(_07823_ ), .Z(_00481_ ) );
MUX2_X1 _15349_ ( .A(_07788_ ), .B(\ICACHE.cache_reg[6][24] ), .S(_07823_ ), .Z(_00482_ ) );
MUX2_X1 _15350_ ( .A(_07791_ ), .B(\ICACHE.cache_reg[6][23] ), .S(_07823_ ), .Z(_00483_ ) );
MUX2_X1 _15351_ ( .A(_07794_ ), .B(\ICACHE.cache_reg[6][22] ), .S(_07823_ ), .Z(_00484_ ) );
NAND3_X1 _15352_ ( .A1(_07544_ ), .A2(_07690_ ), .A3(_07819_ ), .ZN(_07824_ ) );
NOR2_X1 _15353_ ( .A1(_07824_ ), .A2(_07796_ ), .ZN(_07825_ ) );
BUF_X4 _15354_ ( .A(_07825_ ), .Z(_07826_ ) );
MUX2_X1 _15355_ ( .A(\ICACHE.cache_reg[7][31] ), .B(_07689_ ), .S(_07826_ ), .Z(_00485_ ) );
MUX2_X1 _15356_ ( .A(\ICACHE.cache_reg[7][30] ), .B(_07702_ ), .S(_07826_ ), .Z(_00486_ ) );
MUX2_X1 _15357_ ( .A(\ICACHE.cache_reg[7][21] ), .B(_07708_ ), .S(_07826_ ), .Z(_00487_ ) );
MUX2_X1 _15358_ ( .A(\ICACHE.cache_reg[7][20] ), .B(_07711_ ), .S(_07826_ ), .Z(_00488_ ) );
MUX2_X1 _15359_ ( .A(\ICACHE.cache_reg[7][19] ), .B(_07714_ ), .S(_07826_ ), .Z(_00489_ ) );
MUX2_X1 _15360_ ( .A(\ICACHE.cache_reg[7][18] ), .B(_07717_ ), .S(_07826_ ), .Z(_00490_ ) );
MUX2_X1 _15361_ ( .A(\ICACHE.cache_reg[7][17] ), .B(_07721_ ), .S(_07826_ ), .Z(_00491_ ) );
MUX2_X1 _15362_ ( .A(\ICACHE.cache_reg[7][16] ), .B(_07724_ ), .S(_07826_ ), .Z(_00492_ ) );
MUX2_X1 _15363_ ( .A(\ICACHE.cache_reg[7][15] ), .B(_07727_ ), .S(_07826_ ), .Z(_00493_ ) );
MUX2_X1 _15364_ ( .A(\ICACHE.cache_reg[7][14] ), .B(_07731_ ), .S(_07826_ ), .Z(_00494_ ) );
BUF_X4 _15365_ ( .A(_07825_ ), .Z(_07827_ ) );
MUX2_X1 _15366_ ( .A(\ICACHE.cache_reg[7][13] ), .B(_07734_ ), .S(_07827_ ), .Z(_00495_ ) );
MUX2_X1 _15367_ ( .A(\ICACHE.cache_reg[7][12] ), .B(_07738_ ), .S(_07827_ ), .Z(_00496_ ) );
MUX2_X1 _15368_ ( .A(\ICACHE.cache_reg[7][29] ), .B(_07741_ ), .S(_07827_ ), .Z(_00497_ ) );
MUX2_X1 _15369_ ( .A(\ICACHE.cache_reg[7][11] ), .B(_07744_ ), .S(_07827_ ), .Z(_00498_ ) );
MUX2_X1 _15370_ ( .A(\ICACHE.cache_reg[7][10] ), .B(_07747_ ), .S(_07827_ ), .Z(_00499_ ) );
MUX2_X1 _15371_ ( .A(\ICACHE.cache_reg[7][9] ), .B(_07750_ ), .S(_07827_ ), .Z(_00500_ ) );
MUX2_X1 _15372_ ( .A(\ICACHE.cache_reg[7][8] ), .B(_07754_ ), .S(_07827_ ), .Z(_00501_ ) );
MUX2_X1 _15373_ ( .A(\ICACHE.cache_reg[7][7] ), .B(_07757_ ), .S(_07827_ ), .Z(_00502_ ) );
MUX2_X1 _15374_ ( .A(\ICACHE.cache_reg[7][6] ), .B(_07760_ ), .S(_07827_ ), .Z(_00503_ ) );
MUX2_X1 _15375_ ( .A(\ICACHE.cache_reg[7][5] ), .B(_07763_ ), .S(_07827_ ), .Z(_00504_ ) );
BUF_X4 _15376_ ( .A(_07825_ ), .Z(_07828_ ) );
MUX2_X1 _15377_ ( .A(\ICACHE.cache_reg[7][4] ), .B(_07766_ ), .S(_07828_ ), .Z(_00505_ ) );
MUX2_X1 _15378_ ( .A(\ICACHE.cache_reg[7][3] ), .B(_07770_ ), .S(_07828_ ), .Z(_00506_ ) );
MUX2_X1 _15379_ ( .A(\ICACHE.cache_reg[7][2] ), .B(_07773_ ), .S(_07828_ ), .Z(_00507_ ) );
MUX2_X1 _15380_ ( .A(\ICACHE.cache_reg[7][28] ), .B(_07776_ ), .S(_07828_ ), .Z(_00508_ ) );
MUX2_X1 _15381_ ( .A(\ICACHE.cache_reg[7][27] ), .B(_07779_ ), .S(_07828_ ), .Z(_00509_ ) );
MUX2_X1 _15382_ ( .A(\ICACHE.cache_reg[7][26] ), .B(_07782_ ), .S(_07828_ ), .Z(_00510_ ) );
MUX2_X1 _15383_ ( .A(\ICACHE.cache_reg[7][25] ), .B(_07785_ ), .S(_07828_ ), .Z(_00511_ ) );
MUX2_X1 _15384_ ( .A(\ICACHE.cache_reg[7][24] ), .B(_07788_ ), .S(_07828_ ), .Z(_00512_ ) );
MUX2_X1 _15385_ ( .A(\ICACHE.cache_reg[7][23] ), .B(_07791_ ), .S(_07828_ ), .Z(_00513_ ) );
MUX2_X1 _15386_ ( .A(\ICACHE.cache_reg[7][22] ), .B(_07794_ ), .S(_07828_ ), .Z(_00514_ ) );
NOR2_X2 _15387_ ( .A1(fanout_net_11 ), .A2(\ICACHE.s_axi_rready ), .ZN(_07829_ ) );
BUF_X4 _15388_ ( .A(_07829_ ), .Z(_07830_ ) );
MUX2_X1 _15389_ ( .A(\ICACHE.s_axi_araddr [31] ), .B(\BTB.pc_i [31] ), .S(_07830_ ), .Z(_00529_ ) );
MUX2_X1 _15390_ ( .A(\ICACHE.s_axi_araddr [30] ), .B(\BTB.pc_i [30] ), .S(_07830_ ), .Z(_00530_ ) );
MUX2_X1 _15391_ ( .A(\ICACHE.s_axi_araddr [21] ), .B(\BTB.pc_i [21] ), .S(_07830_ ), .Z(_00531_ ) );
MUX2_X1 _15392_ ( .A(\ICACHE.s_axi_araddr [20] ), .B(\BTB.pc_i [20] ), .S(_07830_ ), .Z(_00532_ ) );
MUX2_X1 _15393_ ( .A(\ICACHE.s_axi_araddr [19] ), .B(\BTB.pc_i [19] ), .S(_07830_ ), .Z(_00533_ ) );
MUX2_X1 _15394_ ( .A(\ICACHE.s_axi_araddr [18] ), .B(\BTB.pc_i [18] ), .S(_07830_ ), .Z(_00534_ ) );
MUX2_X1 _15395_ ( .A(\ICACHE.s_axi_araddr [17] ), .B(\BTB.pc_i [17] ), .S(_07830_ ), .Z(_00535_ ) );
MUX2_X1 _15396_ ( .A(\ICACHE.s_axi_araddr [16] ), .B(\BTB.pc_i [16] ), .S(_07830_ ), .Z(_00536_ ) );
MUX2_X1 _15397_ ( .A(\ICACHE.s_axi_araddr [1] ), .B(\BTB.pc_i [1] ), .S(_07830_ ), .Z(_00537_ ) );
MUX2_X1 _15398_ ( .A(\ICACHE.s_axi_araddr [0] ), .B(\BTB.pc_i [0] ), .S(_07830_ ), .Z(_00538_ ) );
MUX2_X1 _15399_ ( .A(\ICACHE.s_axi_araddr [29] ), .B(\BTB.pc_i [29] ), .S(_07829_ ), .Z(_00539_ ) );
MUX2_X1 _15400_ ( .A(\ICACHE.s_axi_araddr [28] ), .B(\BTB.pc_i [28] ), .S(_07829_ ), .Z(_00540_ ) );
MUX2_X1 _15401_ ( .A(\ICACHE.s_axi_araddr [27] ), .B(\BTB.pc_i [27] ), .S(_07829_ ), .Z(_00541_ ) );
MUX2_X1 _15402_ ( .A(\ICACHE.s_axi_araddr [26] ), .B(\BTB.pc_i [26] ), .S(_07829_ ), .Z(_00542_ ) );
MUX2_X1 _15403_ ( .A(\ICACHE.s_axi_araddr [25] ), .B(\BTB.pc_i [25] ), .S(_07829_ ), .Z(_00543_ ) );
MUX2_X1 _15404_ ( .A(\ICACHE.s_axi_araddr [24] ), .B(\BTB.pc_i [24] ), .S(_07829_ ), .Z(_00544_ ) );
MUX2_X1 _15405_ ( .A(\ICACHE.s_axi_araddr [23] ), .B(\BTB.pc_i [23] ), .S(_07829_ ), .Z(_00545_ ) );
MUX2_X1 _15406_ ( .A(\ICACHE.s_axi_araddr [22] ), .B(\BTB.pc_i [22] ), .S(_07829_ ), .Z(_00546_ ) );
BUF_X4 _15407_ ( .A(_04105_ ), .Z(_07831_ ) );
AND3_X1 _15408_ ( .A1(_07540_ ), .A2(io_master_rlast ), .A3(_07831_ ), .ZN(_07832_ ) );
AOI21_X1 _15409_ ( .A(_07660_ ), .B1(_07832_ ), .B2(\ICACHE.s_axi_rready ), .ZN(_07833_ ) );
NOR2_X1 _15410_ ( .A1(_07684_ ), .A2(_07833_ ), .ZN(_07834_ ) );
INV_X1 _15411_ ( .A(\ICACHE.s_axi_arlen [3] ), .ZN(_07835_ ) );
NOR2_X1 _15412_ ( .A1(_07834_ ), .A2(_07835_ ), .ZN(_00547_ ) );
INV_X1 _15413_ ( .A(_07652_ ), .ZN(_07836_ ) );
BUF_X4 _15414_ ( .A(_07836_ ), .Z(_07837_ ) );
INV_X1 _15415_ ( .A(\BTB.pc_i [30] ), .ZN(_07838_ ) );
AND3_X1 _15416_ ( .A1(_07838_ ), .A2(\BTB.pc_i [31] ), .A3(\BTB.pc_i [29] ), .ZN(_07839_ ) );
AND3_X1 _15417_ ( .A1(_07837_ ), .A2(_07535_ ), .A3(_07839_ ), .ZN(_07840_ ) );
MUX2_X1 _15418_ ( .A(\ICACHE.s_axi_arlen [1] ), .B(_07840_ ), .S(_07834_ ), .Z(_00548_ ) );
BUF_X2 _15419_ ( .A(_07645_ ), .Z(_07841_ ) );
AND3_X1 _15420_ ( .A1(_07841_ ), .A2(_07535_ ), .A3(_07839_ ), .ZN(_07842_ ) );
MUX2_X1 _15421_ ( .A(\ICACHE.s_axi_arlen [0] ), .B(_07842_ ), .S(_07834_ ), .Z(_00549_ ) );
BUF_X4 _15422_ ( .A(_07660_ ), .Z(_07843_ ) );
BUF_X4 _15423_ ( .A(_07843_ ), .Z(_07844_ ) );
MUX2_X1 _15424_ ( .A(\ICACHE.tag_check [15] ), .B(\BTB.pc_i [31] ), .S(_07844_ ), .Z(_00552_ ) );
MUX2_X1 _15425_ ( .A(\ICACHE.tag_check [14] ), .B(\BTB.pc_i [30] ), .S(_07844_ ), .Z(_00553_ ) );
MUX2_X1 _15426_ ( .A(\ICACHE.tag_check [5] ), .B(\BTB.pc_i [21] ), .S(_07844_ ), .Z(_00554_ ) );
MUX2_X1 _15427_ ( .A(\ICACHE.tag_check [4] ), .B(\BTB.pc_i [20] ), .S(_07844_ ), .Z(_00555_ ) );
MUX2_X1 _15428_ ( .A(\ICACHE.tag_check [3] ), .B(\BTB.pc_i [19] ), .S(_07844_ ), .Z(_00556_ ) );
MUX2_X1 _15429_ ( .A(\ICACHE.tag_check [2] ), .B(\BTB.pc_i [18] ), .S(_07844_ ), .Z(_00557_ ) );
MUX2_X1 _15430_ ( .A(\ICACHE.tag_check [1] ), .B(\BTB.pc_i [17] ), .S(_07844_ ), .Z(_00558_ ) );
MUX2_X1 _15431_ ( .A(\ICACHE.tag_check [0] ), .B(\BTB.pc_i [16] ), .S(_07844_ ), .Z(_00559_ ) );
MUX2_X1 _15432_ ( .A(\ICACHE.tag_check [13] ), .B(\BTB.pc_i [29] ), .S(_07844_ ), .Z(_00560_ ) );
MUX2_X1 _15433_ ( .A(\ICACHE.tag_check [12] ), .B(\BTB.pc_i [28] ), .S(_07843_ ), .Z(_00561_ ) );
MUX2_X1 _15434_ ( .A(\ICACHE.tag_check [11] ), .B(\BTB.pc_i [27] ), .S(_07843_ ), .Z(_00562_ ) );
MUX2_X1 _15435_ ( .A(\ICACHE.tag_check [10] ), .B(\BTB.pc_i [26] ), .S(_07843_ ), .Z(_00563_ ) );
MUX2_X1 _15436_ ( .A(\ICACHE.tag_check [9] ), .B(\BTB.pc_i [25] ), .S(_07843_ ), .Z(_00564_ ) );
MUX2_X1 _15437_ ( .A(\ICACHE.tag_check [8] ), .B(\BTB.pc_i [24] ), .S(_07843_ ), .Z(_00565_ ) );
MUX2_X1 _15438_ ( .A(\ICACHE.tag_check [7] ), .B(\BTB.pc_i [23] ), .S(_07843_ ), .Z(_00566_ ) );
MUX2_X1 _15439_ ( .A(\ICACHE.tag_check [6] ), .B(\BTB.pc_i [22] ), .S(_07843_ ), .Z(_00567_ ) );
INV_X1 _15440_ ( .A(_07694_ ), .ZN(_07845_ ) );
BUF_X4 _15441_ ( .A(_07845_ ), .Z(_07846_ ) );
NAND3_X1 _15442_ ( .A1(_07846_ ), .A2(\ICACHE.tag_reg[0][10] ), .A3(_04045_ ), .ZN(_07847_ ) );
BUF_X4 _15443_ ( .A(_07845_ ), .Z(_07848_ ) );
OAI21_X1 _15444_ ( .A(_07847_ ), .B1(_07634_ ), .B2(_07848_ ), .ZN(_00568_ ) );
NAND3_X1 _15445_ ( .A1(_07846_ ), .A2(\ICACHE.tag_reg[0][9] ), .A3(_04045_ ), .ZN(_07849_ ) );
OAI21_X1 _15446_ ( .A(_07849_ ), .B1(_07584_ ), .B2(_07848_ ), .ZN(_00569_ ) );
BUF_X4 _15447_ ( .A(_03808_ ), .Z(_07850_ ) );
NAND3_X1 _15448_ ( .A1(_07846_ ), .A2(\ICACHE.tag_reg[0][0] ), .A3(_07850_ ), .ZN(_07851_ ) );
OAI21_X1 _15449_ ( .A(_07851_ ), .B1(_07605_ ), .B2(_07848_ ), .ZN(_00570_ ) );
NAND3_X1 _15450_ ( .A1(_07846_ ), .A2(\ICACHE.tag_reg[0][8] ), .A3(_07850_ ), .ZN(_07852_ ) );
OAI21_X1 _15451_ ( .A(_07852_ ), .B1(_07593_ ), .B2(_07848_ ), .ZN(_00571_ ) );
NAND3_X1 _15452_ ( .A1(_07846_ ), .A2(\ICACHE.tag_reg[0][7] ), .A3(_07850_ ), .ZN(_07853_ ) );
INV_X1 _15453_ ( .A(\ICACHE.s_axi_araddr [12] ), .ZN(_07854_ ) );
OAI21_X1 _15454_ ( .A(_07853_ ), .B1(_07854_ ), .B2(_07848_ ), .ZN(_00572_ ) );
NAND3_X1 _15455_ ( .A1(_07846_ ), .A2(\ICACHE.tag_reg[0][6] ), .A3(_07850_ ), .ZN(_07855_ ) );
OAI21_X1 _15456_ ( .A(_07855_ ), .B1(_07618_ ), .B2(_07848_ ), .ZN(_00573_ ) );
NAND3_X1 _15457_ ( .A1(_07846_ ), .A2(\ICACHE.tag_reg[0][5] ), .A3(_07850_ ), .ZN(_07856_ ) );
OAI21_X1 _15458_ ( .A(_07856_ ), .B1(_07577_ ), .B2(_07848_ ), .ZN(_00574_ ) );
NAND3_X1 _15459_ ( .A1(_07846_ ), .A2(\ICACHE.tag_reg[0][4] ), .A3(_07850_ ), .ZN(_07857_ ) );
OAI21_X1 _15460_ ( .A(_07857_ ), .B1(_07626_ ), .B2(_07848_ ), .ZN(_00575_ ) );
NAND3_X1 _15461_ ( .A1(_07846_ ), .A2(\ICACHE.tag_reg[0][3] ), .A3(_07850_ ), .ZN(_07858_ ) );
OAI21_X1 _15462_ ( .A(_07858_ ), .B1(_07562_ ), .B2(_07848_ ), .ZN(_00576_ ) );
NAND3_X1 _15463_ ( .A1(_07845_ ), .A2(\ICACHE.tag_reg[0][2] ), .A3(_07850_ ), .ZN(_07859_ ) );
INV_X1 _15464_ ( .A(\ICACHE.s_axi_araddr [7] ), .ZN(_07860_ ) );
OAI21_X1 _15465_ ( .A(_07859_ ), .B1(_07860_ ), .B2(_07848_ ), .ZN(_00577_ ) );
NAND3_X1 _15466_ ( .A1(_07845_ ), .A2(\ICACHE.tag_reg[0][1] ), .A3(_07850_ ), .ZN(_07861_ ) );
OAI21_X1 _15467_ ( .A(_07861_ ), .B1(_07555_ ), .B2(_07846_ ), .ZN(_00578_ ) );
NAND2_X1 _15468_ ( .A1(_07692_ ), .A2(_07601_ ), .ZN(_07862_ ) );
BUF_X4 _15469_ ( .A(_07862_ ), .Z(_07863_ ) );
NAND3_X1 _15470_ ( .A1(_07863_ ), .A2(\ICACHE.tag_reg[1][10] ), .A3(_07850_ ), .ZN(_07864_ ) );
BUF_X4 _15471_ ( .A(_07862_ ), .Z(_07865_ ) );
OAI21_X1 _15472_ ( .A(_07864_ ), .B1(_07634_ ), .B2(_07865_ ), .ZN(_00579_ ) );
BUF_X4 _15473_ ( .A(_03808_ ), .Z(_07866_ ) );
NAND3_X1 _15474_ ( .A1(_07863_ ), .A2(\ICACHE.tag_reg[1][9] ), .A3(_07866_ ), .ZN(_07867_ ) );
OAI21_X1 _15475_ ( .A(_07867_ ), .B1(_07584_ ), .B2(_07865_ ), .ZN(_00580_ ) );
NAND3_X1 _15476_ ( .A1(_07863_ ), .A2(\ICACHE.tag_reg[1][0] ), .A3(_07866_ ), .ZN(_07868_ ) );
OAI21_X1 _15477_ ( .A(_07868_ ), .B1(_07605_ ), .B2(_07865_ ), .ZN(_00581_ ) );
NAND3_X1 _15478_ ( .A1(_07863_ ), .A2(\ICACHE.tag_reg[1][8] ), .A3(_07866_ ), .ZN(_07869_ ) );
OAI21_X1 _15479_ ( .A(_07869_ ), .B1(_07593_ ), .B2(_07865_ ), .ZN(_00582_ ) );
NAND3_X1 _15480_ ( .A1(_07863_ ), .A2(\ICACHE.tag_reg[1][7] ), .A3(_07866_ ), .ZN(_07870_ ) );
OAI21_X1 _15481_ ( .A(_07870_ ), .B1(_07854_ ), .B2(_07865_ ), .ZN(_00583_ ) );
NAND3_X1 _15482_ ( .A1(_07863_ ), .A2(\ICACHE.tag_reg[1][6] ), .A3(_07866_ ), .ZN(_07871_ ) );
OAI21_X1 _15483_ ( .A(_07871_ ), .B1(_07618_ ), .B2(_07865_ ), .ZN(_00584_ ) );
NAND3_X1 _15484_ ( .A1(_07863_ ), .A2(\ICACHE.tag_reg[1][5] ), .A3(_07866_ ), .ZN(_07872_ ) );
OAI21_X1 _15485_ ( .A(_07872_ ), .B1(_07577_ ), .B2(_07865_ ), .ZN(_00585_ ) );
NAND3_X1 _15486_ ( .A1(_07863_ ), .A2(\ICACHE.tag_reg[1][4] ), .A3(_07866_ ), .ZN(_07873_ ) );
OAI21_X1 _15487_ ( .A(_07873_ ), .B1(_07626_ ), .B2(_07865_ ), .ZN(_00586_ ) );
NAND3_X1 _15488_ ( .A1(_07863_ ), .A2(\ICACHE.tag_reg[1][3] ), .A3(_07866_ ), .ZN(_07874_ ) );
OAI21_X1 _15489_ ( .A(_07874_ ), .B1(_07562_ ), .B2(_07865_ ), .ZN(_00587_ ) );
NAND3_X1 _15490_ ( .A1(_07862_ ), .A2(\ICACHE.tag_reg[1][2] ), .A3(_07866_ ), .ZN(_07875_ ) );
OAI21_X1 _15491_ ( .A(_07875_ ), .B1(_07860_ ), .B2(_07865_ ), .ZN(_00588_ ) );
NAND3_X1 _15492_ ( .A1(_07862_ ), .A2(\ICACHE.tag_reg[1][1] ), .A3(_07866_ ), .ZN(_07876_ ) );
OAI21_X1 _15493_ ( .A(_07876_ ), .B1(_07555_ ), .B2(_07863_ ), .ZN(_00589_ ) );
INV_X2 _15494_ ( .A(_05509_ ), .ZN(_07877_ ) );
AND4_X1 _15495_ ( .A1(_03732_ ), .A2(_03745_ ), .A3(_03733_ ), .A4(_03722_ ), .ZN(_07878_ ) );
NAND3_X1 _15496_ ( .A1(_07877_ ), .A2(\IDU.state ), .A3(_07878_ ), .ZN(_07879_ ) );
NAND4_X1 _15497_ ( .A1(_07670_ ), .A2(_07675_ ), .A3(_07665_ ), .A4(_07680_ ), .ZN(_07880_ ) );
AOI21_X1 _15498_ ( .A(fanout_net_11 ), .B1(_07880_ ), .B2(_07660_ ), .ZN(_07881_ ) );
NAND2_X2 _15499_ ( .A1(_07879_ ), .A2(_07881_ ), .ZN(_07882_ ) );
NOR2_X1 _15500_ ( .A1(_07882_ ), .A2(_07795_ ), .ZN(_07883_ ) );
AND3_X1 _15501_ ( .A1(_07879_ ), .A2(\ICACHE.valid_reg[0][0] ), .A3(_07881_ ), .ZN(_07884_ ) );
BUF_X4 _15502_ ( .A(_07693_ ), .Z(_07885_ ) );
BUF_X4 _15503_ ( .A(_07885_ ), .Z(_07886_ ) );
OR3_X1 _15504_ ( .A1(_04110_ ), .A2(_04113_ ), .A3(io_master_arready ), .ZN(_07887_ ) );
OAI211_X1 _15505_ ( .A(\CLINT.c_axi_arready_$_NOT__A_Y ), .B(_04091_ ), .C1(_04076_ ), .C2(_04100_ ), .ZN(_07888_ ) );
INV_X1 _15506_ ( .A(\ICACHE.s_axi_arvalid ), .ZN(_07889_ ) );
NOR4_X1 _15507_ ( .A1(_04055_ ), .A2(_07889_ ), .A3(_07535_ ), .A4(\Xbar.state [2] ), .ZN(_07890_ ) );
NAND3_X1 _15508_ ( .A1(_07887_ ), .A2(_07888_ ), .A3(_07890_ ), .ZN(_07891_ ) );
NOR2_X1 _15509_ ( .A1(_07882_ ), .A2(_07891_ ), .ZN(_07892_ ) );
OAI21_X1 _15510_ ( .A(_07886_ ), .B1(_07883_ ), .B2(_07892_ ), .ZN(_07893_ ) );
MUX2_X1 _15511_ ( .A(_07883_ ), .B(_07884_ ), .S(_07893_ ), .Z(_00590_ ) );
NOR2_X1 _15512_ ( .A1(_07882_ ), .A2(_07805_ ), .ZN(_07894_ ) );
AND3_X1 _15513_ ( .A1(_07879_ ), .A2(\ICACHE.valid_reg[0][1] ), .A3(_07881_ ), .ZN(_07895_ ) );
OAI21_X1 _15514_ ( .A(_07886_ ), .B1(_07892_ ), .B2(_07894_ ), .ZN(_07896_ ) );
MUX2_X1 _15515_ ( .A(_07894_ ), .B(_07895_ ), .S(_07896_ ), .Z(_00591_ ) );
NOR2_X1 _15516_ ( .A1(_07882_ ), .A2(_07814_ ), .ZN(_07897_ ) );
AND3_X1 _15517_ ( .A1(_07879_ ), .A2(\ICACHE.valid_reg[0][2] ), .A3(_07881_ ), .ZN(_07898_ ) );
OAI21_X1 _15518_ ( .A(_07886_ ), .B1(_07892_ ), .B2(_07897_ ), .ZN(_07899_ ) );
MUX2_X1 _15519_ ( .A(_07897_ ), .B(_07898_ ), .S(_07899_ ), .Z(_00592_ ) );
NOR2_X1 _15520_ ( .A1(_07882_ ), .A2(_07824_ ), .ZN(_07900_ ) );
AND3_X1 _15521_ ( .A1(_07879_ ), .A2(\ICACHE.valid_reg[0][3] ), .A3(_07881_ ), .ZN(_07901_ ) );
OAI21_X1 _15522_ ( .A(_07886_ ), .B1(_07892_ ), .B2(_07900_ ), .ZN(_07902_ ) );
MUX2_X1 _15523_ ( .A(_07900_ ), .B(_07901_ ), .S(_07902_ ), .Z(_00593_ ) );
AND3_X1 _15524_ ( .A1(_07879_ ), .A2(\ICACHE.valid_reg[1][1] ), .A3(_07881_ ), .ZN(_07903_ ) );
OAI21_X1 _15525_ ( .A(_07601_ ), .B1(_07892_ ), .B2(_07894_ ), .ZN(_07904_ ) );
MUX2_X1 _15526_ ( .A(_07894_ ), .B(_07903_ ), .S(_07904_ ), .Z(_00594_ ) );
AND3_X1 _15527_ ( .A1(_07879_ ), .A2(\ICACHE.valid_reg[1][2] ), .A3(_07881_ ), .ZN(_07905_ ) );
OAI21_X1 _15528_ ( .A(_07601_ ), .B1(_07892_ ), .B2(_07897_ ), .ZN(_07906_ ) );
MUX2_X1 _15529_ ( .A(_07897_ ), .B(_07905_ ), .S(_07906_ ), .Z(_00595_ ) );
AND3_X1 _15530_ ( .A1(_07879_ ), .A2(\ICACHE.valid_reg[1][0] ), .A3(_07881_ ), .ZN(_07907_ ) );
OAI21_X1 _15531_ ( .A(_07601_ ), .B1(_07883_ ), .B2(_07892_ ), .ZN(_07908_ ) );
MUX2_X1 _15532_ ( .A(_07883_ ), .B(_07907_ ), .S(_07908_ ), .Z(_00596_ ) );
AND3_X1 _15533_ ( .A1(_07879_ ), .A2(\ICACHE.valid_reg[1][3] ), .A3(_07881_ ), .ZN(_07909_ ) );
OAI21_X1 _15534_ ( .A(_07601_ ), .B1(_07892_ ), .B2(_07900_ ), .ZN(_07910_ ) );
MUX2_X1 _15535_ ( .A(_07900_ ), .B(_07909_ ), .S(_07910_ ), .Z(_00597_ ) );
MUX2_X1 _15536_ ( .A(\EXU.funct3_i [2] ), .B(\IDU.funct3 [2] ), .S(\IDU.updata ), .Z(_00598_ ) );
MUX2_X1 _15537_ ( .A(\EXU.funct3_i [1] ), .B(\IDU.funct3 [1] ), .S(\IDU.updata ), .Z(_00599_ ) );
MUX2_X1 _15538_ ( .A(\EXU.funct3_i [0] ), .B(\IDU.funct3 [0] ), .S(\IDU.updata ), .Z(_00600_ ) );
BUF_X4 _15539_ ( .A(_05513_ ), .Z(_07911_ ) );
BUF_X4 _15540_ ( .A(_07911_ ), .Z(_07912_ ) );
MUX2_X1 _15541_ ( .A(\EXU.imm_i [31] ), .B(_05479_ ), .S(_07912_ ), .Z(_00601_ ) );
MUX2_X1 _15542_ ( .A(\EXU.imm_i [30] ), .B(_05474_ ), .S(_07912_ ), .Z(_00602_ ) );
MUX2_X1 _15543_ ( .A(\EXU.imm_i [21] ), .B(_05460_ ), .S(_07912_ ), .Z(_00603_ ) );
MUX2_X1 _15544_ ( .A(\EXU.imm_i [20] ), .B(_05462_ ), .S(_07912_ ), .Z(_00604_ ) );
OAI21_X1 _15545_ ( .A(\IDU.immJ [19] ), .B1(_03755_ ), .B2(_03928_ ), .ZN(_07913_ ) );
OAI21_X1 _15546_ ( .A(_07913_ ), .B1(_03741_ ), .B2(_03926_ ), .ZN(_07914_ ) );
MUX2_X1 _15547_ ( .A(\EXU.imm_i [19] ), .B(_07914_ ), .S(_07912_ ), .Z(_00605_ ) );
OAI21_X1 _15548_ ( .A(_03934_ ), .B1(_05497_ ), .B2(_03929_ ), .ZN(_07915_ ) );
MUX2_X1 _15549_ ( .A(\EXU.imm_i [18] ), .B(_07915_ ), .S(_07912_ ), .Z(_00606_ ) );
OAI21_X1 _15550_ ( .A(_03934_ ), .B1(_05502_ ), .B2(_03929_ ), .ZN(_07916_ ) );
MUX2_X1 _15551_ ( .A(\EXU.imm_i [17] ), .B(_07916_ ), .S(_07912_ ), .Z(_00607_ ) );
OAI21_X1 _15552_ ( .A(_03934_ ), .B1(_05505_ ), .B2(_03929_ ), .ZN(_07917_ ) );
MUX2_X1 _15553_ ( .A(\EXU.imm_i [16] ), .B(_07917_ ), .S(_07912_ ), .Z(_00608_ ) );
MUX2_X1 _15554_ ( .A(\EXU.imm_i [15] ), .B(_03951_ ), .S(_07912_ ), .Z(_00609_ ) );
MUX2_X1 _15555_ ( .A(\EXU.imm_i [14] ), .B(_03946_ ), .S(_07912_ ), .Z(_00610_ ) );
AND2_X1 _15556_ ( .A1(_03934_ ), .A2(_03935_ ), .ZN(_07918_ ) );
INV_X1 _15557_ ( .A(_07918_ ), .ZN(_07919_ ) );
BUF_X4 _15558_ ( .A(_07911_ ), .Z(_07920_ ) );
MUX2_X1 _15559_ ( .A(\EXU.imm_i [13] ), .B(_07919_ ), .S(_07920_ ), .Z(_00611_ ) );
INV_X1 _15560_ ( .A(_03932_ ), .ZN(_07921_ ) );
MUX2_X1 _15561_ ( .A(\EXU.imm_i [12] ), .B(_07921_ ), .S(_07920_ ), .Z(_00612_ ) );
MUX2_X1 _15562_ ( .A(\EXU.imm_i [29] ), .B(_05472_ ), .S(_07920_ ), .Z(_00613_ ) );
AND2_X1 _15563_ ( .A1(_03900_ ), .A2(_03901_ ), .ZN(_07922_ ) );
OR4_X1 _15564_ ( .A1(\EXU.state ), .A2(_05509_ ), .A3(_05510_ ), .A4(_07922_ ), .ZN(_07923_ ) );
OAI21_X1 _15565_ ( .A(_07923_ ), .B1(\IDU.updata ), .B2(_04344_ ), .ZN(_00614_ ) );
MUX2_X1 _15566_ ( .A(\EXU.funct7_i ), .B(_03919_ ), .S(_07920_ ), .Z(_00615_ ) );
MUX2_X1 _15567_ ( .A(\EXU.imm_i [9] ), .B(_03915_ ), .S(_07920_ ), .Z(_00616_ ) );
MUX2_X1 _15568_ ( .A(\EXU.imm_i [8] ), .B(_03906_ ), .S(_07920_ ), .Z(_00617_ ) );
MUX2_X1 _15569_ ( .A(\EXU.imm_i [7] ), .B(_03792_ ), .S(_07920_ ), .Z(_00618_ ) );
MUX2_X1 _15570_ ( .A(\EXU.imm_i [6] ), .B(_03788_ ), .S(_07920_ ), .Z(_00619_ ) );
MUX2_X1 _15571_ ( .A(\EXU.imm_i [5] ), .B(_03785_ ), .S(_07920_ ), .Z(_00620_ ) );
MUX2_X1 _15572_ ( .A(\EXU.imm_i [4] ), .B(_05441_ ), .S(_07920_ ), .Z(_00621_ ) );
BUF_X4 _15573_ ( .A(_07911_ ), .Z(_07924_ ) );
MUX2_X1 _15574_ ( .A(\EXU.imm_i [3] ), .B(_03777_ ), .S(_07924_ ), .Z(_00622_ ) );
MUX2_X1 _15575_ ( .A(\EXU.imm_i [2] ), .B(_03772_ ), .S(_07924_ ), .Z(_00623_ ) );
MUX2_X1 _15576_ ( .A(\EXU.imm_i [28] ), .B(_05470_ ), .S(_07924_ ), .Z(_00624_ ) );
MUX2_X1 _15577_ ( .A(\EXU.imm_i [1] ), .B(_03770_ ), .S(_07924_ ), .Z(_00625_ ) );
MUX2_X1 _15578_ ( .A(\EXU.imm_i [0] ), .B(_03835_ ), .S(_07924_ ), .Z(_00626_ ) );
MUX2_X1 _15579_ ( .A(\EXU.imm_i [27] ), .B(_05476_ ), .S(_07924_ ), .Z(_00627_ ) );
MUX2_X1 _15580_ ( .A(\EXU.imm_i [26] ), .B(_05453_ ), .S(_07924_ ), .Z(_00628_ ) );
MUX2_X1 _15581_ ( .A(\EXU.imm_i [25] ), .B(_05451_ ), .S(_07924_ ), .Z(_00629_ ) );
MUX2_X1 _15582_ ( .A(\EXU.imm_i [24] ), .B(_05455_ ), .S(_07924_ ), .Z(_00630_ ) );
MUX2_X1 _15583_ ( .A(\EXU.imm_i [23] ), .B(_05457_ ), .S(_07924_ ), .Z(_00631_ ) );
BUF_X4 _15584_ ( .A(_07911_ ), .Z(_07925_ ) );
MUX2_X1 _15585_ ( .A(\EXU.imm_i [22] ), .B(_05466_ ), .S(_07925_ ), .Z(_00632_ ) );
AND3_X1 _15586_ ( .A1(_03721_ ), .A2(_03733_ ), .A3(_03722_ ), .ZN(_07926_ ) );
AND2_X1 _15587_ ( .A1(_07926_ ), .A2(\IDU.ls_valid_o_$_DFFE_PP__Q_D_$_ANDNOT__Y_B_$_NOR__Y_B_$_ANDNOT__Y_A ), .ZN(_07927_ ) );
OAI221_X1 _15588_ ( .A(\IDU.state ), .B1(_03725_ ), .B2(_07927_ ), .C1(\IDU.updata ), .C2(\IDU.ls_valid_o_$_DFFE_PP__Q_E_$_OR__Y_B ), .ZN(_07928_ ) );
INV_X1 _15589_ ( .A(\IDU.ls_valid_o ), .ZN(_07929_ ) );
OR3_X1 _15590_ ( .A1(_07911_ ), .A2(_07929_ ), .A3(\IDU.ls_valid_o_$_DFFE_PP__Q_E_$_OR__Y_B ), .ZN(_07930_ ) );
NAND2_X1 _15591_ ( .A1(_07928_ ), .A2(_07930_ ), .ZN(_00633_ ) );
MUX2_X1 _15592_ ( .A(\EXU.op_i [4] ), .B(\IDU.inst_i [6] ), .S(_07925_ ), .Z(_00634_ ) );
MUX2_X1 _15593_ ( .A(\EXU.op_i [3] ), .B(\IDU.inst_i [5] ), .S(_07925_ ), .Z(_00635_ ) );
MUX2_X1 _15594_ ( .A(\EXU.op_i [2] ), .B(\IDU.inst_i [4] ), .S(_07925_ ), .Z(_00636_ ) );
MUX2_X1 _15595_ ( .A(\EXU.op_i [1] ), .B(\IDU.inst_i [3] ), .S(_07925_ ), .Z(_00637_ ) );
MUX2_X1 _15596_ ( .A(\EXU.op_i [0] ), .B(\IDU.inst_i [2] ), .S(_07925_ ), .Z(_00638_ ) );
MUX2_X1 _15597_ ( .A(\EXU.pc_i [31] ), .B(\BTB.prepc_tag_i [31] ), .S(_07925_ ), .Z(_00639_ ) );
MUX2_X1 _15598_ ( .A(\EXU.pc_i [30] ), .B(\BTB.prepc_tag_i [30] ), .S(_07925_ ), .Z(_00640_ ) );
MUX2_X1 _15599_ ( .A(\EXU.pc_i [21] ), .B(\BTB.prepc_tag_i [21] ), .S(_07925_ ), .Z(_00641_ ) );
MUX2_X1 _15600_ ( .A(\EXU.pc_i [20] ), .B(\BTB.prepc_tag_i [20] ), .S(_07925_ ), .Z(_00642_ ) );
BUF_X4 _15601_ ( .A(_05514_ ), .Z(_07931_ ) );
MUX2_X1 _15602_ ( .A(\EXU.pc_i [19] ), .B(\BTB.prepc_tag_i [19] ), .S(_07931_ ), .Z(_00643_ ) );
MUX2_X1 _15603_ ( .A(\EXU.pc_i [18] ), .B(\BTB.prepc_tag_i [18] ), .S(_07931_ ), .Z(_00644_ ) );
MUX2_X1 _15604_ ( .A(\EXU.pc_i [17] ), .B(\BTB.prepc_tag_i [17] ), .S(_07931_ ), .Z(_00645_ ) );
MUX2_X1 _15605_ ( .A(\EXU.pc_i [16] ), .B(\BTB.prepc_tag_i [16] ), .S(_07931_ ), .Z(_00646_ ) );
MUX2_X1 _15606_ ( .A(\EXU.pc_i [15] ), .B(\BTB.btag_pre [12] ), .S(_07931_ ), .Z(_00647_ ) );
MUX2_X1 _15607_ ( .A(\EXU.pc_i [14] ), .B(\BTB.btag_pre [11] ), .S(_07931_ ), .Z(_00648_ ) );
MUX2_X1 _15608_ ( .A(\EXU.pc_i [13] ), .B(\BTB.btag_pre [10] ), .S(_07931_ ), .Z(_00649_ ) );
MUX2_X1 _15609_ ( .A(\EXU.pc_i [12] ), .B(\BTB.btag_pre [9] ), .S(_07931_ ), .Z(_00650_ ) );
MUX2_X1 _15610_ ( .A(\EXU.pc_i [29] ), .B(\BTB.prepc_tag_i [29] ), .S(_07931_ ), .Z(_00651_ ) );
MUX2_X1 _15611_ ( .A(\EXU.pc_i [11] ), .B(\BTB.btag_pre [8] ), .S(_07931_ ), .Z(_00652_ ) );
BUF_X4 _15612_ ( .A(_05514_ ), .Z(_07932_ ) );
MUX2_X1 _15613_ ( .A(\EXU.pc_i [10] ), .B(\BTB.btag_pre [7] ), .S(_07932_ ), .Z(_00653_ ) );
MUX2_X1 _15614_ ( .A(\EXU.pc_i [9] ), .B(\BTB.btag_pre [6] ), .S(_07932_ ), .Z(_00654_ ) );
MUX2_X1 _15615_ ( .A(\EXU.pc_i [8] ), .B(\BTB.btag_pre [5] ), .S(_07932_ ), .Z(_00655_ ) );
MUX2_X1 _15616_ ( .A(\EXU.pc_i [7] ), .B(\BTB.btag_pre [4] ), .S(_07932_ ), .Z(_00656_ ) );
MUX2_X1 _15617_ ( .A(\EXU.pc_i [6] ), .B(\BTB.btag_pre [3] ), .S(_07932_ ), .Z(_00657_ ) );
MUX2_X1 _15618_ ( .A(\EXU.pc_i [5] ), .B(\BTB.btag_pre [2] ), .S(_07932_ ), .Z(_00658_ ) );
MUX2_X1 _15619_ ( .A(\EXU.pc_i [4] ), .B(\BTB.btag_pre [1] ), .S(_07932_ ), .Z(_00659_ ) );
MUX2_X1 _15620_ ( .A(\EXU.pc_i [3] ), .B(\BTB.btag_pre [0] ), .S(_07932_ ), .Z(_00660_ ) );
MUX2_X1 _15621_ ( .A(\EXU.pc_i [2] ), .B(\BTB.bindex_pre ), .S(_07932_ ), .Z(_00661_ ) );
MUX2_X1 _15622_ ( .A(\EXU.pc_i [28] ), .B(\BTB.prepc_tag_i [28] ), .S(_07932_ ), .Z(_00662_ ) );
BUF_X4 _15623_ ( .A(_05514_ ), .Z(_07933_ ) );
MUX2_X1 _15624_ ( .A(\EXU.add_pc_4 [1] ), .B(\BTB.prepc_tag_i [1] ), .S(_07933_ ), .Z(_00663_ ) );
MUX2_X1 _15625_ ( .A(\EXU.add_pc_4 [0] ), .B(\BTB.prepc_tag_i [0] ), .S(_07933_ ), .Z(_00664_ ) );
MUX2_X1 _15626_ ( .A(\EXU.pc_i [27] ), .B(\BTB.prepc_tag_i [27] ), .S(_07933_ ), .Z(_00665_ ) );
MUX2_X1 _15627_ ( .A(\EXU.pc_i [26] ), .B(\BTB.prepc_tag_i [26] ), .S(_07933_ ), .Z(_00666_ ) );
MUX2_X1 _15628_ ( .A(\EXU.pc_i [25] ), .B(\BTB.prepc_tag_i [25] ), .S(_07933_ ), .Z(_00667_ ) );
MUX2_X1 _15629_ ( .A(\EXU.pc_i [24] ), .B(\BTB.prepc_tag_i [24] ), .S(_07933_ ), .Z(_00668_ ) );
MUX2_X1 _15630_ ( .A(\EXU.pc_i [23] ), .B(\BTB.prepc_tag_i [23] ), .S(_07933_ ), .Z(_00669_ ) );
MUX2_X1 _15631_ ( .A(\EXU.pc_i [22] ), .B(\BTB.prepc_tag_i [22] ), .S(_07933_ ), .Z(_00670_ ) );
INV_X1 _15632_ ( .A(_05500_ ), .ZN(_07934_ ) );
AND2_X1 _15633_ ( .A1(_07934_ ), .A2(_05506_ ), .ZN(_07935_ ) );
BUF_X4 _15634_ ( .A(_07935_ ), .Z(_07936_ ) );
BUF_X4 _15635_ ( .A(_07936_ ), .Z(_07937_ ) );
AND2_X1 _15636_ ( .A1(_05498_ ), .A2(_05503_ ), .ZN(_07938_ ) );
BUF_X4 _15637_ ( .A(_07938_ ), .Z(_07939_ ) );
BUF_X4 _15638_ ( .A(_07939_ ), .Z(_07940_ ) );
NAND3_X1 _15639_ ( .A1(_07937_ ), .A2(\RFU.rf[14][31] ), .A3(_07940_ ), .ZN(_07941_ ) );
INV_X1 _15640_ ( .A(_05498_ ), .ZN(_07942_ ) );
AND2_X1 _15641_ ( .A1(_07942_ ), .A2(_05503_ ), .ZN(_07943_ ) );
BUF_X4 _15642_ ( .A(_07943_ ), .Z(_07944_ ) );
BUF_X4 _15643_ ( .A(_07944_ ), .Z(_07945_ ) );
NOR2_X2 _15644_ ( .A1(_05500_ ), .A2(_05506_ ), .ZN(_07946_ ) );
BUF_X4 _15645_ ( .A(_07946_ ), .Z(_07947_ ) );
NAND3_X1 _15646_ ( .A1(_07945_ ), .A2(\RFU.rf[4][31] ), .A3(_07947_ ), .ZN(_07948_ ) );
BUF_X4 _15647_ ( .A(_07944_ ), .Z(_07949_ ) );
AND2_X1 _15648_ ( .A1(_05500_ ), .A2(_05506_ ), .ZN(_07950_ ) );
BUF_X4 _15649_ ( .A(_07950_ ), .Z(_07951_ ) );
BUF_X4 _15650_ ( .A(_07951_ ), .Z(_07952_ ) );
NAND3_X1 _15651_ ( .A1(_07949_ ), .A2(\RFU.rf[7][31] ), .A3(_07952_ ), .ZN(_07953_ ) );
BUF_X4 _15652_ ( .A(_07939_ ), .Z(_07954_ ) );
BUF_X4 _15653_ ( .A(_07950_ ), .Z(_07955_ ) );
BUF_X4 _15654_ ( .A(_07955_ ), .Z(_07956_ ) );
NAND3_X1 _15655_ ( .A1(_07954_ ), .A2(_07956_ ), .A3(\RFU.rf[15][31] ), .ZN(_07957_ ) );
NAND4_X1 _15656_ ( .A1(_07941_ ), .A2(_07948_ ), .A3(_07953_ ), .A4(_07957_ ), .ZN(_07958_ ) );
BUF_X2 _15657_ ( .A(_07936_ ), .Z(_07959_ ) );
NOR2_X1 _15658_ ( .A1(_05498_ ), .A2(_05503_ ), .ZN(_07960_ ) );
CLKBUF_X2 _15659_ ( .A(_07960_ ), .Z(_07961_ ) );
AND3_X1 _15660_ ( .A1(_07959_ ), .A2(\RFU.rf[2][31] ), .A3(_07961_ ), .ZN(_07962_ ) );
BUF_X2 _15661_ ( .A(_07944_ ), .Z(_07963_ ) );
CLKBUF_X2 _15662_ ( .A(_07936_ ), .Z(_07964_ ) );
AND3_X1 _15663_ ( .A1(_07963_ ), .A2(_07964_ ), .A3(\RFU.rf[6][31] ), .ZN(_07965_ ) );
BUF_X2 _15664_ ( .A(_07955_ ), .Z(_07966_ ) );
CLKBUF_X2 _15665_ ( .A(_07960_ ), .Z(_07967_ ) );
AND3_X1 _15666_ ( .A1(_07966_ ), .A2(\RFU.rf[3][31] ), .A3(_07967_ ), .ZN(_07968_ ) );
NOR4_X1 _15667_ ( .A1(_07958_ ), .A2(_07962_ ), .A3(_07965_ ), .A4(_07968_ ), .ZN(_07969_ ) );
BUF_X4 _15668_ ( .A(_07943_ ), .Z(_07970_ ) );
BUF_X4 _15669_ ( .A(_07970_ ), .Z(_07971_ ) );
NOR2_X1 _15670_ ( .A1(_07934_ ), .A2(_05506_ ), .ZN(_07972_ ) );
BUF_X8 _15671_ ( .A(_07972_ ), .Z(_07973_ ) );
BUF_X4 _15672_ ( .A(_07973_ ), .Z(_07974_ ) );
NAND3_X1 _15673_ ( .A1(_07971_ ), .A2(_07974_ ), .A3(\RFU.rf[5][31] ), .ZN(_07975_ ) );
BUF_X4 _15674_ ( .A(_07973_ ), .Z(_07976_ ) );
NOR2_X1 _15675_ ( .A1(_07942_ ), .A2(_05503_ ), .ZN(_07977_ ) );
BUF_X4 _15676_ ( .A(_07977_ ), .Z(_07978_ ) );
BUF_X4 _15677_ ( .A(_07978_ ), .Z(_07979_ ) );
NAND3_X1 _15678_ ( .A1(_07976_ ), .A2(_07979_ ), .A3(\RFU.rf[9][31] ), .ZN(_07980_ ) );
BUF_X4 _15679_ ( .A(_07973_ ), .Z(_07981_ ) );
BUF_X4 _15680_ ( .A(_07960_ ), .Z(_07982_ ) );
BUF_X4 _15681_ ( .A(_07982_ ), .Z(_07983_ ) );
NAND3_X1 _15682_ ( .A1(_07981_ ), .A2(\RFU.rf[1][31] ), .A3(_07983_ ), .ZN(_07984_ ) );
BUF_X4 _15683_ ( .A(_07938_ ), .Z(_07985_ ) );
BUF_X4 _15684_ ( .A(_07985_ ), .Z(_07986_ ) );
BUF_X4 _15685_ ( .A(_07946_ ), .Z(_07987_ ) );
BUF_X4 _15686_ ( .A(_07987_ ), .Z(_07988_ ) );
NAND3_X1 _15687_ ( .A1(_07986_ ), .A2(_07988_ ), .A3(\RFU.rf[12][31] ), .ZN(_07989_ ) );
AND4_X1 _15688_ ( .A1(_07975_ ), .A2(_07980_ ), .A3(_07984_ ), .A4(_07989_ ), .ZN(_07990_ ) );
BUF_X4 _15689_ ( .A(_07972_ ), .Z(_07991_ ) );
BUF_X4 _15690_ ( .A(_07991_ ), .Z(_07992_ ) );
BUF_X4 _15691_ ( .A(_07985_ ), .Z(_07993_ ) );
NAND3_X1 _15692_ ( .A1(_07992_ ), .A2(\RFU.rf[13][31] ), .A3(_07993_ ), .ZN(_07994_ ) );
BUF_X4 _15693_ ( .A(_07935_ ), .Z(_07995_ ) );
BUF_X4 _15694_ ( .A(_07995_ ), .Z(_07996_ ) );
BUF_X8 _15695_ ( .A(_07977_ ), .Z(_07997_ ) );
BUF_X4 _15696_ ( .A(_07997_ ), .Z(_07998_ ) );
NAND3_X1 _15697_ ( .A1(_07996_ ), .A2(\RFU.rf[10][31] ), .A3(_07998_ ), .ZN(_07999_ ) );
BUF_X4 _15698_ ( .A(_07997_ ), .Z(_08000_ ) );
BUF_X4 _15699_ ( .A(_07946_ ), .Z(_08001_ ) );
NAND3_X1 _15700_ ( .A1(_08000_ ), .A2(\RFU.rf[8][31] ), .A3(_08001_ ), .ZN(_08002_ ) );
BUF_X4 _15701_ ( .A(_07997_ ), .Z(_08003_ ) );
BUF_X4 _15702_ ( .A(_07951_ ), .Z(_08004_ ) );
NAND3_X1 _15703_ ( .A1(_08003_ ), .A2(\RFU.rf[11][31] ), .A3(_08004_ ), .ZN(_08005_ ) );
AND4_X1 _15704_ ( .A1(_07994_ ), .A2(_07999_ ), .A3(_08002_ ), .A4(_08005_ ), .ZN(_08006_ ) );
NAND3_X1 _15705_ ( .A1(_07969_ ), .A2(_07990_ ), .A3(_08006_ ), .ZN(_08007_ ) );
MUX2_X1 _15706_ ( .A(\EXU.r1_i [31] ), .B(_08007_ ), .S(_07933_ ), .Z(_00671_ ) );
NAND3_X1 _15707_ ( .A1(_07937_ ), .A2(\RFU.rf[14][30] ), .A3(_07940_ ), .ZN(_08008_ ) );
NAND3_X1 _15708_ ( .A1(_07945_ ), .A2(\RFU.rf[4][30] ), .A3(_07947_ ), .ZN(_08009_ ) );
NAND3_X1 _15709_ ( .A1(_07949_ ), .A2(\RFU.rf[7][30] ), .A3(_07952_ ), .ZN(_08010_ ) );
NAND3_X1 _15710_ ( .A1(_07954_ ), .A2(_07956_ ), .A3(\RFU.rf[15][30] ), .ZN(_08011_ ) );
NAND4_X1 _15711_ ( .A1(_08008_ ), .A2(_08009_ ), .A3(_08010_ ), .A4(_08011_ ), .ZN(_08012_ ) );
AND3_X1 _15712_ ( .A1(_07959_ ), .A2(\RFU.rf[2][30] ), .A3(_07961_ ), .ZN(_08013_ ) );
AND3_X1 _15713_ ( .A1(_07963_ ), .A2(_07964_ ), .A3(\RFU.rf[6][30] ), .ZN(_08014_ ) );
AND3_X1 _15714_ ( .A1(_07966_ ), .A2(\RFU.rf[3][30] ), .A3(_07967_ ), .ZN(_08015_ ) );
NOR4_X1 _15715_ ( .A1(_08012_ ), .A2(_08013_ ), .A3(_08014_ ), .A4(_08015_ ), .ZN(_08016_ ) );
NAND3_X1 _15716_ ( .A1(_07971_ ), .A2(_07974_ ), .A3(\RFU.rf[5][30] ), .ZN(_08017_ ) );
NAND3_X1 _15717_ ( .A1(_07976_ ), .A2(_07979_ ), .A3(\RFU.rf[9][30] ), .ZN(_08018_ ) );
NAND3_X1 _15718_ ( .A1(_07981_ ), .A2(\RFU.rf[1][30] ), .A3(_07983_ ), .ZN(_08019_ ) );
NAND3_X1 _15719_ ( .A1(_07986_ ), .A2(_07988_ ), .A3(\RFU.rf[12][30] ), .ZN(_08020_ ) );
AND4_X1 _15720_ ( .A1(_08017_ ), .A2(_08018_ ), .A3(_08019_ ), .A4(_08020_ ), .ZN(_08021_ ) );
NAND3_X1 _15721_ ( .A1(_07992_ ), .A2(\RFU.rf[13][30] ), .A3(_07993_ ), .ZN(_08022_ ) );
NAND3_X1 _15722_ ( .A1(_07996_ ), .A2(\RFU.rf[10][30] ), .A3(_07998_ ), .ZN(_08023_ ) );
NAND3_X1 _15723_ ( .A1(_08000_ ), .A2(\RFU.rf[8][30] ), .A3(_08001_ ), .ZN(_08024_ ) );
NAND3_X1 _15724_ ( .A1(_08003_ ), .A2(\RFU.rf[11][30] ), .A3(_08004_ ), .ZN(_08025_ ) );
AND4_X1 _15725_ ( .A1(_08022_ ), .A2(_08023_ ), .A3(_08024_ ), .A4(_08025_ ), .ZN(_08026_ ) );
NAND3_X1 _15726_ ( .A1(_08016_ ), .A2(_08021_ ), .A3(_08026_ ), .ZN(_08027_ ) );
MUX2_X1 _15727_ ( .A(\EXU.r1_i [30] ), .B(_08027_ ), .S(_07933_ ), .Z(_00672_ ) );
NAND3_X1 _15728_ ( .A1(_07937_ ), .A2(\RFU.rf[14][21] ), .A3(_07940_ ), .ZN(_08028_ ) );
NAND3_X1 _15729_ ( .A1(_07945_ ), .A2(\RFU.rf[4][21] ), .A3(_07947_ ), .ZN(_08029_ ) );
NAND3_X1 _15730_ ( .A1(_07949_ ), .A2(\RFU.rf[7][21] ), .A3(_07952_ ), .ZN(_08030_ ) );
NAND3_X1 _15731_ ( .A1(_07954_ ), .A2(_07956_ ), .A3(\RFU.rf[15][21] ), .ZN(_08031_ ) );
NAND4_X1 _15732_ ( .A1(_08028_ ), .A2(_08029_ ), .A3(_08030_ ), .A4(_08031_ ), .ZN(_08032_ ) );
AND3_X1 _15733_ ( .A1(_07959_ ), .A2(\RFU.rf[2][21] ), .A3(_07961_ ), .ZN(_08033_ ) );
AND3_X1 _15734_ ( .A1(_07963_ ), .A2(_07964_ ), .A3(\RFU.rf[6][21] ), .ZN(_08034_ ) );
AND3_X1 _15735_ ( .A1(_07966_ ), .A2(\RFU.rf[3][21] ), .A3(_07967_ ), .ZN(_08035_ ) );
NOR4_X1 _15736_ ( .A1(_08032_ ), .A2(_08033_ ), .A3(_08034_ ), .A4(_08035_ ), .ZN(_08036_ ) );
NAND3_X1 _15737_ ( .A1(_07971_ ), .A2(_07974_ ), .A3(\RFU.rf[5][21] ), .ZN(_08037_ ) );
NAND3_X1 _15738_ ( .A1(_07976_ ), .A2(_07979_ ), .A3(\RFU.rf[9][21] ), .ZN(_08038_ ) );
NAND3_X1 _15739_ ( .A1(_07981_ ), .A2(\RFU.rf[1][21] ), .A3(_07983_ ), .ZN(_08039_ ) );
NAND3_X1 _15740_ ( .A1(_07986_ ), .A2(_07988_ ), .A3(\RFU.rf[12][21] ), .ZN(_08040_ ) );
AND4_X1 _15741_ ( .A1(_08037_ ), .A2(_08038_ ), .A3(_08039_ ), .A4(_08040_ ), .ZN(_08041_ ) );
NAND3_X1 _15742_ ( .A1(_07992_ ), .A2(\RFU.rf[13][21] ), .A3(_07993_ ), .ZN(_08042_ ) );
NAND3_X1 _15743_ ( .A1(_07996_ ), .A2(\RFU.rf[10][21] ), .A3(_07998_ ), .ZN(_08043_ ) );
NAND3_X1 _15744_ ( .A1(_08000_ ), .A2(\RFU.rf[8][21] ), .A3(_08001_ ), .ZN(_08044_ ) );
NAND3_X1 _15745_ ( .A1(_08003_ ), .A2(\RFU.rf[11][21] ), .A3(_08004_ ), .ZN(_08045_ ) );
AND4_X1 _15746_ ( .A1(_08042_ ), .A2(_08043_ ), .A3(_08044_ ), .A4(_08045_ ), .ZN(_08046_ ) );
NAND3_X1 _15747_ ( .A1(_08036_ ), .A2(_08041_ ), .A3(_08046_ ), .ZN(_08047_ ) );
BUF_X4 _15748_ ( .A(_05514_ ), .Z(_08048_ ) );
MUX2_X1 _15749_ ( .A(\EXU.r1_i [21] ), .B(_08047_ ), .S(_08048_ ), .Z(_00673_ ) );
NAND3_X1 _15750_ ( .A1(_07937_ ), .A2(\RFU.rf[14][20] ), .A3(_07940_ ), .ZN(_08049_ ) );
NAND3_X1 _15751_ ( .A1(_07945_ ), .A2(\RFU.rf[4][20] ), .A3(_07947_ ), .ZN(_08050_ ) );
NAND3_X1 _15752_ ( .A1(_07949_ ), .A2(\RFU.rf[7][20] ), .A3(_07952_ ), .ZN(_08051_ ) );
NAND3_X1 _15753_ ( .A1(_07954_ ), .A2(_07956_ ), .A3(\RFU.rf[15][20] ), .ZN(_08052_ ) );
NAND4_X1 _15754_ ( .A1(_08049_ ), .A2(_08050_ ), .A3(_08051_ ), .A4(_08052_ ), .ZN(_08053_ ) );
AND3_X1 _15755_ ( .A1(_07959_ ), .A2(\RFU.rf[2][20] ), .A3(_07961_ ), .ZN(_08054_ ) );
AND3_X1 _15756_ ( .A1(_07963_ ), .A2(_07964_ ), .A3(\RFU.rf[6][20] ), .ZN(_08055_ ) );
AND3_X1 _15757_ ( .A1(_07966_ ), .A2(\RFU.rf[3][20] ), .A3(_07967_ ), .ZN(_08056_ ) );
NOR4_X1 _15758_ ( .A1(_08053_ ), .A2(_08054_ ), .A3(_08055_ ), .A4(_08056_ ), .ZN(_08057_ ) );
NAND3_X1 _15759_ ( .A1(_07971_ ), .A2(_07974_ ), .A3(\RFU.rf[5][20] ), .ZN(_08058_ ) );
NAND3_X1 _15760_ ( .A1(_07976_ ), .A2(_07979_ ), .A3(\RFU.rf[9][20] ), .ZN(_08059_ ) );
NAND3_X1 _15761_ ( .A1(_07981_ ), .A2(\RFU.rf[1][20] ), .A3(_07983_ ), .ZN(_08060_ ) );
NAND3_X1 _15762_ ( .A1(_07986_ ), .A2(_07988_ ), .A3(\RFU.rf[12][20] ), .ZN(_08061_ ) );
AND4_X1 _15763_ ( .A1(_08058_ ), .A2(_08059_ ), .A3(_08060_ ), .A4(_08061_ ), .ZN(_08062_ ) );
NAND3_X1 _15764_ ( .A1(_07992_ ), .A2(\RFU.rf[13][20] ), .A3(_07993_ ), .ZN(_08063_ ) );
NAND3_X1 _15765_ ( .A1(_07996_ ), .A2(\RFU.rf[10][20] ), .A3(_07998_ ), .ZN(_08064_ ) );
NAND3_X1 _15766_ ( .A1(_08000_ ), .A2(\RFU.rf[8][20] ), .A3(_08001_ ), .ZN(_08065_ ) );
NAND3_X1 _15767_ ( .A1(_08003_ ), .A2(\RFU.rf[11][20] ), .A3(_08004_ ), .ZN(_08066_ ) );
AND4_X1 _15768_ ( .A1(_08063_ ), .A2(_08064_ ), .A3(_08065_ ), .A4(_08066_ ), .ZN(_08067_ ) );
NAND3_X1 _15769_ ( .A1(_08057_ ), .A2(_08062_ ), .A3(_08067_ ), .ZN(_08068_ ) );
MUX2_X1 _15770_ ( .A(\EXU.r1_i [20] ), .B(_08068_ ), .S(_08048_ ), .Z(_00674_ ) );
NAND3_X1 _15771_ ( .A1(_07937_ ), .A2(\RFU.rf[14][19] ), .A3(_07940_ ), .ZN(_08069_ ) );
NAND3_X1 _15772_ ( .A1(_07945_ ), .A2(\RFU.rf[4][19] ), .A3(_07947_ ), .ZN(_08070_ ) );
NAND3_X1 _15773_ ( .A1(_07949_ ), .A2(\RFU.rf[7][19] ), .A3(_07952_ ), .ZN(_08071_ ) );
NAND3_X1 _15774_ ( .A1(_07954_ ), .A2(_07956_ ), .A3(\RFU.rf[15][19] ), .ZN(_08072_ ) );
NAND4_X1 _15775_ ( .A1(_08069_ ), .A2(_08070_ ), .A3(_08071_ ), .A4(_08072_ ), .ZN(_08073_ ) );
AND3_X1 _15776_ ( .A1(_07959_ ), .A2(\RFU.rf[2][19] ), .A3(_07961_ ), .ZN(_08074_ ) );
CLKBUF_X2 _15777_ ( .A(_07936_ ), .Z(_08075_ ) );
AND3_X1 _15778_ ( .A1(_07963_ ), .A2(_08075_ ), .A3(\RFU.rf[6][19] ), .ZN(_08076_ ) );
AND3_X1 _15779_ ( .A1(_07966_ ), .A2(\RFU.rf[3][19] ), .A3(_07967_ ), .ZN(_08077_ ) );
NOR4_X1 _15780_ ( .A1(_08073_ ), .A2(_08074_ ), .A3(_08076_ ), .A4(_08077_ ), .ZN(_08078_ ) );
NAND3_X1 _15781_ ( .A1(_07971_ ), .A2(_07974_ ), .A3(\RFU.rf[5][19] ), .ZN(_08079_ ) );
NAND3_X1 _15782_ ( .A1(_07976_ ), .A2(_07979_ ), .A3(\RFU.rf[9][19] ), .ZN(_08080_ ) );
BUF_X4 _15783_ ( .A(_07973_ ), .Z(_08081_ ) );
NAND3_X1 _15784_ ( .A1(_08081_ ), .A2(\RFU.rf[1][19] ), .A3(_07983_ ), .ZN(_08082_ ) );
NAND3_X1 _15785_ ( .A1(_07986_ ), .A2(_07988_ ), .A3(\RFU.rf[12][19] ), .ZN(_08083_ ) );
AND4_X1 _15786_ ( .A1(_08079_ ), .A2(_08080_ ), .A3(_08082_ ), .A4(_08083_ ), .ZN(_08084_ ) );
NAND3_X1 _15787_ ( .A1(_07992_ ), .A2(\RFU.rf[13][19] ), .A3(_07993_ ), .ZN(_08085_ ) );
BUF_X4 _15788_ ( .A(_07997_ ), .Z(_08086_ ) );
NAND3_X1 _15789_ ( .A1(_07996_ ), .A2(\RFU.rf[10][19] ), .A3(_08086_ ), .ZN(_08087_ ) );
NAND3_X1 _15790_ ( .A1(_08000_ ), .A2(\RFU.rf[8][19] ), .A3(_08001_ ), .ZN(_08088_ ) );
NAND3_X1 _15791_ ( .A1(_08003_ ), .A2(\RFU.rf[11][19] ), .A3(_08004_ ), .ZN(_08089_ ) );
AND4_X1 _15792_ ( .A1(_08085_ ), .A2(_08087_ ), .A3(_08088_ ), .A4(_08089_ ), .ZN(_08090_ ) );
NAND3_X1 _15793_ ( .A1(_08078_ ), .A2(_08084_ ), .A3(_08090_ ), .ZN(_08091_ ) );
MUX2_X1 _15794_ ( .A(\EXU.r1_i [19] ), .B(_08091_ ), .S(_08048_ ), .Z(_00675_ ) );
NAND3_X1 _15795_ ( .A1(_07937_ ), .A2(\RFU.rf[14][18] ), .A3(_07940_ ), .ZN(_08092_ ) );
NAND3_X1 _15796_ ( .A1(_07945_ ), .A2(\RFU.rf[4][18] ), .A3(_07947_ ), .ZN(_08093_ ) );
NAND3_X1 _15797_ ( .A1(_07949_ ), .A2(\RFU.rf[7][18] ), .A3(_07952_ ), .ZN(_08094_ ) );
BUF_X4 _15798_ ( .A(_07939_ ), .Z(_08095_ ) );
NAND3_X1 _15799_ ( .A1(_08095_ ), .A2(_07956_ ), .A3(\RFU.rf[15][18] ), .ZN(_08096_ ) );
NAND4_X1 _15800_ ( .A1(_08092_ ), .A2(_08093_ ), .A3(_08094_ ), .A4(_08096_ ), .ZN(_08097_ ) );
CLKBUF_X2 _15801_ ( .A(_07936_ ), .Z(_08098_ ) );
AND3_X1 _15802_ ( .A1(_08098_ ), .A2(\RFU.rf[2][18] ), .A3(_07961_ ), .ZN(_08099_ ) );
CLKBUF_X2 _15803_ ( .A(_07944_ ), .Z(_08100_ ) );
AND3_X1 _15804_ ( .A1(_08100_ ), .A2(_08075_ ), .A3(\RFU.rf[6][18] ), .ZN(_08101_ ) );
CLKBUF_X2 _15805_ ( .A(_07955_ ), .Z(_08102_ ) );
CLKBUF_X2 _15806_ ( .A(_07960_ ), .Z(_08103_ ) );
AND3_X1 _15807_ ( .A1(_08102_ ), .A2(\RFU.rf[3][18] ), .A3(_08103_ ), .ZN(_08104_ ) );
NOR4_X1 _15808_ ( .A1(_08097_ ), .A2(_08099_ ), .A3(_08101_ ), .A4(_08104_ ), .ZN(_08105_ ) );
NAND3_X1 _15809_ ( .A1(_07971_ ), .A2(_07974_ ), .A3(\RFU.rf[5][18] ), .ZN(_08106_ ) );
NAND3_X1 _15810_ ( .A1(_07976_ ), .A2(_07979_ ), .A3(\RFU.rf[9][18] ), .ZN(_08107_ ) );
NAND3_X1 _15811_ ( .A1(_08081_ ), .A2(\RFU.rf[1][18] ), .A3(_07983_ ), .ZN(_08108_ ) );
NAND3_X1 _15812_ ( .A1(_07986_ ), .A2(_07988_ ), .A3(\RFU.rf[12][18] ), .ZN(_08109_ ) );
AND4_X1 _15813_ ( .A1(_08106_ ), .A2(_08107_ ), .A3(_08108_ ), .A4(_08109_ ), .ZN(_08110_ ) );
NAND3_X1 _15814_ ( .A1(_07992_ ), .A2(\RFU.rf[13][18] ), .A3(_07993_ ), .ZN(_08111_ ) );
NAND3_X1 _15815_ ( .A1(_07996_ ), .A2(\RFU.rf[10][18] ), .A3(_08086_ ), .ZN(_08112_ ) );
NAND3_X1 _15816_ ( .A1(_08000_ ), .A2(\RFU.rf[8][18] ), .A3(_08001_ ), .ZN(_08113_ ) );
NAND3_X1 _15817_ ( .A1(_08003_ ), .A2(\RFU.rf[11][18] ), .A3(_08004_ ), .ZN(_08114_ ) );
AND4_X1 _15818_ ( .A1(_08111_ ), .A2(_08112_ ), .A3(_08113_ ), .A4(_08114_ ), .ZN(_08115_ ) );
NAND3_X1 _15819_ ( .A1(_08105_ ), .A2(_08110_ ), .A3(_08115_ ), .ZN(_08116_ ) );
MUX2_X1 _15820_ ( .A(\EXU.r1_i [18] ), .B(_08116_ ), .S(_08048_ ), .Z(_00676_ ) );
BUF_X4 _15821_ ( .A(_07936_ ), .Z(_08117_ ) );
BUF_X4 _15822_ ( .A(_07939_ ), .Z(_08118_ ) );
NAND3_X1 _15823_ ( .A1(_08117_ ), .A2(\RFU.rf[14][17] ), .A3(_08118_ ), .ZN(_08119_ ) );
BUF_X4 _15824_ ( .A(_07946_ ), .Z(_08120_ ) );
NAND3_X1 _15825_ ( .A1(_07945_ ), .A2(\RFU.rf[4][17] ), .A3(_08120_ ), .ZN(_08121_ ) );
BUF_X4 _15826_ ( .A(_07944_ ), .Z(_08122_ ) );
NAND3_X1 _15827_ ( .A1(_08122_ ), .A2(\RFU.rf[7][17] ), .A3(_07952_ ), .ZN(_08123_ ) );
BUF_X4 _15828_ ( .A(_07955_ ), .Z(_08124_ ) );
NAND3_X1 _15829_ ( .A1(_08095_ ), .A2(_08124_ ), .A3(\RFU.rf[15][17] ), .ZN(_08125_ ) );
NAND4_X1 _15830_ ( .A1(_08119_ ), .A2(_08121_ ), .A3(_08123_ ), .A4(_08125_ ), .ZN(_08126_ ) );
CLKBUF_X2 _15831_ ( .A(_07982_ ), .Z(_08127_ ) );
AND3_X1 _15832_ ( .A1(_08098_ ), .A2(\RFU.rf[2][17] ), .A3(_08127_ ), .ZN(_08128_ ) );
AND3_X1 _15833_ ( .A1(_08100_ ), .A2(_08075_ ), .A3(\RFU.rf[6][17] ), .ZN(_08129_ ) );
AND3_X1 _15834_ ( .A1(_08102_ ), .A2(\RFU.rf[3][17] ), .A3(_08103_ ), .ZN(_08130_ ) );
NOR4_X1 _15835_ ( .A1(_08126_ ), .A2(_08128_ ), .A3(_08129_ ), .A4(_08130_ ), .ZN(_08131_ ) );
NAND3_X1 _15836_ ( .A1(_07971_ ), .A2(_07974_ ), .A3(\RFU.rf[5][17] ), .ZN(_08132_ ) );
BUF_X4 _15837_ ( .A(_07973_ ), .Z(_08133_ ) );
NAND3_X1 _15838_ ( .A1(_08133_ ), .A2(_07979_ ), .A3(\RFU.rf[9][17] ), .ZN(_08134_ ) );
NAND3_X1 _15839_ ( .A1(_08081_ ), .A2(\RFU.rf[1][17] ), .A3(_07983_ ), .ZN(_08135_ ) );
NAND3_X1 _15840_ ( .A1(_07986_ ), .A2(_07988_ ), .A3(\RFU.rf[12][17] ), .ZN(_08136_ ) );
AND4_X1 _15841_ ( .A1(_08132_ ), .A2(_08134_ ), .A3(_08135_ ), .A4(_08136_ ), .ZN(_08137_ ) );
NAND3_X1 _15842_ ( .A1(_07992_ ), .A2(\RFU.rf[13][17] ), .A3(_07993_ ), .ZN(_08138_ ) );
NAND3_X1 _15843_ ( .A1(_07996_ ), .A2(\RFU.rf[10][17] ), .A3(_08086_ ), .ZN(_08139_ ) );
NAND3_X1 _15844_ ( .A1(_08000_ ), .A2(\RFU.rf[8][17] ), .A3(_08001_ ), .ZN(_08140_ ) );
BUF_X4 _15845_ ( .A(_07997_ ), .Z(_08141_ ) );
NAND3_X1 _15846_ ( .A1(_08141_ ), .A2(\RFU.rf[11][17] ), .A3(_08004_ ), .ZN(_08142_ ) );
AND4_X1 _15847_ ( .A1(_08138_ ), .A2(_08139_ ), .A3(_08140_ ), .A4(_08142_ ), .ZN(_08143_ ) );
NAND3_X1 _15848_ ( .A1(_08131_ ), .A2(_08137_ ), .A3(_08143_ ), .ZN(_08144_ ) );
MUX2_X1 _15849_ ( .A(\EXU.r1_i [17] ), .B(_08144_ ), .S(_08048_ ), .Z(_00677_ ) );
NAND3_X1 _15850_ ( .A1(_08117_ ), .A2(\RFU.rf[14][16] ), .A3(_08118_ ), .ZN(_08145_ ) );
BUF_X4 _15851_ ( .A(_07944_ ), .Z(_08146_ ) );
NAND3_X1 _15852_ ( .A1(_08146_ ), .A2(\RFU.rf[4][16] ), .A3(_08120_ ), .ZN(_08147_ ) );
BUF_X4 _15853_ ( .A(_07955_ ), .Z(_08148_ ) );
NAND3_X1 _15854_ ( .A1(_08122_ ), .A2(\RFU.rf[7][16] ), .A3(_08148_ ), .ZN(_08149_ ) );
NAND3_X1 _15855_ ( .A1(_08095_ ), .A2(_08124_ ), .A3(\RFU.rf[15][16] ), .ZN(_08150_ ) );
NAND4_X1 _15856_ ( .A1(_08145_ ), .A2(_08147_ ), .A3(_08149_ ), .A4(_08150_ ), .ZN(_08151_ ) );
AND3_X1 _15857_ ( .A1(_08098_ ), .A2(\RFU.rf[2][16] ), .A3(_08127_ ), .ZN(_08152_ ) );
AND3_X1 _15858_ ( .A1(_08100_ ), .A2(_08075_ ), .A3(\RFU.rf[6][16] ), .ZN(_08153_ ) );
AND3_X1 _15859_ ( .A1(_08102_ ), .A2(\RFU.rf[3][16] ), .A3(_08103_ ), .ZN(_08154_ ) );
NOR4_X1 _15860_ ( .A1(_08151_ ), .A2(_08152_ ), .A3(_08153_ ), .A4(_08154_ ), .ZN(_08155_ ) );
NAND3_X1 _15861_ ( .A1(_07971_ ), .A2(_07974_ ), .A3(\RFU.rf[5][16] ), .ZN(_08156_ ) );
NAND3_X1 _15862_ ( .A1(_08133_ ), .A2(_07979_ ), .A3(\RFU.rf[9][16] ), .ZN(_08157_ ) );
NAND3_X1 _15863_ ( .A1(_08081_ ), .A2(\RFU.rf[1][16] ), .A3(_07983_ ), .ZN(_08158_ ) );
NAND3_X1 _15864_ ( .A1(_07986_ ), .A2(_07988_ ), .A3(\RFU.rf[12][16] ), .ZN(_08159_ ) );
AND4_X1 _15865_ ( .A1(_08156_ ), .A2(_08157_ ), .A3(_08158_ ), .A4(_08159_ ), .ZN(_08160_ ) );
NAND3_X1 _15866_ ( .A1(_07992_ ), .A2(\RFU.rf[13][16] ), .A3(_07993_ ), .ZN(_08161_ ) );
NAND3_X1 _15867_ ( .A1(_07996_ ), .A2(\RFU.rf[10][16] ), .A3(_08086_ ), .ZN(_08162_ ) );
NAND3_X1 _15868_ ( .A1(_08000_ ), .A2(\RFU.rf[8][16] ), .A3(_08001_ ), .ZN(_08163_ ) );
NAND3_X1 _15869_ ( .A1(_08141_ ), .A2(\RFU.rf[11][16] ), .A3(_08004_ ), .ZN(_08164_ ) );
AND4_X1 _15870_ ( .A1(_08161_ ), .A2(_08162_ ), .A3(_08163_ ), .A4(_08164_ ), .ZN(_08165_ ) );
NAND3_X1 _15871_ ( .A1(_08155_ ), .A2(_08160_ ), .A3(_08165_ ), .ZN(_08166_ ) );
MUX2_X1 _15872_ ( .A(\EXU.r1_i [16] ), .B(_08166_ ), .S(_08048_ ), .Z(_00678_ ) );
NAND3_X1 _15873_ ( .A1(_08117_ ), .A2(\RFU.rf[14][15] ), .A3(_08118_ ), .ZN(_08167_ ) );
NAND3_X1 _15874_ ( .A1(_08146_ ), .A2(\RFU.rf[4][15] ), .A3(_08120_ ), .ZN(_08168_ ) );
NAND3_X1 _15875_ ( .A1(_08122_ ), .A2(\RFU.rf[7][15] ), .A3(_08148_ ), .ZN(_08169_ ) );
NAND3_X1 _15876_ ( .A1(_08095_ ), .A2(_08124_ ), .A3(\RFU.rf[15][15] ), .ZN(_08170_ ) );
NAND4_X1 _15877_ ( .A1(_08167_ ), .A2(_08168_ ), .A3(_08169_ ), .A4(_08170_ ), .ZN(_08171_ ) );
AND3_X1 _15878_ ( .A1(_08098_ ), .A2(\RFU.rf[2][15] ), .A3(_08127_ ), .ZN(_08172_ ) );
AND3_X1 _15879_ ( .A1(_08100_ ), .A2(_08075_ ), .A3(\RFU.rf[6][15] ), .ZN(_08173_ ) );
AND3_X1 _15880_ ( .A1(_08102_ ), .A2(\RFU.rf[3][15] ), .A3(_08103_ ), .ZN(_08174_ ) );
NOR4_X1 _15881_ ( .A1(_08171_ ), .A2(_08172_ ), .A3(_08173_ ), .A4(_08174_ ), .ZN(_08175_ ) );
BUF_X4 _15882_ ( .A(_07973_ ), .Z(_08176_ ) );
NAND3_X1 _15883_ ( .A1(_07971_ ), .A2(_08176_ ), .A3(\RFU.rf[5][15] ), .ZN(_08177_ ) );
NAND3_X1 _15884_ ( .A1(_08133_ ), .A2(_07979_ ), .A3(\RFU.rf[9][15] ), .ZN(_08178_ ) );
BUF_X4 _15885_ ( .A(_07982_ ), .Z(_08179_ ) );
NAND3_X1 _15886_ ( .A1(_08081_ ), .A2(\RFU.rf[1][15] ), .A3(_08179_ ), .ZN(_08180_ ) );
BUF_X4 _15887_ ( .A(_07939_ ), .Z(_08181_ ) );
NAND3_X1 _15888_ ( .A1(_08181_ ), .A2(_07988_ ), .A3(\RFU.rf[12][15] ), .ZN(_08182_ ) );
AND4_X1 _15889_ ( .A1(_08177_ ), .A2(_08178_ ), .A3(_08180_ ), .A4(_08182_ ), .ZN(_08183_ ) );
NAND3_X1 _15890_ ( .A1(_07992_ ), .A2(\RFU.rf[13][15] ), .A3(_07993_ ), .ZN(_08184_ ) );
NAND3_X1 _15891_ ( .A1(_07996_ ), .A2(\RFU.rf[10][15] ), .A3(_08086_ ), .ZN(_08185_ ) );
BUF_X4 _15892_ ( .A(_07997_ ), .Z(_08186_ ) );
BUF_X4 _15893_ ( .A(_07987_ ), .Z(_08187_ ) );
NAND3_X1 _15894_ ( .A1(_08186_ ), .A2(\RFU.rf[8][15] ), .A3(_08187_ ), .ZN(_08188_ ) );
NAND3_X1 _15895_ ( .A1(_08141_ ), .A2(\RFU.rf[11][15] ), .A3(_08004_ ), .ZN(_08189_ ) );
AND4_X1 _15896_ ( .A1(_08184_ ), .A2(_08185_ ), .A3(_08188_ ), .A4(_08189_ ), .ZN(_08190_ ) );
NAND3_X1 _15897_ ( .A1(_08175_ ), .A2(_08183_ ), .A3(_08190_ ), .ZN(_08191_ ) );
MUX2_X1 _15898_ ( .A(\EXU.r1_i [15] ), .B(_08191_ ), .S(_08048_ ), .Z(_00679_ ) );
NAND3_X1 _15899_ ( .A1(_08117_ ), .A2(\RFU.rf[14][14] ), .A3(_08118_ ), .ZN(_08192_ ) );
NAND3_X1 _15900_ ( .A1(_08146_ ), .A2(\RFU.rf[4][14] ), .A3(_08120_ ), .ZN(_08193_ ) );
NAND3_X1 _15901_ ( .A1(_08122_ ), .A2(\RFU.rf[7][14] ), .A3(_08148_ ), .ZN(_08194_ ) );
NAND3_X1 _15902_ ( .A1(_08095_ ), .A2(_08124_ ), .A3(\RFU.rf[15][14] ), .ZN(_08195_ ) );
NAND4_X1 _15903_ ( .A1(_08192_ ), .A2(_08193_ ), .A3(_08194_ ), .A4(_08195_ ), .ZN(_08196_ ) );
AND3_X1 _15904_ ( .A1(_08098_ ), .A2(\RFU.rf[2][14] ), .A3(_08127_ ), .ZN(_08197_ ) );
AND3_X1 _15905_ ( .A1(_08100_ ), .A2(_08075_ ), .A3(\RFU.rf[6][14] ), .ZN(_08198_ ) );
AND3_X1 _15906_ ( .A1(_08102_ ), .A2(\RFU.rf[3][14] ), .A3(_08103_ ), .ZN(_08199_ ) );
NOR4_X1 _15907_ ( .A1(_08196_ ), .A2(_08197_ ), .A3(_08198_ ), .A4(_08199_ ), .ZN(_08200_ ) );
NAND3_X1 _15908_ ( .A1(_07971_ ), .A2(_08176_ ), .A3(\RFU.rf[5][14] ), .ZN(_08201_ ) );
NAND3_X1 _15909_ ( .A1(_08133_ ), .A2(_07979_ ), .A3(\RFU.rf[9][14] ), .ZN(_08202_ ) );
NAND3_X1 _15910_ ( .A1(_08081_ ), .A2(\RFU.rf[1][14] ), .A3(_08179_ ), .ZN(_08203_ ) );
NAND3_X1 _15911_ ( .A1(_08181_ ), .A2(_07988_ ), .A3(\RFU.rf[12][14] ), .ZN(_08204_ ) );
AND4_X1 _15912_ ( .A1(_08201_ ), .A2(_08202_ ), .A3(_08203_ ), .A4(_08204_ ), .ZN(_08205_ ) );
NAND3_X1 _15913_ ( .A1(_07992_ ), .A2(\RFU.rf[13][14] ), .A3(_07993_ ), .ZN(_08206_ ) );
BUF_X4 _15914_ ( .A(_07995_ ), .Z(_08207_ ) );
NAND3_X1 _15915_ ( .A1(_08207_ ), .A2(\RFU.rf[10][14] ), .A3(_08086_ ), .ZN(_08208_ ) );
NAND3_X1 _15916_ ( .A1(_08186_ ), .A2(\RFU.rf[8][14] ), .A3(_08187_ ), .ZN(_08209_ ) );
BUF_X4 _15917_ ( .A(_07951_ ), .Z(_08210_ ) );
NAND3_X1 _15918_ ( .A1(_08141_ ), .A2(\RFU.rf[11][14] ), .A3(_08210_ ), .ZN(_08211_ ) );
AND4_X1 _15919_ ( .A1(_08206_ ), .A2(_08208_ ), .A3(_08209_ ), .A4(_08211_ ), .ZN(_08212_ ) );
NAND3_X1 _15920_ ( .A1(_08200_ ), .A2(_08205_ ), .A3(_08212_ ), .ZN(_08213_ ) );
MUX2_X1 _15921_ ( .A(\EXU.r1_i [14] ), .B(_08213_ ), .S(_08048_ ), .Z(_00680_ ) );
NAND3_X1 _15922_ ( .A1(_07996_ ), .A2(\RFU.rf[2][13] ), .A3(_07983_ ), .ZN(_08214_ ) );
NAND3_X1 _15923_ ( .A1(_07970_ ), .A2(\RFU.rf[4][13] ), .A3(_07946_ ), .ZN(_08215_ ) );
NAND3_X1 _15924_ ( .A1(_07936_ ), .A2(\RFU.rf[14][13] ), .A3(_07939_ ), .ZN(_08216_ ) );
NAND3_X1 _15925_ ( .A1(_07944_ ), .A2(\RFU.rf[7][13] ), .A3(_07955_ ), .ZN(_08217_ ) );
NAND3_X1 _15926_ ( .A1(_07939_ ), .A2(_07955_ ), .A3(\RFU.rf[15][13] ), .ZN(_08218_ ) );
AND4_X1 _15927_ ( .A1(_08215_ ), .A2(_08216_ ), .A3(_08217_ ), .A4(_08218_ ), .ZN(_08219_ ) );
NAND3_X1 _15928_ ( .A1(_07945_ ), .A2(_07937_ ), .A3(\RFU.rf[6][13] ), .ZN(_08220_ ) );
NAND3_X1 _15929_ ( .A1(_08004_ ), .A2(_07983_ ), .A3(\RFU.rf[3][13] ), .ZN(_08221_ ) );
AND4_X1 _15930_ ( .A1(_08214_ ), .A2(_08219_ ), .A3(_08220_ ), .A4(_08221_ ), .ZN(_08222_ ) );
BUF_X4 _15931_ ( .A(_07970_ ), .Z(_08223_ ) );
NAND3_X1 _15932_ ( .A1(_08223_ ), .A2(_08176_ ), .A3(\RFU.rf[5][13] ), .ZN(_08224_ ) );
BUF_X4 _15933_ ( .A(_07978_ ), .Z(_08225_ ) );
NAND3_X1 _15934_ ( .A1(_08133_ ), .A2(_08225_ ), .A3(\RFU.rf[9][13] ), .ZN(_08226_ ) );
NAND3_X1 _15935_ ( .A1(_08081_ ), .A2(\RFU.rf[1][13] ), .A3(_08179_ ), .ZN(_08227_ ) );
BUF_X4 _15936_ ( .A(_07987_ ), .Z(_08228_ ) );
NAND3_X1 _15937_ ( .A1(_08181_ ), .A2(_08228_ ), .A3(\RFU.rf[12][13] ), .ZN(_08229_ ) );
AND4_X1 _15938_ ( .A1(_08224_ ), .A2(_08226_ ), .A3(_08227_ ), .A4(_08229_ ), .ZN(_08230_ ) );
BUF_X4 _15939_ ( .A(_07991_ ), .Z(_08231_ ) );
BUF_X4 _15940_ ( .A(_07985_ ), .Z(_08232_ ) );
NAND3_X1 _15941_ ( .A1(_08231_ ), .A2(\RFU.rf[13][13] ), .A3(_08232_ ), .ZN(_08233_ ) );
NAND3_X1 _15942_ ( .A1(_08207_ ), .A2(\RFU.rf[10][13] ), .A3(_08086_ ), .ZN(_08234_ ) );
NAND3_X1 _15943_ ( .A1(_08186_ ), .A2(\RFU.rf[8][13] ), .A3(_08187_ ), .ZN(_08235_ ) );
NAND3_X1 _15944_ ( .A1(_08141_ ), .A2(\RFU.rf[11][13] ), .A3(_08210_ ), .ZN(_08236_ ) );
AND4_X1 _15945_ ( .A1(_08233_ ), .A2(_08234_ ), .A3(_08235_ ), .A4(_08236_ ), .ZN(_08237_ ) );
NAND3_X1 _15946_ ( .A1(_08222_ ), .A2(_08230_ ), .A3(_08237_ ), .ZN(_08238_ ) );
MUX2_X1 _15947_ ( .A(\EXU.r1_i [13] ), .B(_08238_ ), .S(_08048_ ), .Z(_00681_ ) );
NAND3_X1 _15948_ ( .A1(_08117_ ), .A2(\RFU.rf[14][12] ), .A3(_08118_ ), .ZN(_08239_ ) );
NAND3_X1 _15949_ ( .A1(_08146_ ), .A2(\RFU.rf[4][12] ), .A3(_08120_ ), .ZN(_08240_ ) );
NAND3_X1 _15950_ ( .A1(_08122_ ), .A2(\RFU.rf[7][12] ), .A3(_08148_ ), .ZN(_08241_ ) );
NAND3_X1 _15951_ ( .A1(_08095_ ), .A2(_08124_ ), .A3(\RFU.rf[15][12] ), .ZN(_08242_ ) );
NAND4_X1 _15952_ ( .A1(_08239_ ), .A2(_08240_ ), .A3(_08241_ ), .A4(_08242_ ), .ZN(_08243_ ) );
AND3_X1 _15953_ ( .A1(_08098_ ), .A2(\RFU.rf[2][12] ), .A3(_08127_ ), .ZN(_08244_ ) );
AND3_X1 _15954_ ( .A1(_08100_ ), .A2(_08075_ ), .A3(\RFU.rf[6][12] ), .ZN(_08245_ ) );
AND3_X1 _15955_ ( .A1(_08102_ ), .A2(\RFU.rf[3][12] ), .A3(_08103_ ), .ZN(_08246_ ) );
NOR4_X1 _15956_ ( .A1(_08243_ ), .A2(_08244_ ), .A3(_08245_ ), .A4(_08246_ ), .ZN(_08247_ ) );
NAND3_X1 _15957_ ( .A1(_08223_ ), .A2(_08176_ ), .A3(\RFU.rf[5][12] ), .ZN(_08248_ ) );
NAND3_X1 _15958_ ( .A1(_08133_ ), .A2(_08225_ ), .A3(\RFU.rf[9][12] ), .ZN(_08249_ ) );
NAND3_X1 _15959_ ( .A1(_08081_ ), .A2(\RFU.rf[1][12] ), .A3(_08179_ ), .ZN(_08250_ ) );
NAND3_X1 _15960_ ( .A1(_08181_ ), .A2(_08228_ ), .A3(\RFU.rf[12][12] ), .ZN(_08251_ ) );
AND4_X1 _15961_ ( .A1(_08248_ ), .A2(_08249_ ), .A3(_08250_ ), .A4(_08251_ ), .ZN(_08252_ ) );
NAND3_X1 _15962_ ( .A1(_08231_ ), .A2(\RFU.rf[13][12] ), .A3(_08232_ ), .ZN(_08253_ ) );
NAND3_X1 _15963_ ( .A1(_08207_ ), .A2(\RFU.rf[10][12] ), .A3(_08086_ ), .ZN(_08254_ ) );
NAND3_X1 _15964_ ( .A1(_08186_ ), .A2(\RFU.rf[8][12] ), .A3(_08187_ ), .ZN(_08255_ ) );
NAND3_X1 _15965_ ( .A1(_08141_ ), .A2(\RFU.rf[11][12] ), .A3(_08210_ ), .ZN(_08256_ ) );
AND4_X1 _15966_ ( .A1(_08253_ ), .A2(_08254_ ), .A3(_08255_ ), .A4(_08256_ ), .ZN(_08257_ ) );
NAND3_X1 _15967_ ( .A1(_08247_ ), .A2(_08252_ ), .A3(_08257_ ), .ZN(_08258_ ) );
MUX2_X1 _15968_ ( .A(\EXU.r1_i [12] ), .B(_08258_ ), .S(_08048_ ), .Z(_00682_ ) );
NAND3_X1 _15969_ ( .A1(_08117_ ), .A2(\RFU.rf[14][29] ), .A3(_08118_ ), .ZN(_08259_ ) );
NAND3_X1 _15970_ ( .A1(_08146_ ), .A2(\RFU.rf[4][29] ), .A3(_08120_ ), .ZN(_08260_ ) );
NAND3_X1 _15971_ ( .A1(_08122_ ), .A2(\RFU.rf[7][29] ), .A3(_08148_ ), .ZN(_08261_ ) );
NAND3_X1 _15972_ ( .A1(_08095_ ), .A2(_08124_ ), .A3(\RFU.rf[15][29] ), .ZN(_08262_ ) );
NAND4_X1 _15973_ ( .A1(_08259_ ), .A2(_08260_ ), .A3(_08261_ ), .A4(_08262_ ), .ZN(_08263_ ) );
AND3_X1 _15974_ ( .A1(_08098_ ), .A2(\RFU.rf[2][29] ), .A3(_08127_ ), .ZN(_08264_ ) );
AND3_X1 _15975_ ( .A1(_08100_ ), .A2(_08075_ ), .A3(\RFU.rf[6][29] ), .ZN(_08265_ ) );
AND3_X1 _15976_ ( .A1(_08102_ ), .A2(\RFU.rf[3][29] ), .A3(_08103_ ), .ZN(_08266_ ) );
NOR4_X1 _15977_ ( .A1(_08263_ ), .A2(_08264_ ), .A3(_08265_ ), .A4(_08266_ ), .ZN(_08267_ ) );
NAND3_X1 _15978_ ( .A1(_08223_ ), .A2(_08176_ ), .A3(\RFU.rf[5][29] ), .ZN(_08268_ ) );
NAND3_X1 _15979_ ( .A1(_08133_ ), .A2(_08225_ ), .A3(\RFU.rf[9][29] ), .ZN(_08269_ ) );
NAND3_X1 _15980_ ( .A1(_08081_ ), .A2(\RFU.rf[1][29] ), .A3(_08179_ ), .ZN(_08270_ ) );
NAND3_X1 _15981_ ( .A1(_08181_ ), .A2(_08228_ ), .A3(\RFU.rf[12][29] ), .ZN(_08271_ ) );
AND4_X1 _15982_ ( .A1(_08268_ ), .A2(_08269_ ), .A3(_08270_ ), .A4(_08271_ ), .ZN(_08272_ ) );
NAND3_X1 _15983_ ( .A1(_08231_ ), .A2(\RFU.rf[13][29] ), .A3(_08232_ ), .ZN(_08273_ ) );
NAND3_X1 _15984_ ( .A1(_08207_ ), .A2(\RFU.rf[10][29] ), .A3(_08086_ ), .ZN(_08274_ ) );
NAND3_X1 _15985_ ( .A1(_08186_ ), .A2(\RFU.rf[8][29] ), .A3(_08187_ ), .ZN(_08275_ ) );
NAND3_X1 _15986_ ( .A1(_08141_ ), .A2(\RFU.rf[11][29] ), .A3(_08210_ ), .ZN(_08276_ ) );
AND4_X1 _15987_ ( .A1(_08273_ ), .A2(_08274_ ), .A3(_08275_ ), .A4(_08276_ ), .ZN(_08277_ ) );
NAND3_X1 _15988_ ( .A1(_08267_ ), .A2(_08272_ ), .A3(_08277_ ), .ZN(_08278_ ) );
BUF_X4 _15989_ ( .A(_05514_ ), .Z(_08279_ ) );
MUX2_X1 _15990_ ( .A(\EXU.r1_i [29] ), .B(_08278_ ), .S(_08279_ ), .Z(_00683_ ) );
NAND3_X1 _15991_ ( .A1(_08117_ ), .A2(\RFU.rf[14][11] ), .A3(_08118_ ), .ZN(_08280_ ) );
NAND3_X1 _15992_ ( .A1(_08146_ ), .A2(\RFU.rf[4][11] ), .A3(_08120_ ), .ZN(_08281_ ) );
NAND3_X1 _15993_ ( .A1(_08122_ ), .A2(\RFU.rf[7][11] ), .A3(_08148_ ), .ZN(_08282_ ) );
NAND3_X1 _15994_ ( .A1(_08095_ ), .A2(_08124_ ), .A3(\RFU.rf[15][11] ), .ZN(_08283_ ) );
NAND4_X1 _15995_ ( .A1(_08280_ ), .A2(_08281_ ), .A3(_08282_ ), .A4(_08283_ ), .ZN(_08284_ ) );
AND3_X1 _15996_ ( .A1(_08098_ ), .A2(\RFU.rf[2][11] ), .A3(_08127_ ), .ZN(_08285_ ) );
AND3_X1 _15997_ ( .A1(_08100_ ), .A2(_08075_ ), .A3(\RFU.rf[6][11] ), .ZN(_08286_ ) );
AND3_X1 _15998_ ( .A1(_08102_ ), .A2(\RFU.rf[3][11] ), .A3(_08103_ ), .ZN(_08287_ ) );
NOR4_X1 _15999_ ( .A1(_08284_ ), .A2(_08285_ ), .A3(_08286_ ), .A4(_08287_ ), .ZN(_08288_ ) );
NAND3_X1 _16000_ ( .A1(_08223_ ), .A2(_08176_ ), .A3(\RFU.rf[5][11] ), .ZN(_08289_ ) );
NAND3_X1 _16001_ ( .A1(_08133_ ), .A2(_08225_ ), .A3(\RFU.rf[9][11] ), .ZN(_08290_ ) );
NAND3_X1 _16002_ ( .A1(_08081_ ), .A2(\RFU.rf[1][11] ), .A3(_08179_ ), .ZN(_08291_ ) );
NAND3_X1 _16003_ ( .A1(_08181_ ), .A2(_08228_ ), .A3(\RFU.rf[12][11] ), .ZN(_08292_ ) );
AND4_X1 _16004_ ( .A1(_08289_ ), .A2(_08290_ ), .A3(_08291_ ), .A4(_08292_ ), .ZN(_08293_ ) );
NAND3_X1 _16005_ ( .A1(_08231_ ), .A2(\RFU.rf[13][11] ), .A3(_08232_ ), .ZN(_08294_ ) );
NAND3_X1 _16006_ ( .A1(_08207_ ), .A2(\RFU.rf[10][11] ), .A3(_08086_ ), .ZN(_08295_ ) );
NAND3_X1 _16007_ ( .A1(_08186_ ), .A2(\RFU.rf[8][11] ), .A3(_08187_ ), .ZN(_08296_ ) );
NAND3_X1 _16008_ ( .A1(_08141_ ), .A2(\RFU.rf[11][11] ), .A3(_08210_ ), .ZN(_08297_ ) );
AND4_X1 _16009_ ( .A1(_08294_ ), .A2(_08295_ ), .A3(_08296_ ), .A4(_08297_ ), .ZN(_08298_ ) );
NAND3_X1 _16010_ ( .A1(_08288_ ), .A2(_08293_ ), .A3(_08298_ ), .ZN(_08299_ ) );
MUX2_X1 _16011_ ( .A(\EXU.r1_i [11] ), .B(_08299_ ), .S(_08279_ ), .Z(_00684_ ) );
NAND3_X1 _16012_ ( .A1(_08117_ ), .A2(\RFU.rf[14][10] ), .A3(_08118_ ), .ZN(_08300_ ) );
NAND3_X1 _16013_ ( .A1(_08146_ ), .A2(\RFU.rf[4][10] ), .A3(_08120_ ), .ZN(_08301_ ) );
NAND3_X1 _16014_ ( .A1(_08122_ ), .A2(\RFU.rf[7][10] ), .A3(_08148_ ), .ZN(_08302_ ) );
NAND3_X1 _16015_ ( .A1(_08095_ ), .A2(_08124_ ), .A3(\RFU.rf[15][10] ), .ZN(_08303_ ) );
NAND4_X1 _16016_ ( .A1(_08300_ ), .A2(_08301_ ), .A3(_08302_ ), .A4(_08303_ ), .ZN(_08304_ ) );
AND3_X1 _16017_ ( .A1(_08098_ ), .A2(\RFU.rf[2][10] ), .A3(_08127_ ), .ZN(_08305_ ) );
AND3_X1 _16018_ ( .A1(_08100_ ), .A2(_08075_ ), .A3(\RFU.rf[6][10] ), .ZN(_08306_ ) );
AND3_X1 _16019_ ( .A1(_08102_ ), .A2(\RFU.rf[3][10] ), .A3(_08103_ ), .ZN(_08307_ ) );
NOR4_X1 _16020_ ( .A1(_08304_ ), .A2(_08305_ ), .A3(_08306_ ), .A4(_08307_ ), .ZN(_08308_ ) );
NAND3_X1 _16021_ ( .A1(_08223_ ), .A2(_08176_ ), .A3(\RFU.rf[5][10] ), .ZN(_08309_ ) );
NAND3_X1 _16022_ ( .A1(_08133_ ), .A2(_08225_ ), .A3(\RFU.rf[9][10] ), .ZN(_08310_ ) );
BUF_X4 _16023_ ( .A(_07973_ ), .Z(_08311_ ) );
NAND3_X1 _16024_ ( .A1(_08311_ ), .A2(\RFU.rf[1][10] ), .A3(_08179_ ), .ZN(_08312_ ) );
NAND3_X1 _16025_ ( .A1(_08181_ ), .A2(_08228_ ), .A3(\RFU.rf[12][10] ), .ZN(_08313_ ) );
AND4_X1 _16026_ ( .A1(_08309_ ), .A2(_08310_ ), .A3(_08312_ ), .A4(_08313_ ), .ZN(_08314_ ) );
NAND3_X1 _16027_ ( .A1(_08231_ ), .A2(\RFU.rf[13][10] ), .A3(_08232_ ), .ZN(_08315_ ) );
BUF_X4 _16028_ ( .A(_07997_ ), .Z(_08316_ ) );
NAND3_X1 _16029_ ( .A1(_08207_ ), .A2(\RFU.rf[10][10] ), .A3(_08316_ ), .ZN(_08317_ ) );
NAND3_X1 _16030_ ( .A1(_08186_ ), .A2(\RFU.rf[8][10] ), .A3(_08187_ ), .ZN(_08318_ ) );
NAND3_X1 _16031_ ( .A1(_08141_ ), .A2(\RFU.rf[11][10] ), .A3(_08210_ ), .ZN(_08319_ ) );
AND4_X1 _16032_ ( .A1(_08315_ ), .A2(_08317_ ), .A3(_08318_ ), .A4(_08319_ ), .ZN(_08320_ ) );
NAND3_X1 _16033_ ( .A1(_08308_ ), .A2(_08314_ ), .A3(_08320_ ), .ZN(_08321_ ) );
MUX2_X1 _16034_ ( .A(\EXU.r1_i [10] ), .B(_08321_ ), .S(_08279_ ), .Z(_00685_ ) );
NAND3_X1 _16035_ ( .A1(_08117_ ), .A2(\RFU.rf[14][9] ), .A3(_08118_ ), .ZN(_08322_ ) );
NAND3_X1 _16036_ ( .A1(_08146_ ), .A2(\RFU.rf[4][9] ), .A3(_08120_ ), .ZN(_08323_ ) );
NAND3_X1 _16037_ ( .A1(_08122_ ), .A2(\RFU.rf[7][9] ), .A3(_08148_ ), .ZN(_08324_ ) );
NAND3_X1 _16038_ ( .A1(_08095_ ), .A2(_08124_ ), .A3(\RFU.rf[15][9] ), .ZN(_08325_ ) );
NAND4_X1 _16039_ ( .A1(_08322_ ), .A2(_08323_ ), .A3(_08324_ ), .A4(_08325_ ), .ZN(_08326_ ) );
AND3_X1 _16040_ ( .A1(_08098_ ), .A2(\RFU.rf[2][9] ), .A3(_08127_ ), .ZN(_08327_ ) );
CLKBUF_X2 _16041_ ( .A(_07936_ ), .Z(_08328_ ) );
AND3_X1 _16042_ ( .A1(_08100_ ), .A2(_08328_ ), .A3(\RFU.rf[6][9] ), .ZN(_08329_ ) );
AND3_X1 _16043_ ( .A1(_08102_ ), .A2(\RFU.rf[3][9] ), .A3(_08103_ ), .ZN(_08330_ ) );
NOR4_X1 _16044_ ( .A1(_08326_ ), .A2(_08327_ ), .A3(_08329_ ), .A4(_08330_ ), .ZN(_08331_ ) );
NAND3_X1 _16045_ ( .A1(_08223_ ), .A2(_08176_ ), .A3(\RFU.rf[5][9] ), .ZN(_08332_ ) );
NAND3_X1 _16046_ ( .A1(_08133_ ), .A2(_08225_ ), .A3(\RFU.rf[9][9] ), .ZN(_08333_ ) );
NAND3_X1 _16047_ ( .A1(_08311_ ), .A2(\RFU.rf[1][9] ), .A3(_08179_ ), .ZN(_08334_ ) );
NAND3_X1 _16048_ ( .A1(_08181_ ), .A2(_08228_ ), .A3(\RFU.rf[12][9] ), .ZN(_08335_ ) );
AND4_X1 _16049_ ( .A1(_08332_ ), .A2(_08333_ ), .A3(_08334_ ), .A4(_08335_ ), .ZN(_08336_ ) );
NAND3_X1 _16050_ ( .A1(_08231_ ), .A2(\RFU.rf[13][9] ), .A3(_08232_ ), .ZN(_08337_ ) );
NAND3_X1 _16051_ ( .A1(_08207_ ), .A2(\RFU.rf[10][9] ), .A3(_08316_ ), .ZN(_08338_ ) );
NAND3_X1 _16052_ ( .A1(_08186_ ), .A2(\RFU.rf[8][9] ), .A3(_08187_ ), .ZN(_08339_ ) );
NAND3_X1 _16053_ ( .A1(_08141_ ), .A2(\RFU.rf[11][9] ), .A3(_08210_ ), .ZN(_08340_ ) );
AND4_X1 _16054_ ( .A1(_08337_ ), .A2(_08338_ ), .A3(_08339_ ), .A4(_08340_ ), .ZN(_08341_ ) );
NAND3_X1 _16055_ ( .A1(_08331_ ), .A2(_08336_ ), .A3(_08341_ ), .ZN(_08342_ ) );
MUX2_X1 _16056_ ( .A(\EXU.r1_i [9] ), .B(_08342_ ), .S(_08279_ ), .Z(_00686_ ) );
NAND3_X1 _16057_ ( .A1(_08117_ ), .A2(\RFU.rf[14][8] ), .A3(_08118_ ), .ZN(_08343_ ) );
NAND3_X1 _16058_ ( .A1(_08146_ ), .A2(\RFU.rf[4][8] ), .A3(_08120_ ), .ZN(_08344_ ) );
NAND3_X1 _16059_ ( .A1(_08122_ ), .A2(\RFU.rf[7][8] ), .A3(_08148_ ), .ZN(_08345_ ) );
BUF_X4 _16060_ ( .A(_07939_ ), .Z(_08346_ ) );
NAND3_X1 _16061_ ( .A1(_08346_ ), .A2(_08124_ ), .A3(\RFU.rf[15][8] ), .ZN(_08347_ ) );
NAND4_X1 _16062_ ( .A1(_08343_ ), .A2(_08344_ ), .A3(_08345_ ), .A4(_08347_ ), .ZN(_08348_ ) );
CLKBUF_X2 _16063_ ( .A(_07936_ ), .Z(_08349_ ) );
AND3_X1 _16064_ ( .A1(_08349_ ), .A2(\RFU.rf[2][8] ), .A3(_08127_ ), .ZN(_08350_ ) );
CLKBUF_X2 _16065_ ( .A(_07944_ ), .Z(_08351_ ) );
AND3_X1 _16066_ ( .A1(_08351_ ), .A2(_08328_ ), .A3(\RFU.rf[6][8] ), .ZN(_08352_ ) );
CLKBUF_X2 _16067_ ( .A(_07955_ ), .Z(_08353_ ) );
CLKBUF_X2 _16068_ ( .A(_07960_ ), .Z(_08354_ ) );
AND3_X1 _16069_ ( .A1(_08353_ ), .A2(\RFU.rf[3][8] ), .A3(_08354_ ), .ZN(_08355_ ) );
NOR4_X1 _16070_ ( .A1(_08348_ ), .A2(_08350_ ), .A3(_08352_ ), .A4(_08355_ ), .ZN(_08356_ ) );
NAND3_X1 _16071_ ( .A1(_08223_ ), .A2(_08176_ ), .A3(\RFU.rf[5][8] ), .ZN(_08357_ ) );
BUF_X4 _16072_ ( .A(_07973_ ), .Z(_08358_ ) );
NAND3_X1 _16073_ ( .A1(_08358_ ), .A2(_08225_ ), .A3(\RFU.rf[9][8] ), .ZN(_08359_ ) );
NAND3_X1 _16074_ ( .A1(_08311_ ), .A2(\RFU.rf[1][8] ), .A3(_08179_ ), .ZN(_08360_ ) );
NAND3_X1 _16075_ ( .A1(_08181_ ), .A2(_08228_ ), .A3(\RFU.rf[12][8] ), .ZN(_08361_ ) );
AND4_X1 _16076_ ( .A1(_08357_ ), .A2(_08359_ ), .A3(_08360_ ), .A4(_08361_ ), .ZN(_08362_ ) );
NAND3_X1 _16077_ ( .A1(_08231_ ), .A2(\RFU.rf[13][8] ), .A3(_08232_ ), .ZN(_08363_ ) );
NAND3_X1 _16078_ ( .A1(_08207_ ), .A2(\RFU.rf[10][8] ), .A3(_08316_ ), .ZN(_08364_ ) );
NAND3_X1 _16079_ ( .A1(_08186_ ), .A2(\RFU.rf[8][8] ), .A3(_08187_ ), .ZN(_08365_ ) );
BUF_X4 _16080_ ( .A(_07997_ ), .Z(_08366_ ) );
NAND3_X1 _16081_ ( .A1(_08366_ ), .A2(\RFU.rf[11][8] ), .A3(_08210_ ), .ZN(_08367_ ) );
AND4_X1 _16082_ ( .A1(_08363_ ), .A2(_08364_ ), .A3(_08365_ ), .A4(_08367_ ), .ZN(_08368_ ) );
NAND3_X1 _16083_ ( .A1(_08356_ ), .A2(_08362_ ), .A3(_08368_ ), .ZN(_08369_ ) );
MUX2_X1 _16084_ ( .A(\EXU.r1_i [8] ), .B(_08369_ ), .S(_08279_ ), .Z(_00687_ ) );
BUF_X4 _16085_ ( .A(_07936_ ), .Z(_08370_ ) );
BUF_X4 _16086_ ( .A(_07939_ ), .Z(_08371_ ) );
NAND3_X1 _16087_ ( .A1(_08370_ ), .A2(\RFU.rf[14][7] ), .A3(_08371_ ), .ZN(_08372_ ) );
BUF_X4 _16088_ ( .A(_07946_ ), .Z(_08373_ ) );
NAND3_X1 _16089_ ( .A1(_08146_ ), .A2(\RFU.rf[4][7] ), .A3(_08373_ ), .ZN(_08374_ ) );
BUF_X4 _16090_ ( .A(_07944_ ), .Z(_08375_ ) );
NAND3_X1 _16091_ ( .A1(_08375_ ), .A2(\RFU.rf[7][7] ), .A3(_08148_ ), .ZN(_08376_ ) );
BUF_X4 _16092_ ( .A(_07955_ ), .Z(_08377_ ) );
NAND3_X1 _16093_ ( .A1(_08346_ ), .A2(_08377_ ), .A3(\RFU.rf[15][7] ), .ZN(_08378_ ) );
NAND4_X1 _16094_ ( .A1(_08372_ ), .A2(_08374_ ), .A3(_08376_ ), .A4(_08378_ ), .ZN(_08379_ ) );
CLKBUF_X2 _16095_ ( .A(_07960_ ), .Z(_08380_ ) );
AND3_X1 _16096_ ( .A1(_08349_ ), .A2(\RFU.rf[2][7] ), .A3(_08380_ ), .ZN(_08381_ ) );
AND3_X1 _16097_ ( .A1(_08351_ ), .A2(_08328_ ), .A3(\RFU.rf[6][7] ), .ZN(_08382_ ) );
AND3_X1 _16098_ ( .A1(_08353_ ), .A2(\RFU.rf[3][7] ), .A3(_08354_ ), .ZN(_08383_ ) );
NOR4_X1 _16099_ ( .A1(_08379_ ), .A2(_08381_ ), .A3(_08382_ ), .A4(_08383_ ), .ZN(_08384_ ) );
NAND3_X1 _16100_ ( .A1(_08223_ ), .A2(_08176_ ), .A3(\RFU.rf[5][7] ), .ZN(_08385_ ) );
NAND3_X1 _16101_ ( .A1(_08358_ ), .A2(_08225_ ), .A3(\RFU.rf[9][7] ), .ZN(_08386_ ) );
NAND3_X1 _16102_ ( .A1(_08311_ ), .A2(\RFU.rf[1][7] ), .A3(_08179_ ), .ZN(_08387_ ) );
NAND3_X1 _16103_ ( .A1(_08181_ ), .A2(_08228_ ), .A3(\RFU.rf[12][7] ), .ZN(_08388_ ) );
AND4_X1 _16104_ ( .A1(_08385_ ), .A2(_08386_ ), .A3(_08387_ ), .A4(_08388_ ), .ZN(_08389_ ) );
NAND3_X1 _16105_ ( .A1(_08231_ ), .A2(\RFU.rf[13][7] ), .A3(_08232_ ), .ZN(_08390_ ) );
NAND3_X1 _16106_ ( .A1(_08207_ ), .A2(\RFU.rf[10][7] ), .A3(_08316_ ), .ZN(_08391_ ) );
NAND3_X1 _16107_ ( .A1(_08186_ ), .A2(\RFU.rf[8][7] ), .A3(_08187_ ), .ZN(_08392_ ) );
NAND3_X1 _16108_ ( .A1(_08366_ ), .A2(\RFU.rf[11][7] ), .A3(_08210_ ), .ZN(_08393_ ) );
AND4_X1 _16109_ ( .A1(_08390_ ), .A2(_08391_ ), .A3(_08392_ ), .A4(_08393_ ), .ZN(_08394_ ) );
NAND3_X1 _16110_ ( .A1(_08384_ ), .A2(_08389_ ), .A3(_08394_ ), .ZN(_08395_ ) );
MUX2_X1 _16111_ ( .A(\EXU.r1_i [7] ), .B(_08395_ ), .S(_08279_ ), .Z(_00688_ ) );
NAND3_X1 _16112_ ( .A1(_08370_ ), .A2(\RFU.rf[14][6] ), .A3(_08371_ ), .ZN(_08396_ ) );
BUF_X4 _16113_ ( .A(_07944_ ), .Z(_08397_ ) );
NAND3_X1 _16114_ ( .A1(_08397_ ), .A2(\RFU.rf[4][6] ), .A3(_08373_ ), .ZN(_08398_ ) );
BUF_X4 _16115_ ( .A(_07955_ ), .Z(_08399_ ) );
NAND3_X1 _16116_ ( .A1(_08375_ ), .A2(\RFU.rf[7][6] ), .A3(_08399_ ), .ZN(_08400_ ) );
NAND3_X1 _16117_ ( .A1(_08346_ ), .A2(_08377_ ), .A3(\RFU.rf[15][6] ), .ZN(_08401_ ) );
NAND4_X1 _16118_ ( .A1(_08396_ ), .A2(_08398_ ), .A3(_08400_ ), .A4(_08401_ ), .ZN(_08402_ ) );
AND3_X1 _16119_ ( .A1(_08349_ ), .A2(\RFU.rf[2][6] ), .A3(_08380_ ), .ZN(_08403_ ) );
AND3_X1 _16120_ ( .A1(_08351_ ), .A2(_08328_ ), .A3(\RFU.rf[6][6] ), .ZN(_08404_ ) );
AND3_X1 _16121_ ( .A1(_08353_ ), .A2(\RFU.rf[3][6] ), .A3(_08354_ ), .ZN(_08405_ ) );
NOR4_X1 _16122_ ( .A1(_08402_ ), .A2(_08403_ ), .A3(_08404_ ), .A4(_08405_ ), .ZN(_08406_ ) );
BUF_X4 _16123_ ( .A(_07973_ ), .Z(_08407_ ) );
NAND3_X1 _16124_ ( .A1(_08223_ ), .A2(_08407_ ), .A3(\RFU.rf[5][6] ), .ZN(_08408_ ) );
NAND3_X1 _16125_ ( .A1(_08358_ ), .A2(_08225_ ), .A3(\RFU.rf[9][6] ), .ZN(_08409_ ) );
BUF_X4 _16126_ ( .A(_07982_ ), .Z(_08410_ ) );
NAND3_X1 _16127_ ( .A1(_08311_ ), .A2(\RFU.rf[1][6] ), .A3(_08410_ ), .ZN(_08411_ ) );
BUF_X4 _16128_ ( .A(_07939_ ), .Z(_08412_ ) );
NAND3_X1 _16129_ ( .A1(_08412_ ), .A2(_08228_ ), .A3(\RFU.rf[12][6] ), .ZN(_08413_ ) );
AND4_X1 _16130_ ( .A1(_08408_ ), .A2(_08409_ ), .A3(_08411_ ), .A4(_08413_ ), .ZN(_08414_ ) );
NAND3_X1 _16131_ ( .A1(_08231_ ), .A2(\RFU.rf[13][6] ), .A3(_08232_ ), .ZN(_08415_ ) );
NAND3_X1 _16132_ ( .A1(_08207_ ), .A2(\RFU.rf[10][6] ), .A3(_08316_ ), .ZN(_08416_ ) );
BUF_X4 _16133_ ( .A(_07997_ ), .Z(_08417_ ) );
BUF_X4 _16134_ ( .A(_07987_ ), .Z(_08418_ ) );
NAND3_X1 _16135_ ( .A1(_08417_ ), .A2(\RFU.rf[8][6] ), .A3(_08418_ ), .ZN(_08419_ ) );
NAND3_X1 _16136_ ( .A1(_08366_ ), .A2(\RFU.rf[11][6] ), .A3(_08210_ ), .ZN(_08420_ ) );
AND4_X1 _16137_ ( .A1(_08415_ ), .A2(_08416_ ), .A3(_08419_ ), .A4(_08420_ ), .ZN(_08421_ ) );
NAND3_X1 _16138_ ( .A1(_08406_ ), .A2(_08414_ ), .A3(_08421_ ), .ZN(_08422_ ) );
MUX2_X1 _16139_ ( .A(\EXU.r1_i [6] ), .B(_08422_ ), .S(_08279_ ), .Z(_00689_ ) );
NAND3_X1 _16140_ ( .A1(_08370_ ), .A2(\RFU.rf[14][5] ), .A3(_08371_ ), .ZN(_08423_ ) );
NAND3_X1 _16141_ ( .A1(_08397_ ), .A2(\RFU.rf[4][5] ), .A3(_08373_ ), .ZN(_08424_ ) );
NAND3_X1 _16142_ ( .A1(_08375_ ), .A2(\RFU.rf[7][5] ), .A3(_08399_ ), .ZN(_08425_ ) );
NAND3_X1 _16143_ ( .A1(_08346_ ), .A2(_08377_ ), .A3(\RFU.rf[15][5] ), .ZN(_08426_ ) );
NAND4_X1 _16144_ ( .A1(_08423_ ), .A2(_08424_ ), .A3(_08425_ ), .A4(_08426_ ), .ZN(_08427_ ) );
AND3_X1 _16145_ ( .A1(_08349_ ), .A2(\RFU.rf[2][5] ), .A3(_08380_ ), .ZN(_08428_ ) );
AND3_X1 _16146_ ( .A1(_08351_ ), .A2(_08328_ ), .A3(\RFU.rf[6][5] ), .ZN(_08429_ ) );
AND3_X1 _16147_ ( .A1(_08353_ ), .A2(\RFU.rf[3][5] ), .A3(_08354_ ), .ZN(_08430_ ) );
NOR4_X1 _16148_ ( .A1(_08427_ ), .A2(_08428_ ), .A3(_08429_ ), .A4(_08430_ ), .ZN(_08431_ ) );
NAND3_X1 _16149_ ( .A1(_08223_ ), .A2(_08407_ ), .A3(\RFU.rf[5][5] ), .ZN(_08432_ ) );
NAND3_X1 _16150_ ( .A1(_08358_ ), .A2(_08225_ ), .A3(\RFU.rf[9][5] ), .ZN(_08433_ ) );
NAND3_X1 _16151_ ( .A1(_08311_ ), .A2(\RFU.rf[1][5] ), .A3(_08410_ ), .ZN(_08434_ ) );
NAND3_X1 _16152_ ( .A1(_08412_ ), .A2(_08228_ ), .A3(\RFU.rf[12][5] ), .ZN(_08435_ ) );
AND4_X1 _16153_ ( .A1(_08432_ ), .A2(_08433_ ), .A3(_08434_ ), .A4(_08435_ ), .ZN(_08436_ ) );
NAND3_X1 _16154_ ( .A1(_08231_ ), .A2(\RFU.rf[13][5] ), .A3(_08232_ ), .ZN(_08437_ ) );
BUF_X4 _16155_ ( .A(_07995_ ), .Z(_08438_ ) );
NAND3_X1 _16156_ ( .A1(_08438_ ), .A2(\RFU.rf[10][5] ), .A3(_08316_ ), .ZN(_08439_ ) );
NAND3_X1 _16157_ ( .A1(_08417_ ), .A2(\RFU.rf[8][5] ), .A3(_08418_ ), .ZN(_08440_ ) );
BUF_X4 _16158_ ( .A(_07951_ ), .Z(_08441_ ) );
NAND3_X1 _16159_ ( .A1(_08366_ ), .A2(\RFU.rf[11][5] ), .A3(_08441_ ), .ZN(_08442_ ) );
AND4_X1 _16160_ ( .A1(_08437_ ), .A2(_08439_ ), .A3(_08440_ ), .A4(_08442_ ), .ZN(_08443_ ) );
NAND3_X1 _16161_ ( .A1(_08431_ ), .A2(_08436_ ), .A3(_08443_ ), .ZN(_08444_ ) );
MUX2_X1 _16162_ ( .A(\EXU.r1_i [5] ), .B(_08444_ ), .S(_08279_ ), .Z(_00690_ ) );
NAND3_X1 _16163_ ( .A1(_08370_ ), .A2(\RFU.rf[14][4] ), .A3(_08371_ ), .ZN(_08445_ ) );
NAND3_X1 _16164_ ( .A1(_08397_ ), .A2(\RFU.rf[4][4] ), .A3(_08373_ ), .ZN(_08446_ ) );
NAND3_X1 _16165_ ( .A1(_08375_ ), .A2(\RFU.rf[7][4] ), .A3(_08399_ ), .ZN(_08447_ ) );
NAND3_X1 _16166_ ( .A1(_08346_ ), .A2(_08377_ ), .A3(\RFU.rf[15][4] ), .ZN(_08448_ ) );
NAND4_X1 _16167_ ( .A1(_08445_ ), .A2(_08446_ ), .A3(_08447_ ), .A4(_08448_ ), .ZN(_08449_ ) );
AND3_X1 _16168_ ( .A1(_08349_ ), .A2(\RFU.rf[2][4] ), .A3(_08380_ ), .ZN(_08450_ ) );
AND3_X1 _16169_ ( .A1(_08351_ ), .A2(_08328_ ), .A3(\RFU.rf[6][4] ), .ZN(_08451_ ) );
AND3_X1 _16170_ ( .A1(_08353_ ), .A2(\RFU.rf[3][4] ), .A3(_08354_ ), .ZN(_08452_ ) );
NOR4_X1 _16171_ ( .A1(_08449_ ), .A2(_08450_ ), .A3(_08451_ ), .A4(_08452_ ), .ZN(_08453_ ) );
BUF_X4 _16172_ ( .A(_07970_ ), .Z(_08454_ ) );
NAND3_X1 _16173_ ( .A1(_08454_ ), .A2(_08407_ ), .A3(\RFU.rf[5][4] ), .ZN(_08455_ ) );
BUF_X4 _16174_ ( .A(_07997_ ), .Z(_08456_ ) );
NAND3_X1 _16175_ ( .A1(_08358_ ), .A2(_08456_ ), .A3(\RFU.rf[9][4] ), .ZN(_08457_ ) );
NAND3_X1 _16176_ ( .A1(_08311_ ), .A2(\RFU.rf[1][4] ), .A3(_08410_ ), .ZN(_08458_ ) );
BUF_X4 _16177_ ( .A(_07987_ ), .Z(_08459_ ) );
NAND3_X1 _16178_ ( .A1(_08412_ ), .A2(_08459_ ), .A3(\RFU.rf[12][4] ), .ZN(_08460_ ) );
AND4_X1 _16179_ ( .A1(_08455_ ), .A2(_08457_ ), .A3(_08458_ ), .A4(_08460_ ), .ZN(_08461_ ) );
BUF_X4 _16180_ ( .A(_07973_ ), .Z(_08462_ ) );
BUF_X4 _16181_ ( .A(_07985_ ), .Z(_08463_ ) );
NAND3_X1 _16182_ ( .A1(_08462_ ), .A2(\RFU.rf[13][4] ), .A3(_08463_ ), .ZN(_08464_ ) );
NAND3_X1 _16183_ ( .A1(_08438_ ), .A2(\RFU.rf[10][4] ), .A3(_08316_ ), .ZN(_08465_ ) );
NAND3_X1 _16184_ ( .A1(_08417_ ), .A2(\RFU.rf[8][4] ), .A3(_08418_ ), .ZN(_08466_ ) );
NAND3_X1 _16185_ ( .A1(_08366_ ), .A2(\RFU.rf[11][4] ), .A3(_08441_ ), .ZN(_08467_ ) );
AND4_X1 _16186_ ( .A1(_08464_ ), .A2(_08465_ ), .A3(_08466_ ), .A4(_08467_ ), .ZN(_08468_ ) );
NAND3_X1 _16187_ ( .A1(_08453_ ), .A2(_08461_ ), .A3(_08468_ ), .ZN(_08469_ ) );
MUX2_X1 _16188_ ( .A(\EXU.r1_i [4] ), .B(_08469_ ), .S(_08279_ ), .Z(_00691_ ) );
NAND3_X1 _16189_ ( .A1(_08370_ ), .A2(\RFU.rf[14][3] ), .A3(_08371_ ), .ZN(_08470_ ) );
NAND3_X1 _16190_ ( .A1(_08397_ ), .A2(\RFU.rf[4][3] ), .A3(_08373_ ), .ZN(_08471_ ) );
NAND3_X1 _16191_ ( .A1(_08375_ ), .A2(\RFU.rf[7][3] ), .A3(_08399_ ), .ZN(_08472_ ) );
NAND3_X1 _16192_ ( .A1(_08346_ ), .A2(_08377_ ), .A3(\RFU.rf[15][3] ), .ZN(_08473_ ) );
NAND4_X1 _16193_ ( .A1(_08470_ ), .A2(_08471_ ), .A3(_08472_ ), .A4(_08473_ ), .ZN(_08474_ ) );
AND3_X1 _16194_ ( .A1(_08349_ ), .A2(\RFU.rf[2][3] ), .A3(_08380_ ), .ZN(_08475_ ) );
AND3_X1 _16195_ ( .A1(_08351_ ), .A2(_08328_ ), .A3(\RFU.rf[6][3] ), .ZN(_08476_ ) );
AND3_X1 _16196_ ( .A1(_08353_ ), .A2(\RFU.rf[3][3] ), .A3(_08354_ ), .ZN(_08477_ ) );
NOR4_X1 _16197_ ( .A1(_08474_ ), .A2(_08475_ ), .A3(_08476_ ), .A4(_08477_ ), .ZN(_08478_ ) );
NAND3_X1 _16198_ ( .A1(_08454_ ), .A2(_08407_ ), .A3(\RFU.rf[5][3] ), .ZN(_08479_ ) );
NAND3_X1 _16199_ ( .A1(_08358_ ), .A2(_08456_ ), .A3(\RFU.rf[9][3] ), .ZN(_08480_ ) );
NAND3_X1 _16200_ ( .A1(_08311_ ), .A2(\RFU.rf[1][3] ), .A3(_08410_ ), .ZN(_08481_ ) );
NAND3_X1 _16201_ ( .A1(_08412_ ), .A2(_08459_ ), .A3(\RFU.rf[12][3] ), .ZN(_08482_ ) );
AND4_X1 _16202_ ( .A1(_08479_ ), .A2(_08480_ ), .A3(_08481_ ), .A4(_08482_ ), .ZN(_08483_ ) );
NAND3_X1 _16203_ ( .A1(_08462_ ), .A2(\RFU.rf[13][3] ), .A3(_08463_ ), .ZN(_08484_ ) );
NAND3_X1 _16204_ ( .A1(_08438_ ), .A2(\RFU.rf[10][3] ), .A3(_08316_ ), .ZN(_08485_ ) );
NAND3_X1 _16205_ ( .A1(_08417_ ), .A2(\RFU.rf[8][3] ), .A3(_08418_ ), .ZN(_08486_ ) );
NAND3_X1 _16206_ ( .A1(_08366_ ), .A2(\RFU.rf[11][3] ), .A3(_08441_ ), .ZN(_08487_ ) );
AND4_X1 _16207_ ( .A1(_08484_ ), .A2(_08485_ ), .A3(_08486_ ), .A4(_08487_ ), .ZN(_08488_ ) );
NAND3_X1 _16208_ ( .A1(_08478_ ), .A2(_08483_ ), .A3(_08488_ ), .ZN(_08489_ ) );
MUX2_X1 _16209_ ( .A(\EXU.r1_i [3] ), .B(_08489_ ), .S(_08279_ ), .Z(_00692_ ) );
NAND3_X1 _16210_ ( .A1(_08370_ ), .A2(\RFU.rf[14][2] ), .A3(_08371_ ), .ZN(_08490_ ) );
NAND3_X1 _16211_ ( .A1(_08397_ ), .A2(\RFU.rf[4][2] ), .A3(_08373_ ), .ZN(_08491_ ) );
NAND3_X1 _16212_ ( .A1(_08375_ ), .A2(\RFU.rf[7][2] ), .A3(_08399_ ), .ZN(_08492_ ) );
NAND3_X1 _16213_ ( .A1(_08346_ ), .A2(_08377_ ), .A3(\RFU.rf[15][2] ), .ZN(_08493_ ) );
NAND4_X1 _16214_ ( .A1(_08490_ ), .A2(_08491_ ), .A3(_08492_ ), .A4(_08493_ ), .ZN(_08494_ ) );
AND3_X1 _16215_ ( .A1(_08349_ ), .A2(\RFU.rf[2][2] ), .A3(_08380_ ), .ZN(_08495_ ) );
AND3_X1 _16216_ ( .A1(_08351_ ), .A2(_08328_ ), .A3(\RFU.rf[6][2] ), .ZN(_08496_ ) );
AND3_X1 _16217_ ( .A1(_08353_ ), .A2(\RFU.rf[3][2] ), .A3(_08354_ ), .ZN(_08497_ ) );
NOR4_X1 _16218_ ( .A1(_08494_ ), .A2(_08495_ ), .A3(_08496_ ), .A4(_08497_ ), .ZN(_08498_ ) );
NAND3_X1 _16219_ ( .A1(_08454_ ), .A2(_08407_ ), .A3(\RFU.rf[5][2] ), .ZN(_08499_ ) );
NAND3_X1 _16220_ ( .A1(_08358_ ), .A2(_08456_ ), .A3(\RFU.rf[9][2] ), .ZN(_08500_ ) );
NAND3_X1 _16221_ ( .A1(_08311_ ), .A2(\RFU.rf[1][2] ), .A3(_08410_ ), .ZN(_08501_ ) );
NAND3_X1 _16222_ ( .A1(_08412_ ), .A2(_08459_ ), .A3(\RFU.rf[12][2] ), .ZN(_08502_ ) );
AND4_X1 _16223_ ( .A1(_08499_ ), .A2(_08500_ ), .A3(_08501_ ), .A4(_08502_ ), .ZN(_08503_ ) );
NAND3_X1 _16224_ ( .A1(_08462_ ), .A2(\RFU.rf[13][2] ), .A3(_08463_ ), .ZN(_08504_ ) );
NAND3_X1 _16225_ ( .A1(_08438_ ), .A2(\RFU.rf[10][2] ), .A3(_08316_ ), .ZN(_08505_ ) );
NAND3_X1 _16226_ ( .A1(_08417_ ), .A2(\RFU.rf[8][2] ), .A3(_08418_ ), .ZN(_08506_ ) );
NAND3_X1 _16227_ ( .A1(_08366_ ), .A2(\RFU.rf[11][2] ), .A3(_08441_ ), .ZN(_08507_ ) );
AND4_X1 _16228_ ( .A1(_08504_ ), .A2(_08505_ ), .A3(_08506_ ), .A4(_08507_ ), .ZN(_08508_ ) );
NAND3_X1 _16229_ ( .A1(_08498_ ), .A2(_08503_ ), .A3(_08508_ ), .ZN(_08509_ ) );
BUF_X4 _16230_ ( .A(_05514_ ), .Z(_08510_ ) );
MUX2_X1 _16231_ ( .A(\EXU.r1_i [2] ), .B(_08509_ ), .S(_08510_ ), .Z(_00693_ ) );
NAND3_X1 _16232_ ( .A1(_08370_ ), .A2(\RFU.rf[14][28] ), .A3(_08371_ ), .ZN(_08511_ ) );
NAND3_X1 _16233_ ( .A1(_08397_ ), .A2(\RFU.rf[4][28] ), .A3(_08373_ ), .ZN(_08512_ ) );
NAND3_X1 _16234_ ( .A1(_08375_ ), .A2(\RFU.rf[7][28] ), .A3(_08399_ ), .ZN(_08513_ ) );
NAND3_X1 _16235_ ( .A1(_08346_ ), .A2(_08377_ ), .A3(\RFU.rf[15][28] ), .ZN(_08514_ ) );
NAND4_X1 _16236_ ( .A1(_08511_ ), .A2(_08512_ ), .A3(_08513_ ), .A4(_08514_ ), .ZN(_08515_ ) );
AND3_X1 _16237_ ( .A1(_08349_ ), .A2(\RFU.rf[2][28] ), .A3(_08380_ ), .ZN(_08516_ ) );
AND3_X1 _16238_ ( .A1(_08351_ ), .A2(_08328_ ), .A3(\RFU.rf[6][28] ), .ZN(_08517_ ) );
AND3_X1 _16239_ ( .A1(_08353_ ), .A2(\RFU.rf[3][28] ), .A3(_08354_ ), .ZN(_08518_ ) );
NOR4_X1 _16240_ ( .A1(_08515_ ), .A2(_08516_ ), .A3(_08517_ ), .A4(_08518_ ), .ZN(_08519_ ) );
NAND3_X1 _16241_ ( .A1(_08454_ ), .A2(_08407_ ), .A3(\RFU.rf[5][28] ), .ZN(_08520_ ) );
NAND3_X1 _16242_ ( .A1(_08358_ ), .A2(_08456_ ), .A3(\RFU.rf[9][28] ), .ZN(_08521_ ) );
NAND3_X1 _16243_ ( .A1(_08311_ ), .A2(\RFU.rf[1][28] ), .A3(_08410_ ), .ZN(_08522_ ) );
NAND3_X1 _16244_ ( .A1(_08412_ ), .A2(_08459_ ), .A3(\RFU.rf[12][28] ), .ZN(_08523_ ) );
AND4_X1 _16245_ ( .A1(_08520_ ), .A2(_08521_ ), .A3(_08522_ ), .A4(_08523_ ), .ZN(_08524_ ) );
NAND3_X1 _16246_ ( .A1(_08462_ ), .A2(\RFU.rf[13][28] ), .A3(_08463_ ), .ZN(_08525_ ) );
NAND3_X1 _16247_ ( .A1(_08438_ ), .A2(\RFU.rf[10][28] ), .A3(_08316_ ), .ZN(_08526_ ) );
NAND3_X1 _16248_ ( .A1(_08417_ ), .A2(\RFU.rf[8][28] ), .A3(_08418_ ), .ZN(_08527_ ) );
NAND3_X1 _16249_ ( .A1(_08366_ ), .A2(\RFU.rf[11][28] ), .A3(_08441_ ), .ZN(_08528_ ) );
AND4_X1 _16250_ ( .A1(_08525_ ), .A2(_08526_ ), .A3(_08527_ ), .A4(_08528_ ), .ZN(_08529_ ) );
NAND3_X1 _16251_ ( .A1(_08519_ ), .A2(_08524_ ), .A3(_08529_ ), .ZN(_08530_ ) );
MUX2_X1 _16252_ ( .A(\EXU.r1_i [28] ), .B(_08530_ ), .S(_08510_ ), .Z(_00694_ ) );
NAND3_X1 _16253_ ( .A1(_08370_ ), .A2(\RFU.rf[14][1] ), .A3(_08371_ ), .ZN(_08531_ ) );
NAND3_X1 _16254_ ( .A1(_08397_ ), .A2(\RFU.rf[4][1] ), .A3(_08373_ ), .ZN(_08532_ ) );
NAND3_X1 _16255_ ( .A1(_08375_ ), .A2(\RFU.rf[7][1] ), .A3(_08399_ ), .ZN(_08533_ ) );
NAND3_X1 _16256_ ( .A1(_08346_ ), .A2(_08377_ ), .A3(\RFU.rf[15][1] ), .ZN(_08534_ ) );
NAND4_X1 _16257_ ( .A1(_08531_ ), .A2(_08532_ ), .A3(_08533_ ), .A4(_08534_ ), .ZN(_08535_ ) );
AND3_X1 _16258_ ( .A1(_08349_ ), .A2(\RFU.rf[2][1] ), .A3(_08380_ ), .ZN(_08536_ ) );
AND3_X1 _16259_ ( .A1(_08351_ ), .A2(_08328_ ), .A3(\RFU.rf[6][1] ), .ZN(_08537_ ) );
AND3_X1 _16260_ ( .A1(_08353_ ), .A2(\RFU.rf[3][1] ), .A3(_08354_ ), .ZN(_08538_ ) );
NOR4_X1 _16261_ ( .A1(_08535_ ), .A2(_08536_ ), .A3(_08537_ ), .A4(_08538_ ), .ZN(_08539_ ) );
NAND3_X1 _16262_ ( .A1(_08454_ ), .A2(_08407_ ), .A3(\RFU.rf[5][1] ), .ZN(_08540_ ) );
NAND3_X1 _16263_ ( .A1(_08358_ ), .A2(_08456_ ), .A3(\RFU.rf[9][1] ), .ZN(_08541_ ) );
NAND3_X1 _16264_ ( .A1(_07991_ ), .A2(\RFU.rf[1][1] ), .A3(_08410_ ), .ZN(_08542_ ) );
NAND3_X1 _16265_ ( .A1(_08412_ ), .A2(_08459_ ), .A3(\RFU.rf[12][1] ), .ZN(_08543_ ) );
AND4_X1 _16266_ ( .A1(_08540_ ), .A2(_08541_ ), .A3(_08542_ ), .A4(_08543_ ), .ZN(_08544_ ) );
NAND3_X1 _16267_ ( .A1(_08462_ ), .A2(\RFU.rf[13][1] ), .A3(_08463_ ), .ZN(_08545_ ) );
NAND3_X1 _16268_ ( .A1(_08438_ ), .A2(\RFU.rf[10][1] ), .A3(_07978_ ), .ZN(_08546_ ) );
NAND3_X1 _16269_ ( .A1(_08417_ ), .A2(\RFU.rf[8][1] ), .A3(_08418_ ), .ZN(_08547_ ) );
NAND3_X1 _16270_ ( .A1(_08366_ ), .A2(\RFU.rf[11][1] ), .A3(_08441_ ), .ZN(_08548_ ) );
AND4_X1 _16271_ ( .A1(_08545_ ), .A2(_08546_ ), .A3(_08547_ ), .A4(_08548_ ), .ZN(_08549_ ) );
NAND3_X1 _16272_ ( .A1(_08539_ ), .A2(_08544_ ), .A3(_08549_ ), .ZN(_08550_ ) );
MUX2_X1 _16273_ ( .A(\EXU.r1_i [1] ), .B(_08550_ ), .S(_08510_ ), .Z(_00695_ ) );
NAND3_X1 _16274_ ( .A1(_08370_ ), .A2(\RFU.rf[14][0] ), .A3(_08371_ ), .ZN(_08551_ ) );
NAND3_X1 _16275_ ( .A1(_08397_ ), .A2(\RFU.rf[4][0] ), .A3(_08373_ ), .ZN(_08552_ ) );
NAND3_X1 _16276_ ( .A1(_08375_ ), .A2(\RFU.rf[7][0] ), .A3(_08399_ ), .ZN(_08553_ ) );
NAND3_X1 _16277_ ( .A1(_08346_ ), .A2(_08377_ ), .A3(\RFU.rf[15][0] ), .ZN(_08554_ ) );
NAND4_X1 _16278_ ( .A1(_08551_ ), .A2(_08552_ ), .A3(_08553_ ), .A4(_08554_ ), .ZN(_08555_ ) );
AND3_X1 _16279_ ( .A1(_08349_ ), .A2(\RFU.rf[2][0] ), .A3(_08380_ ), .ZN(_08556_ ) );
AND3_X1 _16280_ ( .A1(_08351_ ), .A2(_07995_ ), .A3(\RFU.rf[6][0] ), .ZN(_08557_ ) );
AND3_X1 _16281_ ( .A1(_08353_ ), .A2(\RFU.rf[3][0] ), .A3(_08354_ ), .ZN(_08558_ ) );
NOR4_X1 _16282_ ( .A1(_08555_ ), .A2(_08556_ ), .A3(_08557_ ), .A4(_08558_ ), .ZN(_08559_ ) );
NAND3_X1 _16283_ ( .A1(_08454_ ), .A2(_08407_ ), .A3(\RFU.rf[5][0] ), .ZN(_08560_ ) );
NAND3_X1 _16284_ ( .A1(_08358_ ), .A2(_08456_ ), .A3(\RFU.rf[9][0] ), .ZN(_08561_ ) );
NAND3_X1 _16285_ ( .A1(_07991_ ), .A2(\RFU.rf[1][0] ), .A3(_08410_ ), .ZN(_08562_ ) );
NAND3_X1 _16286_ ( .A1(_08412_ ), .A2(_08459_ ), .A3(\RFU.rf[12][0] ), .ZN(_08563_ ) );
AND4_X1 _16287_ ( .A1(_08560_ ), .A2(_08561_ ), .A3(_08562_ ), .A4(_08563_ ), .ZN(_08564_ ) );
NAND3_X1 _16288_ ( .A1(_08462_ ), .A2(\RFU.rf[13][0] ), .A3(_08463_ ), .ZN(_08565_ ) );
NAND3_X1 _16289_ ( .A1(_08438_ ), .A2(\RFU.rf[10][0] ), .A3(_07978_ ), .ZN(_08566_ ) );
NAND3_X1 _16290_ ( .A1(_08417_ ), .A2(\RFU.rf[8][0] ), .A3(_08418_ ), .ZN(_08567_ ) );
NAND3_X1 _16291_ ( .A1(_08366_ ), .A2(\RFU.rf[11][0] ), .A3(_08441_ ), .ZN(_08568_ ) );
AND4_X1 _16292_ ( .A1(_08565_ ), .A2(_08566_ ), .A3(_08567_ ), .A4(_08568_ ), .ZN(_08569_ ) );
NAND3_X1 _16293_ ( .A1(_08559_ ), .A2(_08564_ ), .A3(_08569_ ), .ZN(_08570_ ) );
MUX2_X1 _16294_ ( .A(\EXU.r1_i [0] ), .B(_08570_ ), .S(_08510_ ), .Z(_00696_ ) );
NAND3_X1 _16295_ ( .A1(_08370_ ), .A2(\RFU.rf[14][27] ), .A3(_08371_ ), .ZN(_08571_ ) );
NAND3_X1 _16296_ ( .A1(_08397_ ), .A2(\RFU.rf[4][27] ), .A3(_08373_ ), .ZN(_08572_ ) );
NAND3_X1 _16297_ ( .A1(_08375_ ), .A2(\RFU.rf[7][27] ), .A3(_08399_ ), .ZN(_08573_ ) );
NAND3_X1 _16298_ ( .A1(_07985_ ), .A2(_08377_ ), .A3(\RFU.rf[15][27] ), .ZN(_08574_ ) );
NAND4_X1 _16299_ ( .A1(_08571_ ), .A2(_08572_ ), .A3(_08573_ ), .A4(_08574_ ), .ZN(_08575_ ) );
AND3_X1 _16300_ ( .A1(_07964_ ), .A2(\RFU.rf[2][27] ), .A3(_08380_ ), .ZN(_08576_ ) );
AND3_X1 _16301_ ( .A1(_07970_ ), .A2(_07995_ ), .A3(\RFU.rf[6][27] ), .ZN(_08577_ ) );
AND3_X1 _16302_ ( .A1(_07951_ ), .A2(\RFU.rf[3][27] ), .A3(_07982_ ), .ZN(_08578_ ) );
NOR4_X1 _16303_ ( .A1(_08575_ ), .A2(_08576_ ), .A3(_08577_ ), .A4(_08578_ ), .ZN(_08579_ ) );
NAND3_X1 _16304_ ( .A1(_08454_ ), .A2(_08407_ ), .A3(\RFU.rf[5][27] ), .ZN(_08580_ ) );
NAND3_X1 _16305_ ( .A1(_07981_ ), .A2(_08456_ ), .A3(\RFU.rf[9][27] ), .ZN(_08581_ ) );
NAND3_X1 _16306_ ( .A1(_07991_ ), .A2(\RFU.rf[1][27] ), .A3(_08410_ ), .ZN(_08582_ ) );
NAND3_X1 _16307_ ( .A1(_08412_ ), .A2(_08459_ ), .A3(\RFU.rf[12][27] ), .ZN(_08583_ ) );
AND4_X1 _16308_ ( .A1(_08580_ ), .A2(_08581_ ), .A3(_08582_ ), .A4(_08583_ ), .ZN(_08584_ ) );
NAND3_X1 _16309_ ( .A1(_08462_ ), .A2(\RFU.rf[13][27] ), .A3(_08463_ ), .ZN(_08585_ ) );
NAND3_X1 _16310_ ( .A1(_08438_ ), .A2(\RFU.rf[10][27] ), .A3(_07978_ ), .ZN(_08586_ ) );
NAND3_X1 _16311_ ( .A1(_08417_ ), .A2(\RFU.rf[8][27] ), .A3(_08418_ ), .ZN(_08587_ ) );
NAND3_X1 _16312_ ( .A1(_07998_ ), .A2(\RFU.rf[11][27] ), .A3(_08441_ ), .ZN(_08588_ ) );
AND4_X1 _16313_ ( .A1(_08585_ ), .A2(_08586_ ), .A3(_08587_ ), .A4(_08588_ ), .ZN(_08589_ ) );
NAND3_X1 _16314_ ( .A1(_08579_ ), .A2(_08584_ ), .A3(_08589_ ), .ZN(_08590_ ) );
MUX2_X1 _16315_ ( .A(\EXU.r1_i [27] ), .B(_08590_ ), .S(_08510_ ), .Z(_00697_ ) );
NAND3_X1 _16316_ ( .A1(_07959_ ), .A2(\RFU.rf[14][26] ), .A3(_07954_ ), .ZN(_08591_ ) );
NAND3_X1 _16317_ ( .A1(_08397_ ), .A2(\RFU.rf[4][26] ), .A3(_07987_ ), .ZN(_08592_ ) );
NAND3_X1 _16318_ ( .A1(_07963_ ), .A2(\RFU.rf[7][26] ), .A3(_08399_ ), .ZN(_08593_ ) );
NAND3_X1 _16319_ ( .A1(_07985_ ), .A2(_07966_ ), .A3(\RFU.rf[15][26] ), .ZN(_08594_ ) );
NAND4_X1 _16320_ ( .A1(_08591_ ), .A2(_08592_ ), .A3(_08593_ ), .A4(_08594_ ), .ZN(_08595_ ) );
AND3_X1 _16321_ ( .A1(_07964_ ), .A2(\RFU.rf[2][26] ), .A3(_07967_ ), .ZN(_08596_ ) );
AND3_X1 _16322_ ( .A1(_07970_ ), .A2(_07995_ ), .A3(\RFU.rf[6][26] ), .ZN(_08597_ ) );
AND3_X1 _16323_ ( .A1(_07951_ ), .A2(\RFU.rf[3][26] ), .A3(_07982_ ), .ZN(_08598_ ) );
NOR4_X1 _16324_ ( .A1(_08595_ ), .A2(_08596_ ), .A3(_08597_ ), .A4(_08598_ ), .ZN(_08599_ ) );
NAND3_X1 _16325_ ( .A1(_08454_ ), .A2(_08407_ ), .A3(\RFU.rf[5][26] ), .ZN(_08600_ ) );
NAND3_X1 _16326_ ( .A1(_07981_ ), .A2(_08456_ ), .A3(\RFU.rf[9][26] ), .ZN(_08601_ ) );
NAND3_X1 _16327_ ( .A1(_07991_ ), .A2(\RFU.rf[1][26] ), .A3(_08410_ ), .ZN(_08602_ ) );
NAND3_X1 _16328_ ( .A1(_08412_ ), .A2(_08459_ ), .A3(\RFU.rf[12][26] ), .ZN(_08603_ ) );
AND4_X1 _16329_ ( .A1(_08600_ ), .A2(_08601_ ), .A3(_08602_ ), .A4(_08603_ ), .ZN(_08604_ ) );
NAND3_X1 _16330_ ( .A1(_08462_ ), .A2(\RFU.rf[13][26] ), .A3(_08463_ ), .ZN(_08605_ ) );
NAND3_X1 _16331_ ( .A1(_08438_ ), .A2(\RFU.rf[10][26] ), .A3(_07978_ ), .ZN(_08606_ ) );
NAND3_X1 _16332_ ( .A1(_08417_ ), .A2(\RFU.rf[8][26] ), .A3(_08418_ ), .ZN(_08607_ ) );
NAND3_X1 _16333_ ( .A1(_07998_ ), .A2(\RFU.rf[11][26] ), .A3(_08441_ ), .ZN(_08608_ ) );
AND4_X1 _16334_ ( .A1(_08605_ ), .A2(_08606_ ), .A3(_08607_ ), .A4(_08608_ ), .ZN(_08609_ ) );
NAND3_X1 _16335_ ( .A1(_08599_ ), .A2(_08604_ ), .A3(_08609_ ), .ZN(_08610_ ) );
MUX2_X1 _16336_ ( .A(\EXU.r1_i [26] ), .B(_08610_ ), .S(_08510_ ), .Z(_00698_ ) );
NAND3_X1 _16337_ ( .A1(_07959_ ), .A2(\RFU.rf[14][25] ), .A3(_07954_ ), .ZN(_08611_ ) );
NAND3_X1 _16338_ ( .A1(_07949_ ), .A2(\RFU.rf[4][25] ), .A3(_07987_ ), .ZN(_08612_ ) );
NAND3_X1 _16339_ ( .A1(_07963_ ), .A2(\RFU.rf[7][25] ), .A3(_07956_ ), .ZN(_08613_ ) );
NAND3_X1 _16340_ ( .A1(_07985_ ), .A2(_07966_ ), .A3(\RFU.rf[15][25] ), .ZN(_08614_ ) );
NAND4_X1 _16341_ ( .A1(_08611_ ), .A2(_08612_ ), .A3(_08613_ ), .A4(_08614_ ), .ZN(_08615_ ) );
AND3_X1 _16342_ ( .A1(_07964_ ), .A2(\RFU.rf[2][25] ), .A3(_07967_ ), .ZN(_08616_ ) );
AND3_X1 _16343_ ( .A1(_07970_ ), .A2(_07995_ ), .A3(\RFU.rf[6][25] ), .ZN(_08617_ ) );
AND3_X1 _16344_ ( .A1(_07951_ ), .A2(\RFU.rf[3][25] ), .A3(_07982_ ), .ZN(_08618_ ) );
NOR4_X1 _16345_ ( .A1(_08615_ ), .A2(_08616_ ), .A3(_08617_ ), .A4(_08618_ ), .ZN(_08619_ ) );
NAND3_X1 _16346_ ( .A1(_08454_ ), .A2(_07976_ ), .A3(\RFU.rf[5][25] ), .ZN(_08620_ ) );
NAND3_X1 _16347_ ( .A1(_07981_ ), .A2(_08456_ ), .A3(\RFU.rf[9][25] ), .ZN(_08621_ ) );
NAND3_X1 _16348_ ( .A1(_07991_ ), .A2(\RFU.rf[1][25] ), .A3(_07961_ ), .ZN(_08622_ ) );
NAND3_X1 _16349_ ( .A1(_07940_ ), .A2(_08459_ ), .A3(\RFU.rf[12][25] ), .ZN(_08623_ ) );
AND4_X1 _16350_ ( .A1(_08620_ ), .A2(_08621_ ), .A3(_08622_ ), .A4(_08623_ ), .ZN(_08624_ ) );
NAND3_X1 _16351_ ( .A1(_08462_ ), .A2(\RFU.rf[13][25] ), .A3(_08463_ ), .ZN(_08625_ ) );
NAND3_X1 _16352_ ( .A1(_08438_ ), .A2(\RFU.rf[10][25] ), .A3(_07978_ ), .ZN(_08626_ ) );
NAND3_X1 _16353_ ( .A1(_08003_ ), .A2(\RFU.rf[8][25] ), .A3(_07947_ ), .ZN(_08627_ ) );
NAND3_X1 _16354_ ( .A1(_07998_ ), .A2(\RFU.rf[11][25] ), .A3(_08441_ ), .ZN(_08628_ ) );
AND4_X1 _16355_ ( .A1(_08625_ ), .A2(_08626_ ), .A3(_08627_ ), .A4(_08628_ ), .ZN(_08629_ ) );
NAND3_X1 _16356_ ( .A1(_08619_ ), .A2(_08624_ ), .A3(_08629_ ), .ZN(_08630_ ) );
MUX2_X1 _16357_ ( .A(\EXU.r1_i [25] ), .B(_08630_ ), .S(_08510_ ), .Z(_00699_ ) );
NAND3_X1 _16358_ ( .A1(_07959_ ), .A2(\RFU.rf[14][24] ), .A3(_07954_ ), .ZN(_08631_ ) );
NAND3_X1 _16359_ ( .A1(_07949_ ), .A2(\RFU.rf[4][24] ), .A3(_07987_ ), .ZN(_08632_ ) );
NAND3_X1 _16360_ ( .A1(_07963_ ), .A2(\RFU.rf[7][24] ), .A3(_07956_ ), .ZN(_08633_ ) );
NAND3_X1 _16361_ ( .A1(_07985_ ), .A2(_07966_ ), .A3(\RFU.rf[15][24] ), .ZN(_08634_ ) );
NAND4_X1 _16362_ ( .A1(_08631_ ), .A2(_08632_ ), .A3(_08633_ ), .A4(_08634_ ), .ZN(_08635_ ) );
AND3_X1 _16363_ ( .A1(_07964_ ), .A2(\RFU.rf[2][24] ), .A3(_07967_ ), .ZN(_08636_ ) );
AND3_X1 _16364_ ( .A1(_07970_ ), .A2(_07995_ ), .A3(\RFU.rf[6][24] ), .ZN(_08637_ ) );
AND3_X1 _16365_ ( .A1(_07951_ ), .A2(\RFU.rf[3][24] ), .A3(_07982_ ), .ZN(_08638_ ) );
NOR4_X1 _16366_ ( .A1(_08635_ ), .A2(_08636_ ), .A3(_08637_ ), .A4(_08638_ ), .ZN(_08639_ ) );
NAND3_X1 _16367_ ( .A1(_08454_ ), .A2(_07976_ ), .A3(\RFU.rf[5][24] ), .ZN(_08640_ ) );
NAND3_X1 _16368_ ( .A1(_07981_ ), .A2(_08456_ ), .A3(\RFU.rf[9][24] ), .ZN(_08641_ ) );
NAND3_X1 _16369_ ( .A1(_07991_ ), .A2(\RFU.rf[1][24] ), .A3(_07961_ ), .ZN(_08642_ ) );
NAND3_X1 _16370_ ( .A1(_07940_ ), .A2(_08459_ ), .A3(\RFU.rf[12][24] ), .ZN(_08643_ ) );
AND4_X1 _16371_ ( .A1(_08640_ ), .A2(_08641_ ), .A3(_08642_ ), .A4(_08643_ ), .ZN(_08644_ ) );
NAND3_X1 _16372_ ( .A1(_08462_ ), .A2(\RFU.rf[13][24] ), .A3(_08463_ ), .ZN(_08645_ ) );
NAND3_X1 _16373_ ( .A1(_07937_ ), .A2(\RFU.rf[10][24] ), .A3(_07978_ ), .ZN(_08646_ ) );
NAND3_X1 _16374_ ( .A1(_08003_ ), .A2(\RFU.rf[8][24] ), .A3(_07947_ ), .ZN(_08647_ ) );
NAND3_X1 _16375_ ( .A1(_07998_ ), .A2(\RFU.rf[11][24] ), .A3(_07952_ ), .ZN(_08648_ ) );
AND4_X1 _16376_ ( .A1(_08645_ ), .A2(_08646_ ), .A3(_08647_ ), .A4(_08648_ ), .ZN(_08649_ ) );
NAND3_X1 _16377_ ( .A1(_08639_ ), .A2(_08644_ ), .A3(_08649_ ), .ZN(_08650_ ) );
MUX2_X1 _16378_ ( .A(\EXU.r1_i [24] ), .B(_08650_ ), .S(_08510_ ), .Z(_00700_ ) );
NAND3_X1 _16379_ ( .A1(_07959_ ), .A2(\RFU.rf[14][23] ), .A3(_07954_ ), .ZN(_08651_ ) );
NAND3_X1 _16380_ ( .A1(_07949_ ), .A2(\RFU.rf[4][23] ), .A3(_07987_ ), .ZN(_08652_ ) );
NAND3_X1 _16381_ ( .A1(_07963_ ), .A2(\RFU.rf[7][23] ), .A3(_07956_ ), .ZN(_08653_ ) );
NAND3_X1 _16382_ ( .A1(_07985_ ), .A2(_07966_ ), .A3(\RFU.rf[15][23] ), .ZN(_08654_ ) );
NAND4_X1 _16383_ ( .A1(_08651_ ), .A2(_08652_ ), .A3(_08653_ ), .A4(_08654_ ), .ZN(_08655_ ) );
AND3_X1 _16384_ ( .A1(_07964_ ), .A2(\RFU.rf[2][23] ), .A3(_07967_ ), .ZN(_08656_ ) );
AND3_X1 _16385_ ( .A1(_07970_ ), .A2(_07995_ ), .A3(\RFU.rf[6][23] ), .ZN(_08657_ ) );
AND3_X1 _16386_ ( .A1(_07951_ ), .A2(\RFU.rf[3][23] ), .A3(_07982_ ), .ZN(_08658_ ) );
NOR4_X1 _16387_ ( .A1(_08655_ ), .A2(_08656_ ), .A3(_08657_ ), .A4(_08658_ ), .ZN(_08659_ ) );
NAND3_X1 _16388_ ( .A1(_07945_ ), .A2(_07976_ ), .A3(\RFU.rf[5][23] ), .ZN(_08660_ ) );
NAND3_X1 _16389_ ( .A1(_07981_ ), .A2(_08000_ ), .A3(\RFU.rf[9][23] ), .ZN(_08661_ ) );
NAND3_X1 _16390_ ( .A1(_07991_ ), .A2(\RFU.rf[1][23] ), .A3(_07961_ ), .ZN(_08662_ ) );
NAND3_X1 _16391_ ( .A1(_07940_ ), .A2(_08001_ ), .A3(\RFU.rf[12][23] ), .ZN(_08663_ ) );
AND4_X1 _16392_ ( .A1(_08660_ ), .A2(_08661_ ), .A3(_08662_ ), .A4(_08663_ ), .ZN(_08664_ ) );
NAND3_X1 _16393_ ( .A1(_07974_ ), .A2(\RFU.rf[13][23] ), .A3(_07986_ ), .ZN(_08665_ ) );
NAND3_X1 _16394_ ( .A1(_07937_ ), .A2(\RFU.rf[10][23] ), .A3(_07978_ ), .ZN(_08666_ ) );
NAND3_X1 _16395_ ( .A1(_08003_ ), .A2(\RFU.rf[8][23] ), .A3(_07947_ ), .ZN(_08667_ ) );
NAND3_X1 _16396_ ( .A1(_07998_ ), .A2(\RFU.rf[11][23] ), .A3(_07952_ ), .ZN(_08668_ ) );
AND4_X1 _16397_ ( .A1(_08665_ ), .A2(_08666_ ), .A3(_08667_ ), .A4(_08668_ ), .ZN(_08669_ ) );
NAND3_X1 _16398_ ( .A1(_08659_ ), .A2(_08664_ ), .A3(_08669_ ), .ZN(_08670_ ) );
MUX2_X1 _16399_ ( .A(\EXU.r1_i [23] ), .B(_08670_ ), .S(_08510_ ), .Z(_00701_ ) );
NAND3_X1 _16400_ ( .A1(_07959_ ), .A2(\RFU.rf[14][22] ), .A3(_07954_ ), .ZN(_08671_ ) );
NAND3_X1 _16401_ ( .A1(_07949_ ), .A2(\RFU.rf[4][22] ), .A3(_07987_ ), .ZN(_08672_ ) );
NAND3_X1 _16402_ ( .A1(_07963_ ), .A2(\RFU.rf[7][22] ), .A3(_07956_ ), .ZN(_08673_ ) );
NAND3_X1 _16403_ ( .A1(_07985_ ), .A2(_07966_ ), .A3(\RFU.rf[15][22] ), .ZN(_08674_ ) );
NAND4_X1 _16404_ ( .A1(_08671_ ), .A2(_08672_ ), .A3(_08673_ ), .A4(_08674_ ), .ZN(_08675_ ) );
AND3_X1 _16405_ ( .A1(_07964_ ), .A2(\RFU.rf[2][22] ), .A3(_07967_ ), .ZN(_08676_ ) );
AND3_X1 _16406_ ( .A1(_07970_ ), .A2(_07995_ ), .A3(\RFU.rf[6][22] ), .ZN(_08677_ ) );
AND3_X1 _16407_ ( .A1(_07951_ ), .A2(\RFU.rf[3][22] ), .A3(_07982_ ), .ZN(_08678_ ) );
NOR4_X1 _16408_ ( .A1(_08675_ ), .A2(_08676_ ), .A3(_08677_ ), .A4(_08678_ ), .ZN(_08679_ ) );
NAND3_X1 _16409_ ( .A1(_07945_ ), .A2(_07976_ ), .A3(\RFU.rf[5][22] ), .ZN(_08680_ ) );
NAND3_X1 _16410_ ( .A1(_07981_ ), .A2(_08000_ ), .A3(\RFU.rf[9][22] ), .ZN(_08681_ ) );
NAND3_X1 _16411_ ( .A1(_07991_ ), .A2(\RFU.rf[1][22] ), .A3(_07961_ ), .ZN(_08682_ ) );
NAND3_X1 _16412_ ( .A1(_07940_ ), .A2(_08001_ ), .A3(\RFU.rf[12][22] ), .ZN(_08683_ ) );
AND4_X1 _16413_ ( .A1(_08680_ ), .A2(_08681_ ), .A3(_08682_ ), .A4(_08683_ ), .ZN(_08684_ ) );
NAND3_X1 _16414_ ( .A1(_07974_ ), .A2(\RFU.rf[13][22] ), .A3(_07986_ ), .ZN(_08685_ ) );
NAND3_X1 _16415_ ( .A1(_07937_ ), .A2(\RFU.rf[10][22] ), .A3(_07978_ ), .ZN(_08686_ ) );
NAND3_X1 _16416_ ( .A1(_08003_ ), .A2(\RFU.rf[8][22] ), .A3(_07947_ ), .ZN(_08687_ ) );
NAND3_X1 _16417_ ( .A1(_07998_ ), .A2(\RFU.rf[11][22] ), .A3(_07952_ ), .ZN(_08688_ ) );
AND4_X1 _16418_ ( .A1(_08685_ ), .A2(_08686_ ), .A3(_08687_ ), .A4(_08688_ ), .ZN(_08689_ ) );
NAND3_X1 _16419_ ( .A1(_08679_ ), .A2(_08684_ ), .A3(_08689_ ), .ZN(_08690_ ) );
MUX2_X1 _16420_ ( .A(\EXU.r1_i [22] ), .B(_08690_ ), .S(_08510_ ), .Z(_00702_ ) );
INV_X1 _16421_ ( .A(_05485_ ), .ZN(_08691_ ) );
NOR2_X1 _16422_ ( .A1(_08691_ ), .A2(_05491_ ), .ZN(_08692_ ) );
BUF_X4 _16423_ ( .A(_08692_ ), .Z(_08693_ ) );
BUF_X4 _16424_ ( .A(_08693_ ), .Z(_08694_ ) );
AND2_X2 _16425_ ( .A1(_05488_ ), .A2(_05494_ ), .ZN(_08695_ ) );
BUF_X4 _16426_ ( .A(_08695_ ), .Z(_08696_ ) );
BUF_X4 _16427_ ( .A(_08696_ ), .Z(_08697_ ) );
NAND3_X1 _16428_ ( .A1(_08694_ ), .A2(\RFU.rf[11][31] ), .A3(_08697_ ), .ZN(_08698_ ) );
AND2_X2 _16429_ ( .A1(_08691_ ), .A2(_05491_ ), .ZN(_08699_ ) );
BUF_X4 _16430_ ( .A(_08699_ ), .Z(_08700_ ) );
BUF_X4 _16431_ ( .A(_08700_ ), .Z(_08701_ ) );
BUF_X8 _16432_ ( .A(_08695_ ), .Z(_08702_ ) );
BUF_X4 _16433_ ( .A(_08702_ ), .Z(_08703_ ) );
NAND3_X1 _16434_ ( .A1(_08701_ ), .A2(\RFU.rf[7][31] ), .A3(_08703_ ), .ZN(_08704_ ) );
BUF_X8 _16435_ ( .A(_08699_ ), .Z(_08705_ ) );
BUF_X4 _16436_ ( .A(_08705_ ), .Z(_08706_ ) );
INV_X1 _16437_ ( .A(_05488_ ), .ZN(_08707_ ) );
NOR2_X1 _16438_ ( .A1(_08707_ ), .A2(_05494_ ), .ZN(_08708_ ) );
BUF_X8 _16439_ ( .A(_08708_ ), .Z(_08709_ ) );
BUF_X4 _16440_ ( .A(_08709_ ), .Z(_08710_ ) );
NAND3_X1 _16441_ ( .A1(_08706_ ), .A2(\RFU.rf[5][31] ), .A3(_08710_ ), .ZN(_08711_ ) );
AND2_X2 _16442_ ( .A1(_08707_ ), .A2(_05494_ ), .ZN(_08712_ ) );
BUF_X8 _16443_ ( .A(_08712_ ), .Z(_08713_ ) );
BUF_X4 _16444_ ( .A(_08713_ ), .Z(_08714_ ) );
BUF_X8 _16445_ ( .A(_08692_ ), .Z(_08715_ ) );
BUF_X4 _16446_ ( .A(_08715_ ), .Z(_08716_ ) );
NAND3_X1 _16447_ ( .A1(_08714_ ), .A2(_08716_ ), .A3(\RFU.rf[10][31] ), .ZN(_08717_ ) );
AND4_X1 _16448_ ( .A1(_08698_ ), .A2(_08704_ ), .A3(_08711_ ), .A4(_08717_ ), .ZN(_08718_ ) );
AND2_X2 _16449_ ( .A1(_05485_ ), .A2(_05491_ ), .ZN(_08719_ ) );
BUF_X4 _16450_ ( .A(_08719_ ), .Z(_08720_ ) );
BUF_X4 _16451_ ( .A(_08720_ ), .Z(_08721_ ) );
OAI21_X2 _16452_ ( .A(_05483_ ), .B1(_05487_ ), .B2(_05493_ ), .ZN(_08722_ ) );
BUF_X4 _16453_ ( .A(_08722_ ), .Z(_08723_ ) );
BUF_X4 _16454_ ( .A(_08723_ ), .Z(_08724_ ) );
NAND3_X1 _16455_ ( .A1(_08721_ ), .A2(\RFU.rf[12][31] ), .A3(_08724_ ), .ZN(_08725_ ) );
BUF_X4 _16456_ ( .A(_08713_ ), .Z(_08726_ ) );
BUF_X4 _16457_ ( .A(_08705_ ), .Z(_08727_ ) );
NAND3_X1 _16458_ ( .A1(_08726_ ), .A2(_08727_ ), .A3(\RFU.rf[6][31] ), .ZN(_08728_ ) );
BUF_X8 _16459_ ( .A(_08719_ ), .Z(_08729_ ) );
BUF_X4 _16460_ ( .A(_08729_ ), .Z(_08730_ ) );
BUF_X4 _16461_ ( .A(_08702_ ), .Z(_08731_ ) );
NAND3_X1 _16462_ ( .A1(_08730_ ), .A2(_08731_ ), .A3(\RFU.rf[15][31] ), .ZN(_08732_ ) );
BUF_X4 _16463_ ( .A(_08715_ ), .Z(_08733_ ) );
BUF_X4 _16464_ ( .A(_08722_ ), .Z(_08734_ ) );
NAND3_X1 _16465_ ( .A1(_08733_ ), .A2(\RFU.rf[8][31] ), .A3(_08734_ ), .ZN(_08735_ ) );
AND4_X1 _16466_ ( .A1(_08725_ ), .A2(_08728_ ), .A3(_08732_ ), .A4(_08735_ ), .ZN(_08736_ ) );
BUF_X4 _16467_ ( .A(_08712_ ), .Z(_08737_ ) );
BUF_X4 _16468_ ( .A(_08737_ ), .Z(_08738_ ) );
BUF_X4 _16469_ ( .A(_08729_ ), .Z(_08739_ ) );
NAND3_X1 _16470_ ( .A1(_08738_ ), .A2(\RFU.rf[14][31] ), .A3(_08739_ ), .ZN(_08740_ ) );
BUF_X4 _16471_ ( .A(_08705_ ), .Z(_08741_ ) );
BUF_X4 _16472_ ( .A(_08723_ ), .Z(_08742_ ) );
NAND3_X1 _16473_ ( .A1(_08741_ ), .A2(\RFU.rf[4][31] ), .A3(_08742_ ), .ZN(_08743_ ) );
BUF_X4 _16474_ ( .A(_08713_ ), .Z(_08744_ ) );
OAI21_X2 _16475_ ( .A(_05483_ ), .B1(_05484_ ), .B2(_05490_ ), .ZN(_08745_ ) );
BUF_X4 _16476_ ( .A(_08745_ ), .Z(_08746_ ) );
NAND3_X1 _16477_ ( .A1(_08744_ ), .A2(\RFU.rf[2][31] ), .A3(_08746_ ), .ZN(_08747_ ) );
BUF_X4 _16478_ ( .A(_08709_ ), .Z(_08748_ ) );
BUF_X4 _16479_ ( .A(_08729_ ), .Z(_08749_ ) );
NAND3_X1 _16480_ ( .A1(_08748_ ), .A2(\RFU.rf[13][31] ), .A3(_08749_ ), .ZN(_08750_ ) );
AND4_X1 _16481_ ( .A1(_08740_ ), .A2(_08743_ ), .A3(_08747_ ), .A4(_08750_ ), .ZN(_08751_ ) );
BUF_X4 _16482_ ( .A(_08708_ ), .Z(_08752_ ) );
BUF_X4 _16483_ ( .A(_08752_ ), .Z(_08753_ ) );
BUF_X4 _16484_ ( .A(_08715_ ), .Z(_08754_ ) );
NAND3_X1 _16485_ ( .A1(_08753_ ), .A2(_08754_ ), .A3(\RFU.rf[9][31] ), .ZN(_08755_ ) );
BUF_X4 _16486_ ( .A(_08709_ ), .Z(_08756_ ) );
BUF_X4 _16487_ ( .A(_08745_ ), .Z(_08757_ ) );
BUF_X4 _16488_ ( .A(_08757_ ), .Z(_08758_ ) );
NAND3_X1 _16489_ ( .A1(_08756_ ), .A2(\RFU.rf[1][31] ), .A3(_08758_ ), .ZN(_08759_ ) );
BUF_X4 _16490_ ( .A(_08702_ ), .Z(_08760_ ) );
BUF_X4 _16491_ ( .A(_08757_ ), .Z(_08761_ ) );
NAND3_X1 _16492_ ( .A1(_08760_ ), .A2(\RFU.rf[3][31] ), .A3(_08761_ ), .ZN(_08762_ ) );
AND3_X1 _16493_ ( .A1(_08755_ ), .A2(_08759_ ), .A3(_08762_ ), .ZN(_08763_ ) );
NAND4_X1 _16494_ ( .A1(_08718_ ), .A2(_08736_ ), .A3(_08751_ ), .A4(_08763_ ), .ZN(_08764_ ) );
BUF_X4 _16495_ ( .A(_05514_ ), .Z(_08765_ ) );
MUX2_X1 _16496_ ( .A(\EXU.r2_i [31] ), .B(_08764_ ), .S(_08765_ ), .Z(_00703_ ) );
NAND3_X1 _16497_ ( .A1(_08694_ ), .A2(\RFU.rf[11][30] ), .A3(_08697_ ), .ZN(_08766_ ) );
NAND3_X1 _16498_ ( .A1(_08701_ ), .A2(\RFU.rf[7][30] ), .A3(_08703_ ), .ZN(_08767_ ) );
NAND3_X1 _16499_ ( .A1(_08706_ ), .A2(\RFU.rf[5][30] ), .A3(_08710_ ), .ZN(_08768_ ) );
BUF_X4 _16500_ ( .A(_08713_ ), .Z(_08769_ ) );
NAND3_X1 _16501_ ( .A1(_08769_ ), .A2(_08716_ ), .A3(\RFU.rf[10][30] ), .ZN(_08770_ ) );
AND4_X1 _16502_ ( .A1(_08766_ ), .A2(_08767_ ), .A3(_08768_ ), .A4(_08770_ ), .ZN(_08771_ ) );
NAND3_X1 _16503_ ( .A1(_08721_ ), .A2(\RFU.rf[12][30] ), .A3(_08724_ ), .ZN(_08772_ ) );
BUF_X4 _16504_ ( .A(_08705_ ), .Z(_08773_ ) );
NAND3_X1 _16505_ ( .A1(_08726_ ), .A2(_08773_ ), .A3(\RFU.rf[6][30] ), .ZN(_08774_ ) );
NAND3_X1 _16506_ ( .A1(_08730_ ), .A2(_08731_ ), .A3(\RFU.rf[15][30] ), .ZN(_08775_ ) );
NAND3_X1 _16507_ ( .A1(_08733_ ), .A2(\RFU.rf[8][30] ), .A3(_08734_ ), .ZN(_08776_ ) );
AND4_X1 _16508_ ( .A1(_08772_ ), .A2(_08774_ ), .A3(_08775_ ), .A4(_08776_ ), .ZN(_08777_ ) );
NAND3_X1 _16509_ ( .A1(_08738_ ), .A2(\RFU.rf[14][30] ), .A3(_08739_ ), .ZN(_08778_ ) );
NAND3_X1 _16510_ ( .A1(_08741_ ), .A2(\RFU.rf[4][30] ), .A3(_08742_ ), .ZN(_08779_ ) );
BUF_X4 _16511_ ( .A(_08713_ ), .Z(_08780_ ) );
NAND3_X1 _16512_ ( .A1(_08780_ ), .A2(\RFU.rf[2][30] ), .A3(_08746_ ), .ZN(_08781_ ) );
BUF_X4 _16513_ ( .A(_08709_ ), .Z(_08782_ ) );
BUF_X4 _16514_ ( .A(_08729_ ), .Z(_08783_ ) );
NAND3_X1 _16515_ ( .A1(_08782_ ), .A2(\RFU.rf[13][30] ), .A3(_08783_ ), .ZN(_08784_ ) );
AND4_X1 _16516_ ( .A1(_08778_ ), .A2(_08779_ ), .A3(_08781_ ), .A4(_08784_ ), .ZN(_08785_ ) );
NAND3_X1 _16517_ ( .A1(_08753_ ), .A2(_08754_ ), .A3(\RFU.rf[9][30] ), .ZN(_08786_ ) );
NAND3_X1 _16518_ ( .A1(_08756_ ), .A2(\RFU.rf[1][30] ), .A3(_08758_ ), .ZN(_08787_ ) );
NAND3_X1 _16519_ ( .A1(_08760_ ), .A2(\RFU.rf[3][30] ), .A3(_08761_ ), .ZN(_08788_ ) );
AND3_X1 _16520_ ( .A1(_08786_ ), .A2(_08787_ ), .A3(_08788_ ), .ZN(_08789_ ) );
NAND4_X1 _16521_ ( .A1(_08771_ ), .A2(_08777_ ), .A3(_08785_ ), .A4(_08789_ ), .ZN(_08790_ ) );
MUX2_X1 _16522_ ( .A(\EXU.r2_i [30] ), .B(_08790_ ), .S(_08765_ ), .Z(_00704_ ) );
NAND3_X1 _16523_ ( .A1(_08694_ ), .A2(\RFU.rf[11][21] ), .A3(_08697_ ), .ZN(_08791_ ) );
NAND3_X1 _16524_ ( .A1(_08701_ ), .A2(\RFU.rf[7][21] ), .A3(_08703_ ), .ZN(_08792_ ) );
NAND3_X1 _16525_ ( .A1(_08706_ ), .A2(\RFU.rf[5][21] ), .A3(_08710_ ), .ZN(_08793_ ) );
NAND3_X1 _16526_ ( .A1(_08769_ ), .A2(_08716_ ), .A3(\RFU.rf[10][21] ), .ZN(_08794_ ) );
AND4_X1 _16527_ ( .A1(_08791_ ), .A2(_08792_ ), .A3(_08793_ ), .A4(_08794_ ), .ZN(_08795_ ) );
NAND3_X1 _16528_ ( .A1(_08721_ ), .A2(\RFU.rf[12][21] ), .A3(_08724_ ), .ZN(_08796_ ) );
BUF_X4 _16529_ ( .A(_08713_ ), .Z(_08797_ ) );
NAND3_X1 _16530_ ( .A1(_08797_ ), .A2(_08773_ ), .A3(\RFU.rf[6][21] ), .ZN(_08798_ ) );
NAND3_X1 _16531_ ( .A1(_08730_ ), .A2(_08731_ ), .A3(\RFU.rf[15][21] ), .ZN(_08799_ ) );
NAND3_X1 _16532_ ( .A1(_08733_ ), .A2(\RFU.rf[8][21] ), .A3(_08734_ ), .ZN(_08800_ ) );
AND4_X1 _16533_ ( .A1(_08796_ ), .A2(_08798_ ), .A3(_08799_ ), .A4(_08800_ ), .ZN(_08801_ ) );
NAND3_X1 _16534_ ( .A1(_08738_ ), .A2(\RFU.rf[14][21] ), .A3(_08739_ ), .ZN(_08802_ ) );
NAND3_X1 _16535_ ( .A1(_08741_ ), .A2(\RFU.rf[4][21] ), .A3(_08742_ ), .ZN(_08803_ ) );
NAND3_X1 _16536_ ( .A1(_08780_ ), .A2(\RFU.rf[2][21] ), .A3(_08746_ ), .ZN(_08804_ ) );
NAND3_X1 _16537_ ( .A1(_08782_ ), .A2(\RFU.rf[13][21] ), .A3(_08783_ ), .ZN(_08805_ ) );
AND4_X1 _16538_ ( .A1(_08802_ ), .A2(_08803_ ), .A3(_08804_ ), .A4(_08805_ ), .ZN(_08806_ ) );
NAND3_X1 _16539_ ( .A1(_08753_ ), .A2(_08754_ ), .A3(\RFU.rf[9][21] ), .ZN(_08807_ ) );
NAND3_X1 _16540_ ( .A1(_08756_ ), .A2(\RFU.rf[1][21] ), .A3(_08758_ ), .ZN(_08808_ ) );
NAND3_X1 _16541_ ( .A1(_08760_ ), .A2(\RFU.rf[3][21] ), .A3(_08761_ ), .ZN(_08809_ ) );
AND3_X1 _16542_ ( .A1(_08807_ ), .A2(_08808_ ), .A3(_08809_ ), .ZN(_08810_ ) );
NAND4_X1 _16543_ ( .A1(_08795_ ), .A2(_08801_ ), .A3(_08806_ ), .A4(_08810_ ), .ZN(_08811_ ) );
MUX2_X1 _16544_ ( .A(\EXU.r2_i [21] ), .B(_08811_ ), .S(_08765_ ), .Z(_00705_ ) );
NAND3_X1 _16545_ ( .A1(_08694_ ), .A2(\RFU.rf[11][20] ), .A3(_08697_ ), .ZN(_08812_ ) );
NAND3_X1 _16546_ ( .A1(_08701_ ), .A2(\RFU.rf[7][20] ), .A3(_08703_ ), .ZN(_08813_ ) );
BUF_X4 _16547_ ( .A(_08709_ ), .Z(_08814_ ) );
NAND3_X1 _16548_ ( .A1(_08706_ ), .A2(\RFU.rf[5][20] ), .A3(_08814_ ), .ZN(_08815_ ) );
NAND3_X1 _16549_ ( .A1(_08769_ ), .A2(_08716_ ), .A3(\RFU.rf[10][20] ), .ZN(_08816_ ) );
AND4_X1 _16550_ ( .A1(_08812_ ), .A2(_08813_ ), .A3(_08815_ ), .A4(_08816_ ), .ZN(_08817_ ) );
NAND3_X1 _16551_ ( .A1(_08721_ ), .A2(\RFU.rf[12][20] ), .A3(_08724_ ), .ZN(_08818_ ) );
NAND3_X1 _16552_ ( .A1(_08797_ ), .A2(_08773_ ), .A3(\RFU.rf[6][20] ), .ZN(_08819_ ) );
BUF_X4 _16553_ ( .A(_08702_ ), .Z(_08820_ ) );
NAND3_X1 _16554_ ( .A1(_08730_ ), .A2(_08820_ ), .A3(\RFU.rf[15][20] ), .ZN(_08821_ ) );
NAND3_X1 _16555_ ( .A1(_08733_ ), .A2(\RFU.rf[8][20] ), .A3(_08734_ ), .ZN(_08822_ ) );
AND4_X1 _16556_ ( .A1(_08818_ ), .A2(_08819_ ), .A3(_08821_ ), .A4(_08822_ ), .ZN(_08823_ ) );
BUF_X4 _16557_ ( .A(_08737_ ), .Z(_08824_ ) );
NAND3_X1 _16558_ ( .A1(_08824_ ), .A2(\RFU.rf[14][20] ), .A3(_08739_ ), .ZN(_08825_ ) );
NAND3_X1 _16559_ ( .A1(_08741_ ), .A2(\RFU.rf[4][20] ), .A3(_08742_ ), .ZN(_08826_ ) );
BUF_X4 _16560_ ( .A(_08745_ ), .Z(_08827_ ) );
NAND3_X1 _16561_ ( .A1(_08780_ ), .A2(\RFU.rf[2][20] ), .A3(_08827_ ), .ZN(_08828_ ) );
NAND3_X1 _16562_ ( .A1(_08782_ ), .A2(\RFU.rf[13][20] ), .A3(_08783_ ), .ZN(_08829_ ) );
AND4_X1 _16563_ ( .A1(_08825_ ), .A2(_08826_ ), .A3(_08828_ ), .A4(_08829_ ), .ZN(_08830_ ) );
NAND3_X1 _16564_ ( .A1(_08753_ ), .A2(_08754_ ), .A3(\RFU.rf[9][20] ), .ZN(_08831_ ) );
NAND3_X1 _16565_ ( .A1(_08756_ ), .A2(\RFU.rf[1][20] ), .A3(_08758_ ), .ZN(_08832_ ) );
NAND3_X1 _16566_ ( .A1(_08760_ ), .A2(\RFU.rf[3][20] ), .A3(_08761_ ), .ZN(_08833_ ) );
AND3_X1 _16567_ ( .A1(_08831_ ), .A2(_08832_ ), .A3(_08833_ ), .ZN(_08834_ ) );
NAND4_X1 _16568_ ( .A1(_08817_ ), .A2(_08823_ ), .A3(_08830_ ), .A4(_08834_ ), .ZN(_08835_ ) );
MUX2_X1 _16569_ ( .A(\EXU.r2_i [20] ), .B(_08835_ ), .S(_08765_ ), .Z(_00706_ ) );
NAND3_X1 _16570_ ( .A1(_08694_ ), .A2(\RFU.rf[11][19] ), .A3(_08697_ ), .ZN(_08836_ ) );
BUF_X4 _16571_ ( .A(_08700_ ), .Z(_08837_ ) );
NAND3_X1 _16572_ ( .A1(_08837_ ), .A2(\RFU.rf[7][19] ), .A3(_08703_ ), .ZN(_08838_ ) );
NAND3_X1 _16573_ ( .A1(_08706_ ), .A2(\RFU.rf[5][19] ), .A3(_08814_ ), .ZN(_08839_ ) );
NAND3_X1 _16574_ ( .A1(_08769_ ), .A2(_08716_ ), .A3(\RFU.rf[10][19] ), .ZN(_08840_ ) );
AND4_X1 _16575_ ( .A1(_08836_ ), .A2(_08838_ ), .A3(_08839_ ), .A4(_08840_ ), .ZN(_08841_ ) );
NAND3_X1 _16576_ ( .A1(_08721_ ), .A2(\RFU.rf[12][19] ), .A3(_08724_ ), .ZN(_08842_ ) );
NAND3_X1 _16577_ ( .A1(_08797_ ), .A2(_08773_ ), .A3(\RFU.rf[6][19] ), .ZN(_08843_ ) );
NAND3_X1 _16578_ ( .A1(_08730_ ), .A2(_08820_ ), .A3(\RFU.rf[15][19] ), .ZN(_08844_ ) );
NAND3_X1 _16579_ ( .A1(_08733_ ), .A2(\RFU.rf[8][19] ), .A3(_08734_ ), .ZN(_08845_ ) );
AND4_X1 _16580_ ( .A1(_08842_ ), .A2(_08843_ ), .A3(_08844_ ), .A4(_08845_ ), .ZN(_08846_ ) );
NAND3_X1 _16581_ ( .A1(_08824_ ), .A2(\RFU.rf[14][19] ), .A3(_08739_ ), .ZN(_08847_ ) );
NAND3_X1 _16582_ ( .A1(_08741_ ), .A2(\RFU.rf[4][19] ), .A3(_08742_ ), .ZN(_08848_ ) );
NAND3_X1 _16583_ ( .A1(_08780_ ), .A2(\RFU.rf[2][19] ), .A3(_08827_ ), .ZN(_08849_ ) );
NAND3_X1 _16584_ ( .A1(_08782_ ), .A2(\RFU.rf[13][19] ), .A3(_08783_ ), .ZN(_08850_ ) );
AND4_X1 _16585_ ( .A1(_08847_ ), .A2(_08848_ ), .A3(_08849_ ), .A4(_08850_ ), .ZN(_08851_ ) );
NAND3_X1 _16586_ ( .A1(_08753_ ), .A2(_08754_ ), .A3(\RFU.rf[9][19] ), .ZN(_08852_ ) );
NAND3_X1 _16587_ ( .A1(_08756_ ), .A2(\RFU.rf[1][19] ), .A3(_08758_ ), .ZN(_08853_ ) );
NAND3_X1 _16588_ ( .A1(_08760_ ), .A2(\RFU.rf[3][19] ), .A3(_08761_ ), .ZN(_08854_ ) );
AND3_X1 _16589_ ( .A1(_08852_ ), .A2(_08853_ ), .A3(_08854_ ), .ZN(_08855_ ) );
NAND4_X1 _16590_ ( .A1(_08841_ ), .A2(_08846_ ), .A3(_08851_ ), .A4(_08855_ ), .ZN(_08856_ ) );
MUX2_X1 _16591_ ( .A(\EXU.r2_i [19] ), .B(_08856_ ), .S(_08765_ ), .Z(_00707_ ) );
NAND3_X1 _16592_ ( .A1(_08701_ ), .A2(\RFU.rf[4][18] ), .A3(_08724_ ), .ZN(_08857_ ) );
BUF_X4 _16593_ ( .A(_08705_ ), .Z(_08858_ ) );
NAND3_X1 _16594_ ( .A1(_08738_ ), .A2(_08858_ ), .A3(\RFU.rf[6][18] ), .ZN(_08859_ ) );
BUF_X4 _16595_ ( .A(_08705_ ), .Z(_08860_ ) );
NAND3_X1 _16596_ ( .A1(_08860_ ), .A2(\RFU.rf[7][18] ), .A3(_08731_ ), .ZN(_08861_ ) );
NAND3_X1 _16597_ ( .A1(_08858_ ), .A2(\RFU.rf[5][18] ), .A3(_08748_ ), .ZN(_08862_ ) );
AND4_X1 _16598_ ( .A1(_08857_ ), .A2(_08859_ ), .A3(_08861_ ), .A4(_08862_ ), .ZN(_08863_ ) );
NAND3_X1 _16599_ ( .A1(_08716_ ), .A2(\RFU.rf[11][18] ), .A3(_08703_ ), .ZN(_08864_ ) );
NAND3_X1 _16600_ ( .A1(_08797_ ), .A2(_08733_ ), .A3(\RFU.rf[10][18] ), .ZN(_08865_ ) );
NAND3_X1 _16601_ ( .A1(_08710_ ), .A2(_08693_ ), .A3(\RFU.rf[9][18] ), .ZN(_08866_ ) );
BUF_X4 _16602_ ( .A(_08715_ ), .Z(_08867_ ) );
NAND3_X1 _16603_ ( .A1(_08867_ ), .A2(\RFU.rf[8][18] ), .A3(_08734_ ), .ZN(_08868_ ) );
AND4_X1 _16604_ ( .A1(_08864_ ), .A2(_08865_ ), .A3(_08866_ ), .A4(_08868_ ), .ZN(_08869_ ) );
NAND3_X1 _16605_ ( .A1(_08824_ ), .A2(\RFU.rf[14][18] ), .A3(_08739_ ), .ZN(_08870_ ) );
NAND3_X1 _16606_ ( .A1(_08710_ ), .A2(\RFU.rf[13][18] ), .A3(_08749_ ), .ZN(_08871_ ) );
NAND3_X1 _16607_ ( .A1(_08749_ ), .A2(\RFU.rf[12][18] ), .A3(_08723_ ), .ZN(_08872_ ) );
NAND3_X1 _16608_ ( .A1(_08749_ ), .A2(_08696_ ), .A3(\RFU.rf[15][18] ), .ZN(_08873_ ) );
AND4_X1 _16609_ ( .A1(_08870_ ), .A2(_08871_ ), .A3(_08872_ ), .A4(_08873_ ), .ZN(_08874_ ) );
NAND3_X1 _16610_ ( .A1(_08738_ ), .A2(\RFU.rf[2][18] ), .A3(_08758_ ), .ZN(_08875_ ) );
NAND3_X1 _16611_ ( .A1(_08756_ ), .A2(\RFU.rf[1][18] ), .A3(_08758_ ), .ZN(_08876_ ) );
NAND3_X1 _16612_ ( .A1(_08760_ ), .A2(\RFU.rf[3][18] ), .A3(_08761_ ), .ZN(_08877_ ) );
AND3_X1 _16613_ ( .A1(_08875_ ), .A2(_08876_ ), .A3(_08877_ ), .ZN(_08878_ ) );
NAND4_X1 _16614_ ( .A1(_08863_ ), .A2(_08869_ ), .A3(_08874_ ), .A4(_08878_ ), .ZN(_08879_ ) );
MUX2_X1 _16615_ ( .A(\EXU.r2_i [18] ), .B(_08879_ ), .S(_08765_ ), .Z(_00708_ ) );
NAND3_X1 _16616_ ( .A1(_08694_ ), .A2(\RFU.rf[11][17] ), .A3(_08697_ ), .ZN(_08880_ ) );
BUF_X4 _16617_ ( .A(_08702_ ), .Z(_08881_ ) );
NAND3_X1 _16618_ ( .A1(_08837_ ), .A2(\RFU.rf[7][17] ), .A3(_08881_ ), .ZN(_08882_ ) );
NAND3_X1 _16619_ ( .A1(_08860_ ), .A2(\RFU.rf[5][17] ), .A3(_08814_ ), .ZN(_08883_ ) );
NAND3_X1 _16620_ ( .A1(_08769_ ), .A2(_08716_ ), .A3(\RFU.rf[10][17] ), .ZN(_08884_ ) );
AND4_X1 _16621_ ( .A1(_08880_ ), .A2(_08882_ ), .A3(_08883_ ), .A4(_08884_ ), .ZN(_08885_ ) );
BUF_X4 _16622_ ( .A(_08723_ ), .Z(_08886_ ) );
NAND3_X1 _16623_ ( .A1(_08721_ ), .A2(\RFU.rf[12][17] ), .A3(_08886_ ), .ZN(_08887_ ) );
NAND3_X1 _16624_ ( .A1(_08797_ ), .A2(_08773_ ), .A3(\RFU.rf[6][17] ), .ZN(_08888_ ) );
NAND3_X1 _16625_ ( .A1(_08730_ ), .A2(_08820_ ), .A3(\RFU.rf[15][17] ), .ZN(_08889_ ) );
NAND3_X1 _16626_ ( .A1(_08867_ ), .A2(\RFU.rf[8][17] ), .A3(_08734_ ), .ZN(_08890_ ) );
AND4_X1 _16627_ ( .A1(_08887_ ), .A2(_08888_ ), .A3(_08889_ ), .A4(_08890_ ), .ZN(_08891_ ) );
NAND3_X1 _16628_ ( .A1(_08824_ ), .A2(\RFU.rf[14][17] ), .A3(_08739_ ), .ZN(_08892_ ) );
NAND3_X1 _16629_ ( .A1(_08741_ ), .A2(\RFU.rf[4][17] ), .A3(_08742_ ), .ZN(_08893_ ) );
NAND3_X1 _16630_ ( .A1(_08780_ ), .A2(\RFU.rf[2][17] ), .A3(_08827_ ), .ZN(_08894_ ) );
NAND3_X1 _16631_ ( .A1(_08782_ ), .A2(\RFU.rf[13][17] ), .A3(_08783_ ), .ZN(_08895_ ) );
AND4_X1 _16632_ ( .A1(_08892_ ), .A2(_08893_ ), .A3(_08894_ ), .A4(_08895_ ), .ZN(_08896_ ) );
NAND3_X1 _16633_ ( .A1(_08753_ ), .A2(_08754_ ), .A3(\RFU.rf[9][17] ), .ZN(_08897_ ) );
NAND3_X1 _16634_ ( .A1(_08756_ ), .A2(\RFU.rf[1][17] ), .A3(_08758_ ), .ZN(_08898_ ) );
NAND3_X1 _16635_ ( .A1(_08760_ ), .A2(\RFU.rf[3][17] ), .A3(_08761_ ), .ZN(_08899_ ) );
AND3_X1 _16636_ ( .A1(_08897_ ), .A2(_08898_ ), .A3(_08899_ ), .ZN(_08900_ ) );
NAND4_X1 _16637_ ( .A1(_08885_ ), .A2(_08891_ ), .A3(_08896_ ), .A4(_08900_ ), .ZN(_08901_ ) );
MUX2_X1 _16638_ ( .A(\EXU.r2_i [17] ), .B(_08901_ ), .S(_08765_ ), .Z(_00709_ ) );
BUF_X4 _16639_ ( .A(_08693_ ), .Z(_08902_ ) );
NAND3_X1 _16640_ ( .A1(_08902_ ), .A2(\RFU.rf[11][16] ), .A3(_08697_ ), .ZN(_08903_ ) );
NAND3_X1 _16641_ ( .A1(_08837_ ), .A2(\RFU.rf[7][16] ), .A3(_08881_ ), .ZN(_08904_ ) );
NAND3_X1 _16642_ ( .A1(_08860_ ), .A2(\RFU.rf[5][16] ), .A3(_08814_ ), .ZN(_08905_ ) );
BUF_X4 _16643_ ( .A(_08715_ ), .Z(_08906_ ) );
NAND3_X1 _16644_ ( .A1(_08769_ ), .A2(_08906_ ), .A3(\RFU.rf[10][16] ), .ZN(_08907_ ) );
AND4_X1 _16645_ ( .A1(_08903_ ), .A2(_08904_ ), .A3(_08905_ ), .A4(_08907_ ), .ZN(_08908_ ) );
BUF_X4 _16646_ ( .A(_08720_ ), .Z(_08909_ ) );
NAND3_X1 _16647_ ( .A1(_08909_ ), .A2(\RFU.rf[12][16] ), .A3(_08886_ ), .ZN(_08910_ ) );
NAND3_X1 _16648_ ( .A1(_08797_ ), .A2(_08773_ ), .A3(\RFU.rf[6][16] ), .ZN(_08911_ ) );
BUF_X4 _16649_ ( .A(_08729_ ), .Z(_08912_ ) );
NAND3_X1 _16650_ ( .A1(_08912_ ), .A2(_08820_ ), .A3(\RFU.rf[15][16] ), .ZN(_08913_ ) );
BUF_X4 _16651_ ( .A(_08722_ ), .Z(_08914_ ) );
NAND3_X1 _16652_ ( .A1(_08867_ ), .A2(\RFU.rf[8][16] ), .A3(_08914_ ), .ZN(_08915_ ) );
AND4_X1 _16653_ ( .A1(_08910_ ), .A2(_08911_ ), .A3(_08913_ ), .A4(_08915_ ), .ZN(_08916_ ) );
BUF_X4 _16654_ ( .A(_08729_ ), .Z(_08917_ ) );
NAND3_X1 _16655_ ( .A1(_08824_ ), .A2(\RFU.rf[14][16] ), .A3(_08917_ ), .ZN(_08918_ ) );
BUF_X4 _16656_ ( .A(_08722_ ), .Z(_08919_ ) );
NAND3_X1 _16657_ ( .A1(_08741_ ), .A2(\RFU.rf[4][16] ), .A3(_08919_ ), .ZN(_08920_ ) );
NAND3_X1 _16658_ ( .A1(_08780_ ), .A2(\RFU.rf[2][16] ), .A3(_08827_ ), .ZN(_08921_ ) );
NAND3_X1 _16659_ ( .A1(_08782_ ), .A2(\RFU.rf[13][16] ), .A3(_08783_ ), .ZN(_08922_ ) );
AND4_X1 _16660_ ( .A1(_08918_ ), .A2(_08920_ ), .A3(_08921_ ), .A4(_08922_ ), .ZN(_08923_ ) );
NAND3_X1 _16661_ ( .A1(_08753_ ), .A2(_08754_ ), .A3(\RFU.rf[9][16] ), .ZN(_08924_ ) );
NAND3_X1 _16662_ ( .A1(_08756_ ), .A2(\RFU.rf[1][16] ), .A3(_08758_ ), .ZN(_08925_ ) );
BUF_X4 _16663_ ( .A(_08745_ ), .Z(_08926_ ) );
NAND3_X1 _16664_ ( .A1(_08760_ ), .A2(\RFU.rf[3][16] ), .A3(_08926_ ), .ZN(_08927_ ) );
AND3_X1 _16665_ ( .A1(_08924_ ), .A2(_08925_ ), .A3(_08927_ ), .ZN(_08928_ ) );
NAND4_X1 _16666_ ( .A1(_08908_ ), .A2(_08916_ ), .A3(_08923_ ), .A4(_08928_ ), .ZN(_08929_ ) );
MUX2_X1 _16667_ ( .A(\EXU.r2_i [16] ), .B(_08929_ ), .S(_08765_ ), .Z(_00710_ ) );
NAND3_X1 _16668_ ( .A1(_08902_ ), .A2(\RFU.rf[11][15] ), .A3(_08697_ ), .ZN(_08930_ ) );
NAND3_X1 _16669_ ( .A1(_08837_ ), .A2(\RFU.rf[7][15] ), .A3(_08881_ ), .ZN(_08931_ ) );
NAND3_X1 _16670_ ( .A1(_08860_ ), .A2(\RFU.rf[5][15] ), .A3(_08814_ ), .ZN(_08932_ ) );
NAND3_X1 _16671_ ( .A1(_08769_ ), .A2(_08906_ ), .A3(\RFU.rf[10][15] ), .ZN(_08933_ ) );
AND4_X1 _16672_ ( .A1(_08930_ ), .A2(_08931_ ), .A3(_08932_ ), .A4(_08933_ ), .ZN(_08934_ ) );
NAND3_X1 _16673_ ( .A1(_08909_ ), .A2(\RFU.rf[12][15] ), .A3(_08886_ ), .ZN(_08935_ ) );
NAND3_X1 _16674_ ( .A1(_08797_ ), .A2(_08773_ ), .A3(\RFU.rf[6][15] ), .ZN(_08936_ ) );
NAND3_X1 _16675_ ( .A1(_08912_ ), .A2(_08820_ ), .A3(\RFU.rf[15][15] ), .ZN(_08937_ ) );
NAND3_X1 _16676_ ( .A1(_08867_ ), .A2(\RFU.rf[8][15] ), .A3(_08914_ ), .ZN(_08938_ ) );
AND4_X1 _16677_ ( .A1(_08935_ ), .A2(_08936_ ), .A3(_08937_ ), .A4(_08938_ ), .ZN(_08939_ ) );
NAND3_X1 _16678_ ( .A1(_08824_ ), .A2(\RFU.rf[14][15] ), .A3(_08917_ ), .ZN(_08940_ ) );
NAND3_X1 _16679_ ( .A1(_08741_ ), .A2(\RFU.rf[4][15] ), .A3(_08919_ ), .ZN(_08941_ ) );
NAND3_X1 _16680_ ( .A1(_08780_ ), .A2(\RFU.rf[2][15] ), .A3(_08827_ ), .ZN(_08942_ ) );
NAND3_X1 _16681_ ( .A1(_08782_ ), .A2(\RFU.rf[13][15] ), .A3(_08783_ ), .ZN(_08943_ ) );
AND4_X1 _16682_ ( .A1(_08940_ ), .A2(_08941_ ), .A3(_08942_ ), .A4(_08943_ ), .ZN(_08944_ ) );
BUF_X4 _16683_ ( .A(_08752_ ), .Z(_08945_ ) );
BUF_X4 _16684_ ( .A(_08715_ ), .Z(_08946_ ) );
NAND3_X1 _16685_ ( .A1(_08945_ ), .A2(_08946_ ), .A3(\RFU.rf[9][15] ), .ZN(_08947_ ) );
BUF_X4 _16686_ ( .A(_08709_ ), .Z(_08948_ ) );
BUF_X4 _16687_ ( .A(_08757_ ), .Z(_08949_ ) );
NAND3_X1 _16688_ ( .A1(_08948_ ), .A2(\RFU.rf[1][15] ), .A3(_08949_ ), .ZN(_08950_ ) );
NAND3_X1 _16689_ ( .A1(_08760_ ), .A2(\RFU.rf[3][15] ), .A3(_08926_ ), .ZN(_08951_ ) );
AND3_X1 _16690_ ( .A1(_08947_ ), .A2(_08950_ ), .A3(_08951_ ), .ZN(_08952_ ) );
NAND4_X1 _16691_ ( .A1(_08934_ ), .A2(_08939_ ), .A3(_08944_ ), .A4(_08952_ ), .ZN(_08953_ ) );
MUX2_X1 _16692_ ( .A(\EXU.r2_i [15] ), .B(_08953_ ), .S(_08765_ ), .Z(_00711_ ) );
BUF_X4 _16693_ ( .A(_08696_ ), .Z(_08954_ ) );
NAND3_X1 _16694_ ( .A1(_08902_ ), .A2(\RFU.rf[11][14] ), .A3(_08954_ ), .ZN(_08955_ ) );
NAND3_X1 _16695_ ( .A1(_08837_ ), .A2(\RFU.rf[7][14] ), .A3(_08881_ ), .ZN(_08956_ ) );
NAND3_X1 _16696_ ( .A1(_08860_ ), .A2(\RFU.rf[5][14] ), .A3(_08814_ ), .ZN(_08957_ ) );
NAND3_X1 _16697_ ( .A1(_08769_ ), .A2(_08906_ ), .A3(\RFU.rf[10][14] ), .ZN(_08958_ ) );
AND4_X1 _16698_ ( .A1(_08955_ ), .A2(_08956_ ), .A3(_08957_ ), .A4(_08958_ ), .ZN(_08959_ ) );
NAND3_X1 _16699_ ( .A1(_08909_ ), .A2(\RFU.rf[12][14] ), .A3(_08886_ ), .ZN(_08960_ ) );
NAND3_X1 _16700_ ( .A1(_08797_ ), .A2(_08773_ ), .A3(\RFU.rf[6][14] ), .ZN(_08961_ ) );
NAND3_X1 _16701_ ( .A1(_08912_ ), .A2(_08820_ ), .A3(\RFU.rf[15][14] ), .ZN(_08962_ ) );
NAND3_X1 _16702_ ( .A1(_08867_ ), .A2(\RFU.rf[8][14] ), .A3(_08914_ ), .ZN(_08963_ ) );
AND4_X1 _16703_ ( .A1(_08960_ ), .A2(_08961_ ), .A3(_08962_ ), .A4(_08963_ ), .ZN(_08964_ ) );
NAND3_X1 _16704_ ( .A1(_08824_ ), .A2(\RFU.rf[14][14] ), .A3(_08917_ ), .ZN(_08965_ ) );
NAND3_X1 _16705_ ( .A1(_08741_ ), .A2(\RFU.rf[4][14] ), .A3(_08919_ ), .ZN(_08966_ ) );
NAND3_X1 _16706_ ( .A1(_08780_ ), .A2(\RFU.rf[2][14] ), .A3(_08827_ ), .ZN(_08967_ ) );
NAND3_X1 _16707_ ( .A1(_08782_ ), .A2(\RFU.rf[13][14] ), .A3(_08783_ ), .ZN(_08968_ ) );
AND4_X1 _16708_ ( .A1(_08965_ ), .A2(_08966_ ), .A3(_08967_ ), .A4(_08968_ ), .ZN(_08969_ ) );
NAND3_X1 _16709_ ( .A1(_08945_ ), .A2(_08946_ ), .A3(\RFU.rf[9][14] ), .ZN(_08970_ ) );
NAND3_X1 _16710_ ( .A1(_08948_ ), .A2(\RFU.rf[1][14] ), .A3(_08949_ ), .ZN(_08971_ ) );
BUF_X4 _16711_ ( .A(_08702_ ), .Z(_08972_ ) );
NAND3_X1 _16712_ ( .A1(_08972_ ), .A2(\RFU.rf[3][14] ), .A3(_08926_ ), .ZN(_08973_ ) );
AND3_X1 _16713_ ( .A1(_08970_ ), .A2(_08971_ ), .A3(_08973_ ), .ZN(_08974_ ) );
NAND4_X1 _16714_ ( .A1(_08959_ ), .A2(_08964_ ), .A3(_08969_ ), .A4(_08974_ ), .ZN(_08975_ ) );
MUX2_X1 _16715_ ( .A(\EXU.r2_i [14] ), .B(_08975_ ), .S(_08765_ ), .Z(_00712_ ) );
NAND3_X1 _16716_ ( .A1(_08902_ ), .A2(\RFU.rf[11][13] ), .A3(_08954_ ), .ZN(_08976_ ) );
NAND3_X1 _16717_ ( .A1(_08837_ ), .A2(\RFU.rf[7][13] ), .A3(_08881_ ), .ZN(_08977_ ) );
NAND3_X1 _16718_ ( .A1(_08860_ ), .A2(\RFU.rf[5][13] ), .A3(_08814_ ), .ZN(_08978_ ) );
NAND3_X1 _16719_ ( .A1(_08769_ ), .A2(_08906_ ), .A3(\RFU.rf[10][13] ), .ZN(_08979_ ) );
AND4_X1 _16720_ ( .A1(_08976_ ), .A2(_08977_ ), .A3(_08978_ ), .A4(_08979_ ), .ZN(_08980_ ) );
NAND3_X1 _16721_ ( .A1(_08909_ ), .A2(\RFU.rf[12][13] ), .A3(_08886_ ), .ZN(_08981_ ) );
NAND3_X1 _16722_ ( .A1(_08797_ ), .A2(_08773_ ), .A3(\RFU.rf[6][13] ), .ZN(_08982_ ) );
NAND3_X1 _16723_ ( .A1(_08912_ ), .A2(_08820_ ), .A3(\RFU.rf[15][13] ), .ZN(_08983_ ) );
NAND3_X1 _16724_ ( .A1(_08867_ ), .A2(\RFU.rf[8][13] ), .A3(_08914_ ), .ZN(_08984_ ) );
AND4_X1 _16725_ ( .A1(_08981_ ), .A2(_08982_ ), .A3(_08983_ ), .A4(_08984_ ), .ZN(_08985_ ) );
NAND3_X1 _16726_ ( .A1(_08824_ ), .A2(\RFU.rf[14][13] ), .A3(_08917_ ), .ZN(_08986_ ) );
NAND3_X1 _16727_ ( .A1(_08741_ ), .A2(\RFU.rf[4][13] ), .A3(_08919_ ), .ZN(_08987_ ) );
NAND3_X1 _16728_ ( .A1(_08780_ ), .A2(\RFU.rf[2][13] ), .A3(_08827_ ), .ZN(_08988_ ) );
NAND3_X1 _16729_ ( .A1(_08782_ ), .A2(\RFU.rf[13][13] ), .A3(_08783_ ), .ZN(_08989_ ) );
AND4_X1 _16730_ ( .A1(_08986_ ), .A2(_08987_ ), .A3(_08988_ ), .A4(_08989_ ), .ZN(_08990_ ) );
NAND3_X1 _16731_ ( .A1(_08945_ ), .A2(_08946_ ), .A3(\RFU.rf[9][13] ), .ZN(_08991_ ) );
NAND3_X1 _16732_ ( .A1(_08948_ ), .A2(\RFU.rf[1][13] ), .A3(_08949_ ), .ZN(_08992_ ) );
NAND3_X1 _16733_ ( .A1(_08972_ ), .A2(\RFU.rf[3][13] ), .A3(_08926_ ), .ZN(_08993_ ) );
AND3_X1 _16734_ ( .A1(_08991_ ), .A2(_08992_ ), .A3(_08993_ ), .ZN(_08994_ ) );
NAND4_X1 _16735_ ( .A1(_08980_ ), .A2(_08985_ ), .A3(_08990_ ), .A4(_08994_ ), .ZN(_08995_ ) );
BUF_X4 _16736_ ( .A(_05514_ ), .Z(_08996_ ) );
MUX2_X1 _16737_ ( .A(\EXU.r2_i [13] ), .B(_08995_ ), .S(_08996_ ), .Z(_00713_ ) );
NAND3_X1 _16738_ ( .A1(_08902_ ), .A2(\RFU.rf[11][12] ), .A3(_08954_ ), .ZN(_08997_ ) );
NAND3_X1 _16739_ ( .A1(_08837_ ), .A2(\RFU.rf[7][12] ), .A3(_08881_ ), .ZN(_08998_ ) );
NAND3_X1 _16740_ ( .A1(_08860_ ), .A2(\RFU.rf[5][12] ), .A3(_08814_ ), .ZN(_08999_ ) );
NAND3_X1 _16741_ ( .A1(_08769_ ), .A2(_08906_ ), .A3(\RFU.rf[10][12] ), .ZN(_09000_ ) );
AND4_X1 _16742_ ( .A1(_08997_ ), .A2(_08998_ ), .A3(_08999_ ), .A4(_09000_ ), .ZN(_09001_ ) );
NAND3_X1 _16743_ ( .A1(_08909_ ), .A2(\RFU.rf[12][12] ), .A3(_08886_ ), .ZN(_09002_ ) );
NAND3_X1 _16744_ ( .A1(_08797_ ), .A2(_08773_ ), .A3(\RFU.rf[6][12] ), .ZN(_09003_ ) );
NAND3_X1 _16745_ ( .A1(_08912_ ), .A2(_08820_ ), .A3(\RFU.rf[15][12] ), .ZN(_09004_ ) );
NAND3_X1 _16746_ ( .A1(_08867_ ), .A2(\RFU.rf[8][12] ), .A3(_08914_ ), .ZN(_09005_ ) );
AND4_X1 _16747_ ( .A1(_09002_ ), .A2(_09003_ ), .A3(_09004_ ), .A4(_09005_ ), .ZN(_09006_ ) );
NAND3_X1 _16748_ ( .A1(_08824_ ), .A2(\RFU.rf[14][12] ), .A3(_08917_ ), .ZN(_09007_ ) );
BUF_X4 _16749_ ( .A(_08705_ ), .Z(_09008_ ) );
NAND3_X1 _16750_ ( .A1(_09008_ ), .A2(\RFU.rf[4][12] ), .A3(_08919_ ), .ZN(_09009_ ) );
NAND3_X1 _16751_ ( .A1(_08780_ ), .A2(\RFU.rf[2][12] ), .A3(_08827_ ), .ZN(_09010_ ) );
NAND3_X1 _16752_ ( .A1(_08782_ ), .A2(\RFU.rf[13][12] ), .A3(_08783_ ), .ZN(_09011_ ) );
AND4_X1 _16753_ ( .A1(_09007_ ), .A2(_09009_ ), .A3(_09010_ ), .A4(_09011_ ), .ZN(_09012_ ) );
NAND3_X1 _16754_ ( .A1(_08945_ ), .A2(_08946_ ), .A3(\RFU.rf[9][12] ), .ZN(_09013_ ) );
NAND3_X1 _16755_ ( .A1(_08948_ ), .A2(\RFU.rf[1][12] ), .A3(_08949_ ), .ZN(_09014_ ) );
NAND3_X1 _16756_ ( .A1(_08972_ ), .A2(\RFU.rf[3][12] ), .A3(_08926_ ), .ZN(_09015_ ) );
AND3_X1 _16757_ ( .A1(_09013_ ), .A2(_09014_ ), .A3(_09015_ ), .ZN(_09016_ ) );
NAND4_X1 _16758_ ( .A1(_09001_ ), .A2(_09006_ ), .A3(_09012_ ), .A4(_09016_ ), .ZN(_09017_ ) );
MUX2_X1 _16759_ ( .A(\EXU.r2_i [12] ), .B(_09017_ ), .S(_08996_ ), .Z(_00714_ ) );
NAND3_X1 _16760_ ( .A1(_08902_ ), .A2(\RFU.rf[11][29] ), .A3(_08954_ ), .ZN(_09018_ ) );
NAND3_X1 _16761_ ( .A1(_08837_ ), .A2(\RFU.rf[7][29] ), .A3(_08881_ ), .ZN(_09019_ ) );
NAND3_X1 _16762_ ( .A1(_08860_ ), .A2(\RFU.rf[5][29] ), .A3(_08814_ ), .ZN(_09020_ ) );
BUF_X4 _16763_ ( .A(_08713_ ), .Z(_09021_ ) );
NAND3_X1 _16764_ ( .A1(_09021_ ), .A2(_08906_ ), .A3(\RFU.rf[10][29] ), .ZN(_09022_ ) );
AND4_X1 _16765_ ( .A1(_09018_ ), .A2(_09019_ ), .A3(_09020_ ), .A4(_09022_ ), .ZN(_09023_ ) );
NAND3_X1 _16766_ ( .A1(_08909_ ), .A2(\RFU.rf[12][29] ), .A3(_08886_ ), .ZN(_09024_ ) );
BUF_X4 _16767_ ( .A(_08713_ ), .Z(_09025_ ) );
BUF_X4 _16768_ ( .A(_08705_ ), .Z(_09026_ ) );
NAND3_X1 _16769_ ( .A1(_09025_ ), .A2(_09026_ ), .A3(\RFU.rf[6][29] ), .ZN(_09027_ ) );
NAND3_X1 _16770_ ( .A1(_08912_ ), .A2(_08820_ ), .A3(\RFU.rf[15][29] ), .ZN(_09028_ ) );
NAND3_X1 _16771_ ( .A1(_08867_ ), .A2(\RFU.rf[8][29] ), .A3(_08914_ ), .ZN(_09029_ ) );
AND4_X1 _16772_ ( .A1(_09024_ ), .A2(_09027_ ), .A3(_09028_ ), .A4(_09029_ ), .ZN(_09030_ ) );
NAND3_X1 _16773_ ( .A1(_08824_ ), .A2(\RFU.rf[14][29] ), .A3(_08917_ ), .ZN(_09031_ ) );
NAND3_X1 _16774_ ( .A1(_09008_ ), .A2(\RFU.rf[4][29] ), .A3(_08919_ ), .ZN(_09032_ ) );
BUF_X4 _16775_ ( .A(_08713_ ), .Z(_09033_ ) );
NAND3_X1 _16776_ ( .A1(_09033_ ), .A2(\RFU.rf[2][29] ), .A3(_08827_ ), .ZN(_09034_ ) );
BUF_X4 _16777_ ( .A(_08709_ ), .Z(_09035_ ) );
BUF_X4 _16778_ ( .A(_08729_ ), .Z(_09036_ ) );
NAND3_X1 _16779_ ( .A1(_09035_ ), .A2(\RFU.rf[13][29] ), .A3(_09036_ ), .ZN(_09037_ ) );
AND4_X1 _16780_ ( .A1(_09031_ ), .A2(_09032_ ), .A3(_09034_ ), .A4(_09037_ ), .ZN(_09038_ ) );
NAND3_X1 _16781_ ( .A1(_08945_ ), .A2(_08946_ ), .A3(\RFU.rf[9][29] ), .ZN(_09039_ ) );
NAND3_X1 _16782_ ( .A1(_08948_ ), .A2(\RFU.rf[1][29] ), .A3(_08949_ ), .ZN(_09040_ ) );
NAND3_X1 _16783_ ( .A1(_08972_ ), .A2(\RFU.rf[3][29] ), .A3(_08926_ ), .ZN(_09041_ ) );
AND3_X1 _16784_ ( .A1(_09039_ ), .A2(_09040_ ), .A3(_09041_ ), .ZN(_09042_ ) );
NAND4_X1 _16785_ ( .A1(_09023_ ), .A2(_09030_ ), .A3(_09038_ ), .A4(_09042_ ), .ZN(_09043_ ) );
MUX2_X1 _16786_ ( .A(\EXU.r2_i [29] ), .B(_09043_ ), .S(_08996_ ), .Z(_00715_ ) );
NAND3_X1 _16787_ ( .A1(_08902_ ), .A2(\RFU.rf[11][11] ), .A3(_08954_ ), .ZN(_09044_ ) );
NAND3_X1 _16788_ ( .A1(_08837_ ), .A2(\RFU.rf[7][11] ), .A3(_08881_ ), .ZN(_09045_ ) );
NAND3_X1 _16789_ ( .A1(_08860_ ), .A2(\RFU.rf[5][11] ), .A3(_08814_ ), .ZN(_09046_ ) );
NAND3_X1 _16790_ ( .A1(_09021_ ), .A2(_08906_ ), .A3(\RFU.rf[10][11] ), .ZN(_09047_ ) );
AND4_X1 _16791_ ( .A1(_09044_ ), .A2(_09045_ ), .A3(_09046_ ), .A4(_09047_ ), .ZN(_09048_ ) );
NAND3_X1 _16792_ ( .A1(_08909_ ), .A2(\RFU.rf[12][11] ), .A3(_08886_ ), .ZN(_09049_ ) );
NAND3_X1 _16793_ ( .A1(_09025_ ), .A2(_09026_ ), .A3(\RFU.rf[6][11] ), .ZN(_09050_ ) );
NAND3_X1 _16794_ ( .A1(_08912_ ), .A2(_08820_ ), .A3(\RFU.rf[15][11] ), .ZN(_09051_ ) );
NAND3_X1 _16795_ ( .A1(_08867_ ), .A2(\RFU.rf[8][11] ), .A3(_08914_ ), .ZN(_09052_ ) );
AND4_X1 _16796_ ( .A1(_09049_ ), .A2(_09050_ ), .A3(_09051_ ), .A4(_09052_ ), .ZN(_09053_ ) );
BUF_X4 _16797_ ( .A(_08713_ ), .Z(_09054_ ) );
NAND3_X1 _16798_ ( .A1(_09054_ ), .A2(\RFU.rf[14][11] ), .A3(_08917_ ), .ZN(_09055_ ) );
NAND3_X1 _16799_ ( .A1(_09008_ ), .A2(\RFU.rf[4][11] ), .A3(_08919_ ), .ZN(_09056_ ) );
NAND3_X1 _16800_ ( .A1(_09033_ ), .A2(\RFU.rf[2][11] ), .A3(_08827_ ), .ZN(_09057_ ) );
NAND3_X1 _16801_ ( .A1(_09035_ ), .A2(\RFU.rf[13][11] ), .A3(_09036_ ), .ZN(_09058_ ) );
AND4_X1 _16802_ ( .A1(_09055_ ), .A2(_09056_ ), .A3(_09057_ ), .A4(_09058_ ), .ZN(_09059_ ) );
NAND3_X1 _16803_ ( .A1(_08945_ ), .A2(_08946_ ), .A3(\RFU.rf[9][11] ), .ZN(_09060_ ) );
NAND3_X1 _16804_ ( .A1(_08948_ ), .A2(\RFU.rf[1][11] ), .A3(_08949_ ), .ZN(_09061_ ) );
NAND3_X1 _16805_ ( .A1(_08972_ ), .A2(\RFU.rf[3][11] ), .A3(_08926_ ), .ZN(_09062_ ) );
AND3_X1 _16806_ ( .A1(_09060_ ), .A2(_09061_ ), .A3(_09062_ ), .ZN(_09063_ ) );
NAND4_X1 _16807_ ( .A1(_09048_ ), .A2(_09053_ ), .A3(_09059_ ), .A4(_09063_ ), .ZN(_09064_ ) );
MUX2_X1 _16808_ ( .A(\EXU.r2_i [11] ), .B(_09064_ ), .S(_08996_ ), .Z(_00716_ ) );
NAND3_X1 _16809_ ( .A1(_08902_ ), .A2(\RFU.rf[11][10] ), .A3(_08954_ ), .ZN(_09065_ ) );
NAND3_X1 _16810_ ( .A1(_08837_ ), .A2(\RFU.rf[7][10] ), .A3(_08881_ ), .ZN(_09066_ ) );
BUF_X4 _16811_ ( .A(_08709_ ), .Z(_09067_ ) );
NAND3_X1 _16812_ ( .A1(_08860_ ), .A2(\RFU.rf[5][10] ), .A3(_09067_ ), .ZN(_09068_ ) );
NAND3_X1 _16813_ ( .A1(_09021_ ), .A2(_08906_ ), .A3(\RFU.rf[10][10] ), .ZN(_09069_ ) );
AND4_X1 _16814_ ( .A1(_09065_ ), .A2(_09066_ ), .A3(_09068_ ), .A4(_09069_ ), .ZN(_09070_ ) );
NAND3_X1 _16815_ ( .A1(_08909_ ), .A2(\RFU.rf[12][10] ), .A3(_08886_ ), .ZN(_09071_ ) );
NAND3_X1 _16816_ ( .A1(_09025_ ), .A2(_09026_ ), .A3(\RFU.rf[6][10] ), .ZN(_09072_ ) );
BUF_X4 _16817_ ( .A(_08702_ ), .Z(_09073_ ) );
NAND3_X1 _16818_ ( .A1(_08912_ ), .A2(_09073_ ), .A3(\RFU.rf[15][10] ), .ZN(_09074_ ) );
NAND3_X1 _16819_ ( .A1(_08867_ ), .A2(\RFU.rf[8][10] ), .A3(_08914_ ), .ZN(_09075_ ) );
AND4_X1 _16820_ ( .A1(_09071_ ), .A2(_09072_ ), .A3(_09074_ ), .A4(_09075_ ), .ZN(_09076_ ) );
NAND3_X1 _16821_ ( .A1(_09054_ ), .A2(\RFU.rf[14][10] ), .A3(_08917_ ), .ZN(_09077_ ) );
NAND3_X1 _16822_ ( .A1(_09008_ ), .A2(\RFU.rf[4][10] ), .A3(_08919_ ), .ZN(_09078_ ) );
BUF_X4 _16823_ ( .A(_08745_ ), .Z(_09079_ ) );
NAND3_X1 _16824_ ( .A1(_09033_ ), .A2(\RFU.rf[2][10] ), .A3(_09079_ ), .ZN(_09080_ ) );
NAND3_X1 _16825_ ( .A1(_09035_ ), .A2(\RFU.rf[13][10] ), .A3(_09036_ ), .ZN(_09081_ ) );
AND4_X1 _16826_ ( .A1(_09077_ ), .A2(_09078_ ), .A3(_09080_ ), .A4(_09081_ ), .ZN(_09082_ ) );
NAND3_X1 _16827_ ( .A1(_08945_ ), .A2(_08946_ ), .A3(\RFU.rf[9][10] ), .ZN(_09083_ ) );
NAND3_X1 _16828_ ( .A1(_08948_ ), .A2(\RFU.rf[1][10] ), .A3(_08949_ ), .ZN(_09084_ ) );
NAND3_X1 _16829_ ( .A1(_08972_ ), .A2(\RFU.rf[3][10] ), .A3(_08926_ ), .ZN(_09085_ ) );
AND3_X1 _16830_ ( .A1(_09083_ ), .A2(_09084_ ), .A3(_09085_ ), .ZN(_09086_ ) );
NAND4_X1 _16831_ ( .A1(_09070_ ), .A2(_09076_ ), .A3(_09082_ ), .A4(_09086_ ), .ZN(_09087_ ) );
MUX2_X1 _16832_ ( .A(\EXU.r2_i [10] ), .B(_09087_ ), .S(_08996_ ), .Z(_00717_ ) );
NAND3_X1 _16833_ ( .A1(_08902_ ), .A2(\RFU.rf[11][9] ), .A3(_08954_ ), .ZN(_09088_ ) );
BUF_X4 _16834_ ( .A(_08705_ ), .Z(_09089_ ) );
NAND3_X1 _16835_ ( .A1(_09089_ ), .A2(\RFU.rf[7][9] ), .A3(_08881_ ), .ZN(_09090_ ) );
BUF_X4 _16836_ ( .A(_08705_ ), .Z(_09091_ ) );
NAND3_X1 _16837_ ( .A1(_09091_ ), .A2(\RFU.rf[5][9] ), .A3(_09067_ ), .ZN(_09092_ ) );
NAND3_X1 _16838_ ( .A1(_09021_ ), .A2(_08906_ ), .A3(\RFU.rf[10][9] ), .ZN(_09093_ ) );
AND4_X1 _16839_ ( .A1(_09088_ ), .A2(_09090_ ), .A3(_09092_ ), .A4(_09093_ ), .ZN(_09094_ ) );
NAND3_X1 _16840_ ( .A1(_08909_ ), .A2(\RFU.rf[12][9] ), .A3(_08886_ ), .ZN(_09095_ ) );
NAND3_X1 _16841_ ( .A1(_09025_ ), .A2(_09026_ ), .A3(\RFU.rf[6][9] ), .ZN(_09096_ ) );
NAND3_X1 _16842_ ( .A1(_08912_ ), .A2(_09073_ ), .A3(\RFU.rf[15][9] ), .ZN(_09097_ ) );
BUF_X4 _16843_ ( .A(_08715_ ), .Z(_09098_ ) );
NAND3_X1 _16844_ ( .A1(_09098_ ), .A2(\RFU.rf[8][9] ), .A3(_08914_ ), .ZN(_09099_ ) );
AND4_X1 _16845_ ( .A1(_09095_ ), .A2(_09096_ ), .A3(_09097_ ), .A4(_09099_ ), .ZN(_09100_ ) );
NAND3_X1 _16846_ ( .A1(_09054_ ), .A2(\RFU.rf[14][9] ), .A3(_08917_ ), .ZN(_09101_ ) );
NAND3_X1 _16847_ ( .A1(_09008_ ), .A2(\RFU.rf[4][9] ), .A3(_08919_ ), .ZN(_09102_ ) );
NAND3_X1 _16848_ ( .A1(_09033_ ), .A2(\RFU.rf[2][9] ), .A3(_09079_ ), .ZN(_09103_ ) );
NAND3_X1 _16849_ ( .A1(_09035_ ), .A2(\RFU.rf[13][9] ), .A3(_09036_ ), .ZN(_09104_ ) );
AND4_X1 _16850_ ( .A1(_09101_ ), .A2(_09102_ ), .A3(_09103_ ), .A4(_09104_ ), .ZN(_09105_ ) );
NAND3_X1 _16851_ ( .A1(_08945_ ), .A2(_08946_ ), .A3(\RFU.rf[9][9] ), .ZN(_09106_ ) );
NAND3_X1 _16852_ ( .A1(_08948_ ), .A2(\RFU.rf[1][9] ), .A3(_08949_ ), .ZN(_09107_ ) );
NAND3_X1 _16853_ ( .A1(_08972_ ), .A2(\RFU.rf[3][9] ), .A3(_08926_ ), .ZN(_09108_ ) );
AND3_X1 _16854_ ( .A1(_09106_ ), .A2(_09107_ ), .A3(_09108_ ), .ZN(_09109_ ) );
NAND4_X1 _16855_ ( .A1(_09094_ ), .A2(_09100_ ), .A3(_09105_ ), .A4(_09109_ ), .ZN(_09110_ ) );
MUX2_X1 _16856_ ( .A(\EXU.r2_i [9] ), .B(_09110_ ), .S(_08996_ ), .Z(_00718_ ) );
NAND3_X1 _16857_ ( .A1(_08902_ ), .A2(\RFU.rf[11][8] ), .A3(_08954_ ), .ZN(_09111_ ) );
BUF_X4 _16858_ ( .A(_08702_ ), .Z(_09112_ ) );
NAND3_X1 _16859_ ( .A1(_09089_ ), .A2(\RFU.rf[7][8] ), .A3(_09112_ ), .ZN(_09113_ ) );
NAND3_X1 _16860_ ( .A1(_09091_ ), .A2(\RFU.rf[5][8] ), .A3(_09067_ ), .ZN(_09114_ ) );
NAND3_X1 _16861_ ( .A1(_09021_ ), .A2(_08906_ ), .A3(\RFU.rf[10][8] ), .ZN(_09115_ ) );
AND4_X1 _16862_ ( .A1(_09111_ ), .A2(_09113_ ), .A3(_09114_ ), .A4(_09115_ ), .ZN(_09116_ ) );
BUF_X4 _16863_ ( .A(_08723_ ), .Z(_09117_ ) );
NAND3_X1 _16864_ ( .A1(_08909_ ), .A2(\RFU.rf[12][8] ), .A3(_09117_ ), .ZN(_09118_ ) );
NAND3_X1 _16865_ ( .A1(_09025_ ), .A2(_09026_ ), .A3(\RFU.rf[6][8] ), .ZN(_09119_ ) );
NAND3_X1 _16866_ ( .A1(_08912_ ), .A2(_09073_ ), .A3(\RFU.rf[15][8] ), .ZN(_09120_ ) );
NAND3_X1 _16867_ ( .A1(_09098_ ), .A2(\RFU.rf[8][8] ), .A3(_08914_ ), .ZN(_09121_ ) );
AND4_X1 _16868_ ( .A1(_09118_ ), .A2(_09119_ ), .A3(_09120_ ), .A4(_09121_ ), .ZN(_09122_ ) );
NAND3_X1 _16869_ ( .A1(_09054_ ), .A2(\RFU.rf[14][8] ), .A3(_08917_ ), .ZN(_09123_ ) );
NAND3_X1 _16870_ ( .A1(_09008_ ), .A2(\RFU.rf[4][8] ), .A3(_08919_ ), .ZN(_09124_ ) );
NAND3_X1 _16871_ ( .A1(_09033_ ), .A2(\RFU.rf[2][8] ), .A3(_09079_ ), .ZN(_09125_ ) );
NAND3_X1 _16872_ ( .A1(_09035_ ), .A2(\RFU.rf[13][8] ), .A3(_09036_ ), .ZN(_09126_ ) );
AND4_X1 _16873_ ( .A1(_09123_ ), .A2(_09124_ ), .A3(_09125_ ), .A4(_09126_ ), .ZN(_09127_ ) );
NAND3_X1 _16874_ ( .A1(_08945_ ), .A2(_08946_ ), .A3(\RFU.rf[9][8] ), .ZN(_09128_ ) );
NAND3_X1 _16875_ ( .A1(_08948_ ), .A2(\RFU.rf[1][8] ), .A3(_08949_ ), .ZN(_09129_ ) );
NAND3_X1 _16876_ ( .A1(_08972_ ), .A2(\RFU.rf[3][8] ), .A3(_08926_ ), .ZN(_09130_ ) );
AND3_X1 _16877_ ( .A1(_09128_ ), .A2(_09129_ ), .A3(_09130_ ), .ZN(_09131_ ) );
NAND4_X1 _16878_ ( .A1(_09116_ ), .A2(_09122_ ), .A3(_09127_ ), .A4(_09131_ ), .ZN(_09132_ ) );
MUX2_X1 _16879_ ( .A(\EXU.r2_i [8] ), .B(_09132_ ), .S(_08996_ ), .Z(_00719_ ) );
BUF_X4 _16880_ ( .A(_08715_ ), .Z(_09133_ ) );
NAND3_X1 _16881_ ( .A1(_09133_ ), .A2(\RFU.rf[11][7] ), .A3(_08954_ ), .ZN(_09134_ ) );
NAND3_X1 _16882_ ( .A1(_09089_ ), .A2(\RFU.rf[7][7] ), .A3(_09112_ ), .ZN(_09135_ ) );
NAND3_X1 _16883_ ( .A1(_09091_ ), .A2(\RFU.rf[5][7] ), .A3(_09067_ ), .ZN(_09136_ ) );
BUF_X4 _16884_ ( .A(_08715_ ), .Z(_09137_ ) );
NAND3_X1 _16885_ ( .A1(_09021_ ), .A2(_09137_ ), .A3(\RFU.rf[10][7] ), .ZN(_09138_ ) );
AND4_X1 _16886_ ( .A1(_09134_ ), .A2(_09135_ ), .A3(_09136_ ), .A4(_09138_ ), .ZN(_09139_ ) );
BUF_X4 _16887_ ( .A(_08729_ ), .Z(_09140_ ) );
NAND3_X1 _16888_ ( .A1(_09140_ ), .A2(\RFU.rf[12][7] ), .A3(_09117_ ), .ZN(_09141_ ) );
NAND3_X1 _16889_ ( .A1(_09025_ ), .A2(_09026_ ), .A3(\RFU.rf[6][7] ), .ZN(_09142_ ) );
BUF_X4 _16890_ ( .A(_08729_ ), .Z(_09143_ ) );
NAND3_X1 _16891_ ( .A1(_09143_ ), .A2(_09073_ ), .A3(\RFU.rf[15][7] ), .ZN(_09144_ ) );
BUF_X4 _16892_ ( .A(_08722_ ), .Z(_09145_ ) );
NAND3_X1 _16893_ ( .A1(_09098_ ), .A2(\RFU.rf[8][7] ), .A3(_09145_ ), .ZN(_09146_ ) );
AND4_X1 _16894_ ( .A1(_09141_ ), .A2(_09142_ ), .A3(_09144_ ), .A4(_09146_ ), .ZN(_09147_ ) );
BUF_X4 _16895_ ( .A(_08729_ ), .Z(_09148_ ) );
NAND3_X1 _16896_ ( .A1(_09054_ ), .A2(\RFU.rf[14][7] ), .A3(_09148_ ), .ZN(_09149_ ) );
BUF_X4 _16897_ ( .A(_08722_ ), .Z(_09150_ ) );
NAND3_X1 _16898_ ( .A1(_09008_ ), .A2(\RFU.rf[4][7] ), .A3(_09150_ ), .ZN(_09151_ ) );
NAND3_X1 _16899_ ( .A1(_09033_ ), .A2(\RFU.rf[2][7] ), .A3(_09079_ ), .ZN(_09152_ ) );
NAND3_X1 _16900_ ( .A1(_09035_ ), .A2(\RFU.rf[13][7] ), .A3(_09036_ ), .ZN(_09153_ ) );
AND4_X1 _16901_ ( .A1(_09149_ ), .A2(_09151_ ), .A3(_09152_ ), .A4(_09153_ ), .ZN(_09154_ ) );
NAND3_X1 _16902_ ( .A1(_08945_ ), .A2(_08946_ ), .A3(\RFU.rf[9][7] ), .ZN(_09155_ ) );
NAND3_X1 _16903_ ( .A1(_08948_ ), .A2(\RFU.rf[1][7] ), .A3(_08949_ ), .ZN(_09156_ ) );
BUF_X4 _16904_ ( .A(_08745_ ), .Z(_09157_ ) );
NAND3_X1 _16905_ ( .A1(_08972_ ), .A2(\RFU.rf[3][7] ), .A3(_09157_ ), .ZN(_09158_ ) );
AND3_X1 _16906_ ( .A1(_09155_ ), .A2(_09156_ ), .A3(_09158_ ), .ZN(_09159_ ) );
NAND4_X1 _16907_ ( .A1(_09139_ ), .A2(_09147_ ), .A3(_09154_ ), .A4(_09159_ ), .ZN(_09160_ ) );
MUX2_X1 _16908_ ( .A(\EXU.r2_i [7] ), .B(_09160_ ), .S(_08996_ ), .Z(_00720_ ) );
NAND3_X1 _16909_ ( .A1(_09133_ ), .A2(\RFU.rf[11][6] ), .A3(_08954_ ), .ZN(_09161_ ) );
NAND3_X1 _16910_ ( .A1(_09089_ ), .A2(\RFU.rf[7][6] ), .A3(_09112_ ), .ZN(_09162_ ) );
NAND3_X1 _16911_ ( .A1(_09091_ ), .A2(\RFU.rf[5][6] ), .A3(_09067_ ), .ZN(_09163_ ) );
NAND3_X1 _16912_ ( .A1(_09021_ ), .A2(_09137_ ), .A3(\RFU.rf[10][6] ), .ZN(_09164_ ) );
AND4_X1 _16913_ ( .A1(_09161_ ), .A2(_09162_ ), .A3(_09163_ ), .A4(_09164_ ), .ZN(_09165_ ) );
NAND3_X1 _16914_ ( .A1(_09140_ ), .A2(\RFU.rf[12][6] ), .A3(_09117_ ), .ZN(_09166_ ) );
NAND3_X1 _16915_ ( .A1(_09025_ ), .A2(_09026_ ), .A3(\RFU.rf[6][6] ), .ZN(_09167_ ) );
NAND3_X1 _16916_ ( .A1(_09143_ ), .A2(_09073_ ), .A3(\RFU.rf[15][6] ), .ZN(_09168_ ) );
NAND3_X1 _16917_ ( .A1(_09098_ ), .A2(\RFU.rf[8][6] ), .A3(_09145_ ), .ZN(_09169_ ) );
AND4_X1 _16918_ ( .A1(_09166_ ), .A2(_09167_ ), .A3(_09168_ ), .A4(_09169_ ), .ZN(_09170_ ) );
NAND3_X1 _16919_ ( .A1(_09054_ ), .A2(\RFU.rf[14][6] ), .A3(_09148_ ), .ZN(_09171_ ) );
NAND3_X1 _16920_ ( .A1(_09008_ ), .A2(\RFU.rf[4][6] ), .A3(_09150_ ), .ZN(_09172_ ) );
NAND3_X1 _16921_ ( .A1(_09033_ ), .A2(\RFU.rf[2][6] ), .A3(_09079_ ), .ZN(_09173_ ) );
NAND3_X1 _16922_ ( .A1(_09035_ ), .A2(\RFU.rf[13][6] ), .A3(_09036_ ), .ZN(_09174_ ) );
AND4_X1 _16923_ ( .A1(_09171_ ), .A2(_09172_ ), .A3(_09173_ ), .A4(_09174_ ), .ZN(_09175_ ) );
BUF_X4 _16924_ ( .A(_08709_ ), .Z(_09176_ ) );
BUF_X4 _16925_ ( .A(_08715_ ), .Z(_09177_ ) );
NAND3_X1 _16926_ ( .A1(_09176_ ), .A2(_09177_ ), .A3(\RFU.rf[9][6] ), .ZN(_09178_ ) );
BUF_X4 _16927_ ( .A(_08709_ ), .Z(_09179_ ) );
BUF_X4 _16928_ ( .A(_08757_ ), .Z(_09180_ ) );
NAND3_X1 _16929_ ( .A1(_09179_ ), .A2(\RFU.rf[1][6] ), .A3(_09180_ ), .ZN(_09181_ ) );
NAND3_X1 _16930_ ( .A1(_08972_ ), .A2(\RFU.rf[3][6] ), .A3(_09157_ ), .ZN(_09182_ ) );
AND3_X1 _16931_ ( .A1(_09178_ ), .A2(_09181_ ), .A3(_09182_ ), .ZN(_09183_ ) );
NAND4_X1 _16932_ ( .A1(_09165_ ), .A2(_09170_ ), .A3(_09175_ ), .A4(_09183_ ), .ZN(_09184_ ) );
MUX2_X1 _16933_ ( .A(\EXU.r2_i [6] ), .B(_09184_ ), .S(_08996_ ), .Z(_00721_ ) );
BUF_X4 _16934_ ( .A(_08702_ ), .Z(_09185_ ) );
NAND3_X1 _16935_ ( .A1(_09133_ ), .A2(\RFU.rf[11][5] ), .A3(_09185_ ), .ZN(_09186_ ) );
NAND3_X1 _16936_ ( .A1(_09089_ ), .A2(\RFU.rf[7][5] ), .A3(_09112_ ), .ZN(_09187_ ) );
NAND3_X1 _16937_ ( .A1(_09091_ ), .A2(\RFU.rf[5][5] ), .A3(_09067_ ), .ZN(_09188_ ) );
NAND3_X1 _16938_ ( .A1(_09021_ ), .A2(_09137_ ), .A3(\RFU.rf[10][5] ), .ZN(_09189_ ) );
AND4_X1 _16939_ ( .A1(_09186_ ), .A2(_09187_ ), .A3(_09188_ ), .A4(_09189_ ), .ZN(_09190_ ) );
NAND3_X1 _16940_ ( .A1(_09140_ ), .A2(\RFU.rf[12][5] ), .A3(_09117_ ), .ZN(_09191_ ) );
NAND3_X1 _16941_ ( .A1(_09025_ ), .A2(_09026_ ), .A3(\RFU.rf[6][5] ), .ZN(_09192_ ) );
NAND3_X1 _16942_ ( .A1(_09143_ ), .A2(_09073_ ), .A3(\RFU.rf[15][5] ), .ZN(_09193_ ) );
NAND3_X1 _16943_ ( .A1(_09098_ ), .A2(\RFU.rf[8][5] ), .A3(_09145_ ), .ZN(_09194_ ) );
AND4_X1 _16944_ ( .A1(_09191_ ), .A2(_09192_ ), .A3(_09193_ ), .A4(_09194_ ), .ZN(_09195_ ) );
NAND3_X1 _16945_ ( .A1(_09054_ ), .A2(\RFU.rf[14][5] ), .A3(_09148_ ), .ZN(_09196_ ) );
NAND3_X1 _16946_ ( .A1(_09008_ ), .A2(\RFU.rf[4][5] ), .A3(_09150_ ), .ZN(_09197_ ) );
NAND3_X1 _16947_ ( .A1(_09033_ ), .A2(\RFU.rf[2][5] ), .A3(_09079_ ), .ZN(_09198_ ) );
NAND3_X1 _16948_ ( .A1(_09035_ ), .A2(\RFU.rf[13][5] ), .A3(_09036_ ), .ZN(_09199_ ) );
AND4_X1 _16949_ ( .A1(_09196_ ), .A2(_09197_ ), .A3(_09198_ ), .A4(_09199_ ), .ZN(_09200_ ) );
NAND3_X1 _16950_ ( .A1(_09176_ ), .A2(_09177_ ), .A3(\RFU.rf[9][5] ), .ZN(_09201_ ) );
NAND3_X1 _16951_ ( .A1(_09179_ ), .A2(\RFU.rf[1][5] ), .A3(_09180_ ), .ZN(_09202_ ) );
BUF_X4 _16952_ ( .A(_08702_ ), .Z(_09203_ ) );
NAND3_X1 _16953_ ( .A1(_09203_ ), .A2(\RFU.rf[3][5] ), .A3(_09157_ ), .ZN(_09204_ ) );
AND3_X1 _16954_ ( .A1(_09201_ ), .A2(_09202_ ), .A3(_09204_ ), .ZN(_09205_ ) );
NAND4_X1 _16955_ ( .A1(_09190_ ), .A2(_09195_ ), .A3(_09200_ ), .A4(_09205_ ), .ZN(_09206_ ) );
MUX2_X1 _16956_ ( .A(\EXU.r2_i [5] ), .B(_09206_ ), .S(_08996_ ), .Z(_00722_ ) );
NAND3_X1 _16957_ ( .A1(_09133_ ), .A2(\RFU.rf[11][4] ), .A3(_09185_ ), .ZN(_09207_ ) );
NAND3_X1 _16958_ ( .A1(_09089_ ), .A2(\RFU.rf[7][4] ), .A3(_09112_ ), .ZN(_09208_ ) );
NAND3_X1 _16959_ ( .A1(_09091_ ), .A2(\RFU.rf[5][4] ), .A3(_09067_ ), .ZN(_09209_ ) );
NAND3_X1 _16960_ ( .A1(_09021_ ), .A2(_09137_ ), .A3(\RFU.rf[10][4] ), .ZN(_09210_ ) );
AND4_X1 _16961_ ( .A1(_09207_ ), .A2(_09208_ ), .A3(_09209_ ), .A4(_09210_ ), .ZN(_09211_ ) );
NAND3_X1 _16962_ ( .A1(_09140_ ), .A2(\RFU.rf[12][4] ), .A3(_09117_ ), .ZN(_09212_ ) );
NAND3_X1 _16963_ ( .A1(_09025_ ), .A2(_09026_ ), .A3(\RFU.rf[6][4] ), .ZN(_09213_ ) );
NAND3_X1 _16964_ ( .A1(_09143_ ), .A2(_09073_ ), .A3(\RFU.rf[15][4] ), .ZN(_09214_ ) );
NAND3_X1 _16965_ ( .A1(_09098_ ), .A2(\RFU.rf[8][4] ), .A3(_09145_ ), .ZN(_09215_ ) );
AND4_X1 _16966_ ( .A1(_09212_ ), .A2(_09213_ ), .A3(_09214_ ), .A4(_09215_ ), .ZN(_09216_ ) );
NAND3_X1 _16967_ ( .A1(_09054_ ), .A2(\RFU.rf[14][4] ), .A3(_09148_ ), .ZN(_09217_ ) );
NAND3_X1 _16968_ ( .A1(_09008_ ), .A2(\RFU.rf[4][4] ), .A3(_09150_ ), .ZN(_09218_ ) );
NAND3_X1 _16969_ ( .A1(_09033_ ), .A2(\RFU.rf[2][4] ), .A3(_09079_ ), .ZN(_09219_ ) );
NAND3_X1 _16970_ ( .A1(_09035_ ), .A2(\RFU.rf[13][4] ), .A3(_09036_ ), .ZN(_09220_ ) );
AND4_X1 _16971_ ( .A1(_09217_ ), .A2(_09218_ ), .A3(_09219_ ), .A4(_09220_ ), .ZN(_09221_ ) );
NAND3_X1 _16972_ ( .A1(_09176_ ), .A2(_09177_ ), .A3(\RFU.rf[9][4] ), .ZN(_09222_ ) );
NAND3_X1 _16973_ ( .A1(_09179_ ), .A2(\RFU.rf[1][4] ), .A3(_09180_ ), .ZN(_09223_ ) );
NAND3_X1 _16974_ ( .A1(_09203_ ), .A2(\RFU.rf[3][4] ), .A3(_09157_ ), .ZN(_09224_ ) );
AND3_X1 _16975_ ( .A1(_09222_ ), .A2(_09223_ ), .A3(_09224_ ), .ZN(_09225_ ) );
NAND4_X1 _16976_ ( .A1(_09211_ ), .A2(_09216_ ), .A3(_09221_ ), .A4(_09225_ ), .ZN(_09226_ ) );
BUF_X4 _16977_ ( .A(_05514_ ), .Z(_09227_ ) );
MUX2_X1 _16978_ ( .A(\EXU.r2_i [4] ), .B(_09226_ ), .S(_09227_ ), .Z(_00723_ ) );
NAND3_X1 _16979_ ( .A1(_09133_ ), .A2(\RFU.rf[11][3] ), .A3(_09185_ ), .ZN(_09228_ ) );
NAND3_X1 _16980_ ( .A1(_09089_ ), .A2(\RFU.rf[7][3] ), .A3(_09112_ ), .ZN(_09229_ ) );
NAND3_X1 _16981_ ( .A1(_09091_ ), .A2(\RFU.rf[5][3] ), .A3(_09067_ ), .ZN(_09230_ ) );
NAND3_X1 _16982_ ( .A1(_09021_ ), .A2(_09137_ ), .A3(\RFU.rf[10][3] ), .ZN(_09231_ ) );
AND4_X1 _16983_ ( .A1(_09228_ ), .A2(_09229_ ), .A3(_09230_ ), .A4(_09231_ ), .ZN(_09232_ ) );
NAND3_X1 _16984_ ( .A1(_09140_ ), .A2(\RFU.rf[12][3] ), .A3(_09117_ ), .ZN(_09233_ ) );
NAND3_X1 _16985_ ( .A1(_09025_ ), .A2(_09026_ ), .A3(\RFU.rf[6][3] ), .ZN(_09234_ ) );
NAND3_X1 _16986_ ( .A1(_09143_ ), .A2(_09073_ ), .A3(\RFU.rf[15][3] ), .ZN(_09235_ ) );
NAND3_X1 _16987_ ( .A1(_09098_ ), .A2(\RFU.rf[8][3] ), .A3(_09145_ ), .ZN(_09236_ ) );
AND4_X1 _16988_ ( .A1(_09233_ ), .A2(_09234_ ), .A3(_09235_ ), .A4(_09236_ ), .ZN(_09237_ ) );
NAND3_X1 _16989_ ( .A1(_09054_ ), .A2(\RFU.rf[14][3] ), .A3(_09148_ ), .ZN(_09238_ ) );
NAND3_X1 _16990_ ( .A1(_08727_ ), .A2(\RFU.rf[4][3] ), .A3(_09150_ ), .ZN(_09239_ ) );
NAND3_X1 _16991_ ( .A1(_09033_ ), .A2(\RFU.rf[2][3] ), .A3(_09079_ ), .ZN(_09240_ ) );
NAND3_X1 _16992_ ( .A1(_09035_ ), .A2(\RFU.rf[13][3] ), .A3(_09036_ ), .ZN(_09241_ ) );
AND4_X1 _16993_ ( .A1(_09238_ ), .A2(_09239_ ), .A3(_09240_ ), .A4(_09241_ ), .ZN(_09242_ ) );
NAND3_X1 _16994_ ( .A1(_09176_ ), .A2(_09177_ ), .A3(\RFU.rf[9][3] ), .ZN(_09243_ ) );
NAND3_X1 _16995_ ( .A1(_09179_ ), .A2(\RFU.rf[1][3] ), .A3(_09180_ ), .ZN(_09244_ ) );
NAND3_X1 _16996_ ( .A1(_09203_ ), .A2(\RFU.rf[3][3] ), .A3(_09157_ ), .ZN(_09245_ ) );
AND3_X1 _16997_ ( .A1(_09243_ ), .A2(_09244_ ), .A3(_09245_ ), .ZN(_09246_ ) );
NAND4_X1 _16998_ ( .A1(_09232_ ), .A2(_09237_ ), .A3(_09242_ ), .A4(_09246_ ), .ZN(_09247_ ) );
MUX2_X1 _16999_ ( .A(\EXU.r2_i [3] ), .B(_09247_ ), .S(_09227_ ), .Z(_00724_ ) );
NAND3_X1 _17000_ ( .A1(_09133_ ), .A2(\RFU.rf[11][2] ), .A3(_09185_ ), .ZN(_09248_ ) );
NAND3_X1 _17001_ ( .A1(_09089_ ), .A2(\RFU.rf[7][2] ), .A3(_09112_ ), .ZN(_09249_ ) );
NAND3_X1 _17002_ ( .A1(_09091_ ), .A2(\RFU.rf[5][2] ), .A3(_09067_ ), .ZN(_09250_ ) );
NAND3_X1 _17003_ ( .A1(_08726_ ), .A2(_09137_ ), .A3(\RFU.rf[10][2] ), .ZN(_09251_ ) );
AND4_X1 _17004_ ( .A1(_09248_ ), .A2(_09249_ ), .A3(_09250_ ), .A4(_09251_ ), .ZN(_09252_ ) );
NAND3_X1 _17005_ ( .A1(_09140_ ), .A2(\RFU.rf[12][2] ), .A3(_09117_ ), .ZN(_09253_ ) );
NAND3_X1 _17006_ ( .A1(_08744_ ), .A2(_08700_ ), .A3(\RFU.rf[6][2] ), .ZN(_09254_ ) );
NAND3_X1 _17007_ ( .A1(_09143_ ), .A2(_09073_ ), .A3(\RFU.rf[15][2] ), .ZN(_09255_ ) );
NAND3_X1 _17008_ ( .A1(_09098_ ), .A2(\RFU.rf[8][2] ), .A3(_09145_ ), .ZN(_09256_ ) );
AND4_X1 _17009_ ( .A1(_09253_ ), .A2(_09254_ ), .A3(_09255_ ), .A4(_09256_ ), .ZN(_09257_ ) );
NAND3_X1 _17010_ ( .A1(_09054_ ), .A2(\RFU.rf[14][2] ), .A3(_09148_ ), .ZN(_09258_ ) );
NAND3_X1 _17011_ ( .A1(_08727_ ), .A2(\RFU.rf[4][2] ), .A3(_09150_ ), .ZN(_09259_ ) );
NAND3_X1 _17012_ ( .A1(_08737_ ), .A2(\RFU.rf[2][2] ), .A3(_09079_ ), .ZN(_09260_ ) );
NAND3_X1 _17013_ ( .A1(_08752_ ), .A2(\RFU.rf[13][2] ), .A3(_08720_ ), .ZN(_09261_ ) );
AND4_X1 _17014_ ( .A1(_09258_ ), .A2(_09259_ ), .A3(_09260_ ), .A4(_09261_ ), .ZN(_09262_ ) );
NAND3_X1 _17015_ ( .A1(_09176_ ), .A2(_09177_ ), .A3(\RFU.rf[9][2] ), .ZN(_09263_ ) );
NAND3_X1 _17016_ ( .A1(_09179_ ), .A2(\RFU.rf[1][2] ), .A3(_09180_ ), .ZN(_09264_ ) );
NAND3_X1 _17017_ ( .A1(_09203_ ), .A2(\RFU.rf[3][2] ), .A3(_09157_ ), .ZN(_09265_ ) );
AND3_X1 _17018_ ( .A1(_09263_ ), .A2(_09264_ ), .A3(_09265_ ), .ZN(_09266_ ) );
NAND4_X1 _17019_ ( .A1(_09252_ ), .A2(_09257_ ), .A3(_09262_ ), .A4(_09266_ ), .ZN(_09267_ ) );
MUX2_X1 _17020_ ( .A(\EXU.r2_i [2] ), .B(_09267_ ), .S(_09227_ ), .Z(_00725_ ) );
NAND3_X1 _17021_ ( .A1(_09133_ ), .A2(\RFU.rf[11][28] ), .A3(_09185_ ), .ZN(_09268_ ) );
NAND3_X1 _17022_ ( .A1(_09089_ ), .A2(\RFU.rf[7][28] ), .A3(_09112_ ), .ZN(_09269_ ) );
NAND3_X1 _17023_ ( .A1(_09091_ ), .A2(\RFU.rf[5][28] ), .A3(_09067_ ), .ZN(_09270_ ) );
NAND3_X1 _17024_ ( .A1(_08726_ ), .A2(_09137_ ), .A3(\RFU.rf[10][28] ), .ZN(_09271_ ) );
AND4_X1 _17025_ ( .A1(_09268_ ), .A2(_09269_ ), .A3(_09270_ ), .A4(_09271_ ), .ZN(_09272_ ) );
NAND3_X1 _17026_ ( .A1(_09140_ ), .A2(\RFU.rf[12][28] ), .A3(_09117_ ), .ZN(_09273_ ) );
NAND3_X1 _17027_ ( .A1(_08744_ ), .A2(_08700_ ), .A3(\RFU.rf[6][28] ), .ZN(_09274_ ) );
NAND3_X1 _17028_ ( .A1(_09143_ ), .A2(_09073_ ), .A3(\RFU.rf[15][28] ), .ZN(_09275_ ) );
NAND3_X1 _17029_ ( .A1(_09098_ ), .A2(\RFU.rf[8][28] ), .A3(_09145_ ), .ZN(_09276_ ) );
AND4_X1 _17030_ ( .A1(_09273_ ), .A2(_09274_ ), .A3(_09275_ ), .A4(_09276_ ), .ZN(_09277_ ) );
NAND3_X1 _17031_ ( .A1(_08714_ ), .A2(\RFU.rf[14][28] ), .A3(_09148_ ), .ZN(_09278_ ) );
NAND3_X1 _17032_ ( .A1(_08727_ ), .A2(\RFU.rf[4][28] ), .A3(_09150_ ), .ZN(_09279_ ) );
NAND3_X1 _17033_ ( .A1(_08737_ ), .A2(\RFU.rf[2][28] ), .A3(_09079_ ), .ZN(_09280_ ) );
NAND3_X1 _17034_ ( .A1(_08752_ ), .A2(\RFU.rf[13][28] ), .A3(_08720_ ), .ZN(_09281_ ) );
AND4_X1 _17035_ ( .A1(_09278_ ), .A2(_09279_ ), .A3(_09280_ ), .A4(_09281_ ), .ZN(_09282_ ) );
NAND3_X1 _17036_ ( .A1(_09176_ ), .A2(_09177_ ), .A3(\RFU.rf[9][28] ), .ZN(_09283_ ) );
NAND3_X1 _17037_ ( .A1(_09179_ ), .A2(\RFU.rf[1][28] ), .A3(_09180_ ), .ZN(_09284_ ) );
NAND3_X1 _17038_ ( .A1(_09203_ ), .A2(\RFU.rf[3][28] ), .A3(_09157_ ), .ZN(_09285_ ) );
AND3_X1 _17039_ ( .A1(_09283_ ), .A2(_09284_ ), .A3(_09285_ ), .ZN(_09286_ ) );
NAND4_X1 _17040_ ( .A1(_09272_ ), .A2(_09277_ ), .A3(_09282_ ), .A4(_09286_ ), .ZN(_09287_ ) );
MUX2_X1 _17041_ ( .A(\EXU.r2_i [28] ), .B(_09287_ ), .S(_09227_ ), .Z(_00726_ ) );
NAND3_X1 _17042_ ( .A1(_08701_ ), .A2(\RFU.rf[4][1] ), .A3(_08724_ ), .ZN(_09288_ ) );
NAND3_X1 _17043_ ( .A1(_08738_ ), .A2(_08858_ ), .A3(\RFU.rf[6][1] ), .ZN(_09289_ ) );
NAND3_X1 _17044_ ( .A1(_09091_ ), .A2(\RFU.rf[7][1] ), .A3(_08731_ ), .ZN(_09290_ ) );
NAND3_X1 _17045_ ( .A1(_08858_ ), .A2(\RFU.rf[5][1] ), .A3(_08748_ ), .ZN(_09291_ ) );
AND4_X1 _17046_ ( .A1(_09288_ ), .A2(_09289_ ), .A3(_09290_ ), .A4(_09291_ ), .ZN(_09292_ ) );
NAND3_X1 _17047_ ( .A1(_08716_ ), .A2(\RFU.rf[11][1] ), .A3(_08703_ ), .ZN(_09293_ ) );
NAND3_X1 _17048_ ( .A1(_08744_ ), .A2(_08733_ ), .A3(\RFU.rf[10][1] ), .ZN(_09294_ ) );
NAND3_X1 _17049_ ( .A1(_08710_ ), .A2(_08693_ ), .A3(\RFU.rf[9][1] ), .ZN(_09295_ ) );
NAND3_X1 _17050_ ( .A1(_09098_ ), .A2(\RFU.rf[8][1] ), .A3(_09145_ ), .ZN(_09296_ ) );
AND4_X1 _17051_ ( .A1(_09293_ ), .A2(_09294_ ), .A3(_09295_ ), .A4(_09296_ ), .ZN(_09297_ ) );
NAND3_X1 _17052_ ( .A1(_08714_ ), .A2(\RFU.rf[14][1] ), .A3(_09148_ ), .ZN(_09298_ ) );
NAND3_X1 _17053_ ( .A1(_08710_ ), .A2(\RFU.rf[13][1] ), .A3(_08749_ ), .ZN(_09299_ ) );
NAND3_X1 _17054_ ( .A1(_08749_ ), .A2(\RFU.rf[12][1] ), .A3(_08723_ ), .ZN(_09300_ ) );
NAND3_X1 _17055_ ( .A1(_08749_ ), .A2(_08696_ ), .A3(\RFU.rf[15][1] ), .ZN(_09301_ ) );
AND4_X1 _17056_ ( .A1(_09298_ ), .A2(_09299_ ), .A3(_09300_ ), .A4(_09301_ ), .ZN(_09302_ ) );
NAND3_X1 _17057_ ( .A1(_08738_ ), .A2(\RFU.rf[2][1] ), .A3(_08758_ ), .ZN(_09303_ ) );
NAND3_X1 _17058_ ( .A1(_09179_ ), .A2(\RFU.rf[1][1] ), .A3(_09180_ ), .ZN(_09304_ ) );
NAND3_X1 _17059_ ( .A1(_09203_ ), .A2(\RFU.rf[3][1] ), .A3(_09157_ ), .ZN(_09305_ ) );
AND3_X1 _17060_ ( .A1(_09303_ ), .A2(_09304_ ), .A3(_09305_ ), .ZN(_09306_ ) );
NAND4_X1 _17061_ ( .A1(_09292_ ), .A2(_09297_ ), .A3(_09302_ ), .A4(_09306_ ), .ZN(_09307_ ) );
MUX2_X1 _17062_ ( .A(\EXU.r2_i [1] ), .B(_09307_ ), .S(_09227_ ), .Z(_00727_ ) );
NAND3_X1 _17063_ ( .A1(_09133_ ), .A2(\RFU.rf[11][0] ), .A3(_09185_ ), .ZN(_09308_ ) );
NAND3_X1 _17064_ ( .A1(_09089_ ), .A2(\RFU.rf[7][0] ), .A3(_09112_ ), .ZN(_09309_ ) );
NAND3_X1 _17065_ ( .A1(_08858_ ), .A2(\RFU.rf[5][0] ), .A3(_08748_ ), .ZN(_09310_ ) );
NAND3_X1 _17066_ ( .A1(_08726_ ), .A2(_09137_ ), .A3(\RFU.rf[10][0] ), .ZN(_09311_ ) );
AND4_X1 _17067_ ( .A1(_09308_ ), .A2(_09309_ ), .A3(_09310_ ), .A4(_09311_ ), .ZN(_09312_ ) );
NAND3_X1 _17068_ ( .A1(_09140_ ), .A2(\RFU.rf[12][0] ), .A3(_09117_ ), .ZN(_09313_ ) );
NAND3_X1 _17069_ ( .A1(_08744_ ), .A2(_08700_ ), .A3(\RFU.rf[6][0] ), .ZN(_09314_ ) );
NAND3_X1 _17070_ ( .A1(_09143_ ), .A2(_08696_ ), .A3(\RFU.rf[15][0] ), .ZN(_09315_ ) );
NAND3_X1 _17071_ ( .A1(_08693_ ), .A2(\RFU.rf[8][0] ), .A3(_09145_ ), .ZN(_09316_ ) );
AND4_X1 _17072_ ( .A1(_09313_ ), .A2(_09314_ ), .A3(_09315_ ), .A4(_09316_ ), .ZN(_09317_ ) );
NAND3_X1 _17073_ ( .A1(_08714_ ), .A2(\RFU.rf[14][0] ), .A3(_09148_ ), .ZN(_09318_ ) );
NAND3_X1 _17074_ ( .A1(_08727_ ), .A2(\RFU.rf[4][0] ), .A3(_09150_ ), .ZN(_09319_ ) );
NAND3_X1 _17075_ ( .A1(_08737_ ), .A2(\RFU.rf[2][0] ), .A3(_08757_ ), .ZN(_09320_ ) );
NAND3_X1 _17076_ ( .A1(_08752_ ), .A2(\RFU.rf[13][0] ), .A3(_08720_ ), .ZN(_09321_ ) );
AND4_X1 _17077_ ( .A1(_09318_ ), .A2(_09319_ ), .A3(_09320_ ), .A4(_09321_ ), .ZN(_09322_ ) );
NAND3_X1 _17078_ ( .A1(_09176_ ), .A2(_09177_ ), .A3(\RFU.rf[9][0] ), .ZN(_09323_ ) );
NAND3_X1 _17079_ ( .A1(_09179_ ), .A2(\RFU.rf[1][0] ), .A3(_09180_ ), .ZN(_09324_ ) );
NAND3_X1 _17080_ ( .A1(_09203_ ), .A2(\RFU.rf[3][0] ), .A3(_09157_ ), .ZN(_09325_ ) );
AND3_X1 _17081_ ( .A1(_09323_ ), .A2(_09324_ ), .A3(_09325_ ), .ZN(_09326_ ) );
NAND4_X1 _17082_ ( .A1(_09312_ ), .A2(_09317_ ), .A3(_09322_ ), .A4(_09326_ ), .ZN(_09327_ ) );
MUX2_X1 _17083_ ( .A(\EXU.r2_i [0] ), .B(_09327_ ), .S(_09227_ ), .Z(_00728_ ) );
NAND3_X1 _17084_ ( .A1(_09133_ ), .A2(\RFU.rf[11][27] ), .A3(_09185_ ), .ZN(_09328_ ) );
NAND3_X1 _17085_ ( .A1(_08706_ ), .A2(\RFU.rf[7][27] ), .A3(_09112_ ), .ZN(_09329_ ) );
NAND3_X1 _17086_ ( .A1(_08858_ ), .A2(\RFU.rf[5][27] ), .A3(_08748_ ), .ZN(_09330_ ) );
NAND3_X1 _17087_ ( .A1(_08726_ ), .A2(_09137_ ), .A3(\RFU.rf[10][27] ), .ZN(_09331_ ) );
AND4_X1 _17088_ ( .A1(_09328_ ), .A2(_09329_ ), .A3(_09330_ ), .A4(_09331_ ), .ZN(_09332_ ) );
NAND3_X1 _17089_ ( .A1(_09140_ ), .A2(\RFU.rf[12][27] ), .A3(_09117_ ), .ZN(_09333_ ) );
NAND3_X1 _17090_ ( .A1(_08744_ ), .A2(_08700_ ), .A3(\RFU.rf[6][27] ), .ZN(_09334_ ) );
NAND3_X1 _17091_ ( .A1(_09143_ ), .A2(_08696_ ), .A3(\RFU.rf[15][27] ), .ZN(_09335_ ) );
NAND3_X1 _17092_ ( .A1(_08693_ ), .A2(\RFU.rf[8][27] ), .A3(_09145_ ), .ZN(_09336_ ) );
AND4_X1 _17093_ ( .A1(_09333_ ), .A2(_09334_ ), .A3(_09335_ ), .A4(_09336_ ), .ZN(_09337_ ) );
NAND3_X1 _17094_ ( .A1(_08714_ ), .A2(\RFU.rf[14][27] ), .A3(_09148_ ), .ZN(_09338_ ) );
NAND3_X1 _17095_ ( .A1(_08727_ ), .A2(\RFU.rf[4][27] ), .A3(_09150_ ), .ZN(_09339_ ) );
NAND3_X1 _17096_ ( .A1(_08737_ ), .A2(\RFU.rf[2][27] ), .A3(_08757_ ), .ZN(_09340_ ) );
NAND3_X1 _17097_ ( .A1(_08752_ ), .A2(\RFU.rf[13][27] ), .A3(_08720_ ), .ZN(_09341_ ) );
AND4_X1 _17098_ ( .A1(_09338_ ), .A2(_09339_ ), .A3(_09340_ ), .A4(_09341_ ), .ZN(_09342_ ) );
NAND3_X1 _17099_ ( .A1(_09176_ ), .A2(_09177_ ), .A3(\RFU.rf[9][27] ), .ZN(_09343_ ) );
NAND3_X1 _17100_ ( .A1(_09179_ ), .A2(\RFU.rf[1][27] ), .A3(_09180_ ), .ZN(_09344_ ) );
NAND3_X1 _17101_ ( .A1(_09203_ ), .A2(\RFU.rf[3][27] ), .A3(_09157_ ), .ZN(_09345_ ) );
AND3_X1 _17102_ ( .A1(_09343_ ), .A2(_09344_ ), .A3(_09345_ ), .ZN(_09346_ ) );
NAND4_X1 _17103_ ( .A1(_09332_ ), .A2(_09337_ ), .A3(_09342_ ), .A4(_09346_ ), .ZN(_09347_ ) );
MUX2_X1 _17104_ ( .A(\EXU.r2_i [27] ), .B(_09347_ ), .S(_09227_ ), .Z(_00729_ ) );
NAND3_X1 _17105_ ( .A1(_09133_ ), .A2(\RFU.rf[11][26] ), .A3(_09185_ ), .ZN(_09348_ ) );
NAND3_X1 _17106_ ( .A1(_08706_ ), .A2(\RFU.rf[7][26] ), .A3(_08731_ ), .ZN(_09349_ ) );
NAND3_X1 _17107_ ( .A1(_08858_ ), .A2(\RFU.rf[5][26] ), .A3(_08748_ ), .ZN(_09350_ ) );
NAND3_X1 _17108_ ( .A1(_08726_ ), .A2(_09137_ ), .A3(\RFU.rf[10][26] ), .ZN(_09351_ ) );
AND4_X1 _17109_ ( .A1(_09348_ ), .A2(_09349_ ), .A3(_09350_ ), .A4(_09351_ ), .ZN(_09352_ ) );
NAND3_X1 _17110_ ( .A1(_09140_ ), .A2(\RFU.rf[12][26] ), .A3(_08742_ ), .ZN(_09353_ ) );
NAND3_X1 _17111_ ( .A1(_08744_ ), .A2(_08700_ ), .A3(\RFU.rf[6][26] ), .ZN(_09354_ ) );
NAND3_X1 _17112_ ( .A1(_09143_ ), .A2(_08696_ ), .A3(\RFU.rf[15][26] ), .ZN(_09355_ ) );
NAND3_X1 _17113_ ( .A1(_08693_ ), .A2(\RFU.rf[8][26] ), .A3(_08723_ ), .ZN(_09356_ ) );
AND4_X1 _17114_ ( .A1(_09353_ ), .A2(_09354_ ), .A3(_09355_ ), .A4(_09356_ ), .ZN(_09357_ ) );
NAND3_X1 _17115_ ( .A1(_08714_ ), .A2(\RFU.rf[14][26] ), .A3(_08730_ ), .ZN(_09358_ ) );
NAND3_X1 _17116_ ( .A1(_08727_ ), .A2(\RFU.rf[4][26] ), .A3(_09150_ ), .ZN(_09359_ ) );
NAND3_X1 _17117_ ( .A1(_08737_ ), .A2(\RFU.rf[2][26] ), .A3(_08757_ ), .ZN(_09360_ ) );
NAND3_X1 _17118_ ( .A1(_08752_ ), .A2(\RFU.rf[13][26] ), .A3(_08720_ ), .ZN(_09361_ ) );
AND4_X1 _17119_ ( .A1(_09358_ ), .A2(_09359_ ), .A3(_09360_ ), .A4(_09361_ ), .ZN(_09362_ ) );
NAND3_X1 _17120_ ( .A1(_09176_ ), .A2(_09177_ ), .A3(\RFU.rf[9][26] ), .ZN(_09363_ ) );
NAND3_X1 _17121_ ( .A1(_09179_ ), .A2(\RFU.rf[1][26] ), .A3(_09180_ ), .ZN(_09364_ ) );
NAND3_X1 _17122_ ( .A1(_09203_ ), .A2(\RFU.rf[3][26] ), .A3(_08746_ ), .ZN(_09365_ ) );
AND3_X1 _17123_ ( .A1(_09363_ ), .A2(_09364_ ), .A3(_09365_ ), .ZN(_09366_ ) );
NAND4_X1 _17124_ ( .A1(_09352_ ), .A2(_09357_ ), .A3(_09362_ ), .A4(_09366_ ), .ZN(_09367_ ) );
MUX2_X1 _17125_ ( .A(\EXU.r2_i [26] ), .B(_09367_ ), .S(_09227_ ), .Z(_00730_ ) );
NAND3_X1 _17126_ ( .A1(_08754_ ), .A2(\RFU.rf[11][25] ), .A3(_09185_ ), .ZN(_09368_ ) );
NAND3_X1 _17127_ ( .A1(_08706_ ), .A2(\RFU.rf[7][25] ), .A3(_08731_ ), .ZN(_09369_ ) );
NAND3_X1 _17128_ ( .A1(_08858_ ), .A2(\RFU.rf[5][25] ), .A3(_08748_ ), .ZN(_09370_ ) );
NAND3_X1 _17129_ ( .A1(_08726_ ), .A2(_08733_ ), .A3(\RFU.rf[10][25] ), .ZN(_09371_ ) );
AND4_X1 _17130_ ( .A1(_09368_ ), .A2(_09369_ ), .A3(_09370_ ), .A4(_09371_ ), .ZN(_09372_ ) );
NAND3_X1 _17131_ ( .A1(_08739_ ), .A2(\RFU.rf[12][25] ), .A3(_08742_ ), .ZN(_09373_ ) );
NAND3_X1 _17132_ ( .A1(_08744_ ), .A2(_08700_ ), .A3(\RFU.rf[6][25] ), .ZN(_09374_ ) );
NAND3_X1 _17133_ ( .A1(_08749_ ), .A2(_08696_ ), .A3(\RFU.rf[15][25] ), .ZN(_09375_ ) );
NAND3_X1 _17134_ ( .A1(_08693_ ), .A2(\RFU.rf[8][25] ), .A3(_08723_ ), .ZN(_09376_ ) );
AND4_X1 _17135_ ( .A1(_09373_ ), .A2(_09374_ ), .A3(_09375_ ), .A4(_09376_ ), .ZN(_09377_ ) );
NAND3_X1 _17136_ ( .A1(_08714_ ), .A2(\RFU.rf[14][25] ), .A3(_08730_ ), .ZN(_09378_ ) );
NAND3_X1 _17137_ ( .A1(_08727_ ), .A2(\RFU.rf[4][25] ), .A3(_08734_ ), .ZN(_09379_ ) );
NAND3_X1 _17138_ ( .A1(_08737_ ), .A2(\RFU.rf[2][25] ), .A3(_08757_ ), .ZN(_09380_ ) );
NAND3_X1 _17139_ ( .A1(_08752_ ), .A2(\RFU.rf[13][25] ), .A3(_08720_ ), .ZN(_09381_ ) );
AND4_X1 _17140_ ( .A1(_09378_ ), .A2(_09379_ ), .A3(_09380_ ), .A4(_09381_ ), .ZN(_09382_ ) );
NAND3_X1 _17141_ ( .A1(_09176_ ), .A2(_09177_ ), .A3(\RFU.rf[9][25] ), .ZN(_09383_ ) );
NAND3_X1 _17142_ ( .A1(_08710_ ), .A2(\RFU.rf[1][25] ), .A3(_08761_ ), .ZN(_09384_ ) );
NAND3_X1 _17143_ ( .A1(_09203_ ), .A2(\RFU.rf[3][25] ), .A3(_08746_ ), .ZN(_09385_ ) );
AND3_X1 _17144_ ( .A1(_09383_ ), .A2(_09384_ ), .A3(_09385_ ), .ZN(_09386_ ) );
NAND4_X1 _17145_ ( .A1(_09372_ ), .A2(_09377_ ), .A3(_09382_ ), .A4(_09386_ ), .ZN(_09387_ ) );
MUX2_X1 _17146_ ( .A(\EXU.r2_i [25] ), .B(_09387_ ), .S(_09227_ ), .Z(_00731_ ) );
NAND3_X1 _17147_ ( .A1(_08754_ ), .A2(\RFU.rf[11][24] ), .A3(_09185_ ), .ZN(_09388_ ) );
NAND3_X1 _17148_ ( .A1(_08706_ ), .A2(\RFU.rf[7][24] ), .A3(_08731_ ), .ZN(_09389_ ) );
NAND3_X1 _17149_ ( .A1(_08858_ ), .A2(\RFU.rf[5][24] ), .A3(_08748_ ), .ZN(_09390_ ) );
NAND3_X1 _17150_ ( .A1(_08726_ ), .A2(_08733_ ), .A3(\RFU.rf[10][24] ), .ZN(_09391_ ) );
AND4_X1 _17151_ ( .A1(_09388_ ), .A2(_09389_ ), .A3(_09390_ ), .A4(_09391_ ), .ZN(_09392_ ) );
NAND3_X1 _17152_ ( .A1(_08739_ ), .A2(\RFU.rf[12][24] ), .A3(_08742_ ), .ZN(_09393_ ) );
NAND3_X1 _17153_ ( .A1(_08744_ ), .A2(_08700_ ), .A3(\RFU.rf[6][24] ), .ZN(_09394_ ) );
NAND3_X1 _17154_ ( .A1(_08749_ ), .A2(_08696_ ), .A3(\RFU.rf[15][24] ), .ZN(_09395_ ) );
NAND3_X1 _17155_ ( .A1(_08693_ ), .A2(\RFU.rf[8][24] ), .A3(_08723_ ), .ZN(_09396_ ) );
AND4_X1 _17156_ ( .A1(_09393_ ), .A2(_09394_ ), .A3(_09395_ ), .A4(_09396_ ), .ZN(_09397_ ) );
NAND3_X1 _17157_ ( .A1(_08714_ ), .A2(\RFU.rf[14][24] ), .A3(_08730_ ), .ZN(_09398_ ) );
NAND3_X1 _17158_ ( .A1(_08727_ ), .A2(\RFU.rf[4][24] ), .A3(_08734_ ), .ZN(_09399_ ) );
NAND3_X1 _17159_ ( .A1(_08737_ ), .A2(\RFU.rf[2][24] ), .A3(_08757_ ), .ZN(_09400_ ) );
NAND3_X1 _17160_ ( .A1(_08752_ ), .A2(\RFU.rf[13][24] ), .A3(_08720_ ), .ZN(_09401_ ) );
AND4_X1 _17161_ ( .A1(_09398_ ), .A2(_09399_ ), .A3(_09400_ ), .A4(_09401_ ), .ZN(_09402_ ) );
NAND3_X1 _17162_ ( .A1(_08756_ ), .A2(_08716_ ), .A3(\RFU.rf[9][24] ), .ZN(_09403_ ) );
NAND3_X1 _17163_ ( .A1(_08710_ ), .A2(\RFU.rf[1][24] ), .A3(_08761_ ), .ZN(_09404_ ) );
NAND3_X1 _17164_ ( .A1(_08703_ ), .A2(\RFU.rf[3][24] ), .A3(_08746_ ), .ZN(_09405_ ) );
AND3_X1 _17165_ ( .A1(_09403_ ), .A2(_09404_ ), .A3(_09405_ ), .ZN(_09406_ ) );
NAND4_X1 _17166_ ( .A1(_09392_ ), .A2(_09397_ ), .A3(_09402_ ), .A4(_09406_ ), .ZN(_09407_ ) );
MUX2_X1 _17167_ ( .A(\EXU.r2_i [24] ), .B(_09407_ ), .S(_09227_ ), .Z(_00732_ ) );
NAND3_X1 _17168_ ( .A1(_08738_ ), .A2(\RFU.rf[14][23] ), .A3(_08721_ ), .ZN(_09408_ ) );
NAND3_X1 _17169_ ( .A1(_08753_ ), .A2(\RFU.rf[13][23] ), .A3(_08721_ ), .ZN(_09409_ ) );
NAND3_X1 _17170_ ( .A1(_08721_ ), .A2(\RFU.rf[12][23] ), .A3(_08724_ ), .ZN(_09410_ ) );
NAND3_X1 _17171_ ( .A1(_08721_ ), .A2(_08703_ ), .A3(\RFU.rf[15][23] ), .ZN(_09411_ ) );
AND4_X1 _17172_ ( .A1(_09408_ ), .A2(_09409_ ), .A3(_09410_ ), .A4(_09411_ ), .ZN(_09412_ ) );
NAND3_X1 _17173_ ( .A1(_08738_ ), .A2(_08694_ ), .A3(\RFU.rf[10][23] ), .ZN(_09413_ ) );
NAND3_X1 _17174_ ( .A1(_08753_ ), .A2(_08694_ ), .A3(\RFU.rf[9][23] ), .ZN(_09414_ ) );
NAND3_X1 _17175_ ( .A1(_08694_ ), .A2(\RFU.rf[8][23] ), .A3(_08724_ ), .ZN(_09415_ ) );
AND3_X1 _17176_ ( .A1(_09413_ ), .A2(_09414_ ), .A3(_09415_ ), .ZN(_09416_ ) );
NAND3_X1 _17177_ ( .A1(_08694_ ), .A2(\RFU.rf[11][23] ), .A3(_08697_ ), .ZN(_09417_ ) );
NAND3_X1 _17178_ ( .A1(_09412_ ), .A2(_09416_ ), .A3(_09417_ ), .ZN(_09418_ ) );
NAND3_X1 _17179_ ( .A1(_08701_ ), .A2(\RFU.rf[4][23] ), .A3(_08724_ ), .ZN(_09419_ ) );
NAND3_X1 _17180_ ( .A1(_08714_ ), .A2(\RFU.rf[2][23] ), .A3(_08746_ ), .ZN(_09420_ ) );
NAND3_X1 _17181_ ( .A1(_08731_ ), .A2(\RFU.rf[3][23] ), .A3(_08746_ ), .ZN(_09421_ ) );
NAND3_X1 _17182_ ( .A1(_08748_ ), .A2(\RFU.rf[1][23] ), .A3(_08746_ ), .ZN(_09422_ ) );
AND4_X1 _17183_ ( .A1(_09419_ ), .A2(_09420_ ), .A3(_09421_ ), .A4(_09422_ ), .ZN(_09423_ ) );
NAND3_X1 _17184_ ( .A1(_08701_ ), .A2(\RFU.rf[7][23] ), .A3(_08697_ ), .ZN(_09424_ ) );
NAND3_X1 _17185_ ( .A1(_08701_ ), .A2(\RFU.rf[5][23] ), .A3(_08753_ ), .ZN(_09425_ ) );
NAND3_X1 _17186_ ( .A1(_08738_ ), .A2(_08701_ ), .A3(\RFU.rf[6][23] ), .ZN(_09426_ ) );
NAND4_X1 _17187_ ( .A1(_09423_ ), .A2(_09424_ ), .A3(_09425_ ), .A4(_09426_ ), .ZN(_09427_ ) );
OAI21_X1 _17188_ ( .A(\IDU.updata ), .B1(_09418_ ), .B2(_09427_ ), .ZN(_09428_ ) );
INV_X1 _17189_ ( .A(\EXU.r2_i [23] ), .ZN(_09429_ ) );
OAI21_X1 _17190_ ( .A(_09428_ ), .B1(_09429_ ), .B2(\IDU.updata ), .ZN(_00733_ ) );
NAND3_X1 _17191_ ( .A1(_08754_ ), .A2(\RFU.rf[11][22] ), .A3(_08760_ ), .ZN(_09430_ ) );
NAND3_X1 _17192_ ( .A1(_08706_ ), .A2(\RFU.rf[7][22] ), .A3(_08731_ ), .ZN(_09431_ ) );
NAND3_X1 _17193_ ( .A1(_08858_ ), .A2(\RFU.rf[5][22] ), .A3(_08748_ ), .ZN(_09432_ ) );
NAND3_X1 _17194_ ( .A1(_08726_ ), .A2(_08733_ ), .A3(\RFU.rf[10][22] ), .ZN(_09433_ ) );
AND4_X1 _17195_ ( .A1(_09430_ ), .A2(_09431_ ), .A3(_09432_ ), .A4(_09433_ ), .ZN(_09434_ ) );
NAND3_X1 _17196_ ( .A1(_08739_ ), .A2(\RFU.rf[12][22] ), .A3(_08742_ ), .ZN(_09435_ ) );
NAND3_X1 _17197_ ( .A1(_08744_ ), .A2(_08700_ ), .A3(\RFU.rf[6][22] ), .ZN(_09436_ ) );
NAND3_X1 _17198_ ( .A1(_08749_ ), .A2(_08696_ ), .A3(\RFU.rf[15][22] ), .ZN(_09437_ ) );
NAND3_X1 _17199_ ( .A1(_08693_ ), .A2(\RFU.rf[8][22] ), .A3(_08723_ ), .ZN(_09438_ ) );
AND4_X1 _17200_ ( .A1(_09435_ ), .A2(_09436_ ), .A3(_09437_ ), .A4(_09438_ ), .ZN(_09439_ ) );
NAND3_X1 _17201_ ( .A1(_08714_ ), .A2(\RFU.rf[14][22] ), .A3(_08730_ ), .ZN(_09440_ ) );
NAND3_X1 _17202_ ( .A1(_08727_ ), .A2(\RFU.rf[4][22] ), .A3(_08734_ ), .ZN(_09441_ ) );
NAND3_X1 _17203_ ( .A1(_08737_ ), .A2(\RFU.rf[2][22] ), .A3(_08757_ ), .ZN(_09442_ ) );
NAND3_X1 _17204_ ( .A1(_08752_ ), .A2(\RFU.rf[13][22] ), .A3(_08720_ ), .ZN(_09443_ ) );
AND4_X1 _17205_ ( .A1(_09440_ ), .A2(_09441_ ), .A3(_09442_ ), .A4(_09443_ ), .ZN(_09444_ ) );
NAND3_X1 _17206_ ( .A1(_08756_ ), .A2(_08716_ ), .A3(\RFU.rf[9][22] ), .ZN(_09445_ ) );
NAND3_X1 _17207_ ( .A1(_08710_ ), .A2(\RFU.rf[1][22] ), .A3(_08761_ ), .ZN(_09446_ ) );
NAND3_X1 _17208_ ( .A1(_08703_ ), .A2(\RFU.rf[3][22] ), .A3(_08746_ ), .ZN(_09447_ ) );
AND3_X1 _17209_ ( .A1(_09445_ ), .A2(_09446_ ), .A3(_09447_ ), .ZN(_09448_ ) );
NAND4_X1 _17210_ ( .A1(_09434_ ), .A2(_09439_ ), .A3(_09444_ ), .A4(_09448_ ), .ZN(_09449_ ) );
MUX2_X1 _17211_ ( .A(\EXU.r2_i [22] ), .B(_09449_ ), .S(_07911_ ), .Z(_00734_ ) );
NOR4_X1 _17212_ ( .A1(_07927_ ), .A2(_03731_ ), .A3(_03736_ ), .A4(_03739_ ), .ZN(_09450_ ) );
NAND2_X1 _17213_ ( .A1(_09450_ ), .A2(_03929_ ), .ZN(_09451_ ) );
AND2_X1 _17214_ ( .A1(_09451_ ), .A2(\IDU.immB [3] ), .ZN(_09452_ ) );
MUX2_X1 _17215_ ( .A(\EXU.rd_i [3] ), .B(_09452_ ), .S(_07911_ ), .Z(_00735_ ) );
AND2_X1 _17216_ ( .A1(_09451_ ), .A2(\IDU.immB [2] ), .ZN(_01579_ ) );
MUX2_X1 _17217_ ( .A(\EXU.rd_i [2] ), .B(_01579_ ), .S(_07911_ ), .Z(_00736_ ) );
AND2_X1 _17218_ ( .A1(_09451_ ), .A2(\IDU.immB [1] ), .ZN(_01580_ ) );
MUX2_X1 _17219_ ( .A(\EXU.rd_i [1] ), .B(_01580_ ), .S(_07911_ ), .Z(_00737_ ) );
AND2_X1 _17220_ ( .A1(_09451_ ), .A2(\IDU.immB [11] ), .ZN(_01581_ ) );
MUX2_X1 _17221_ ( .A(\EXU.rd_i [0] ), .B(_01581_ ), .S(_07911_ ), .Z(_00738_ ) );
INV_X1 _17222_ ( .A(\IFU.state_$_NOT__A_Y ), .ZN(_01582_ ) );
NOR3_X1 _17223_ ( .A1(_07622_ ), .A2(_07660_ ), .A3(_07658_ ), .ZN(_01583_ ) );
INV_X1 _17224_ ( .A(\ICACHE.s_axi_arlen [0] ), .ZN(_01584_ ) );
NOR2_X1 _17225_ ( .A1(\ICACHE.s_axi_arlen [3] ), .A2(\ICACHE.s_axi_arlen [1] ), .ZN(_01585_ ) );
NAND3_X1 _17226_ ( .A1(_01583_ ), .A2(_01584_ ), .A3(_01585_ ), .ZN(_01586_ ) );
NAND2_X1 _17227_ ( .A1(_01585_ ), .A2(_01584_ ), .ZN(_01587_ ) );
NAND4_X1 _17228_ ( .A1(_07540_ ), .A2(io_master_rlast ), .A3(_07831_ ), .A4(_01587_ ), .ZN(_01588_ ) );
AOI21_X1 _17229_ ( .A(\ICACHE.axi_rvalid_enable ), .B1(_01586_ ), .B2(_01588_ ), .ZN(_01589_ ) );
AND4_X1 _17230_ ( .A1(_01582_ ), .A2(_01589_ ), .A3(\ICACHE.m_axi_rready ), .A4(\ICACHE.burst_counter_$_DFFE_PP__Q_E_$_ANDNOT__Y_B_$_MUX__Y_A ), .ZN(_01590_ ) );
OAI21_X1 _17231_ ( .A(_05252_ ), .B1(_01590_ ), .B2(\IDU.if_valid_i ), .ZN(_01591_ ) );
AND2_X2 _17232_ ( .A1(_05510_ ), .A2(\IDU.if_valid_i ), .ZN(_01592_ ) );
INV_X1 _17233_ ( .A(_01592_ ), .ZN(_01593_ ) );
NOR2_X1 _17234_ ( .A1(_05509_ ), .A2(_01593_ ), .ZN(_01594_ ) );
BUF_X4 _17235_ ( .A(_01594_ ), .Z(_01595_ ) );
BUF_X2 _17236_ ( .A(_01595_ ), .Z(\IFU.updata ) );
AOI21_X1 _17237_ ( .A(_01591_ ), .B1(\IFU.updata ), .B2(_01582_ ), .ZN(_00742_ ) );
BUF_X4 _17238_ ( .A(_07877_ ), .Z(_01596_ ) );
BUF_X4 _17239_ ( .A(_01592_ ), .Z(_01597_ ) );
INV_X1 _17240_ ( .A(_07659_ ), .ZN(_01598_ ) );
BUF_X4 _17241_ ( .A(_01598_ ), .Z(_01599_ ) );
BUF_X4 _17242_ ( .A(_07652_ ), .Z(_01600_ ) );
BUF_X2 _17243_ ( .A(_07646_ ), .Z(_01601_ ) );
NAND2_X1 _17244_ ( .A1(_07886_ ), .A2(\ICACHE.cache_reg[4][31] ), .ZN(_01602_ ) );
BUF_X8 _17245_ ( .A(_07548_ ), .Z(_01603_ ) );
BUF_X4 _17246_ ( .A(_01603_ ), .Z(_01604_ ) );
BUF_X8 _17247_ ( .A(_07550_ ), .Z(_01605_ ) );
BUF_X4 _17248_ ( .A(_01605_ ), .Z(_01606_ ) );
NAND3_X1 _17249_ ( .A1(_01604_ ), .A2(_01606_ ), .A3(\ICACHE.cache_reg[5][31] ), .ZN(_01607_ ) );
AOI21_X1 _17250_ ( .A(_01601_ ), .B1(_01602_ ), .B2(_01607_ ), .ZN(_01608_ ) );
BUF_X4 _17251_ ( .A(_07693_ ), .Z(_01609_ ) );
NAND2_X1 _17252_ ( .A1(_01609_ ), .A2(\ICACHE.cache_reg[6][31] ), .ZN(_01610_ ) );
BUF_X4 _17253_ ( .A(_01603_ ), .Z(_01611_ ) );
BUF_X4 _17254_ ( .A(_01605_ ), .Z(_01612_ ) );
NAND3_X1 _17255_ ( .A1(_01611_ ), .A2(_01612_ ), .A3(\ICACHE.cache_reg[7][31] ), .ZN(_01613_ ) );
AOI21_X1 _17256_ ( .A(_07841_ ), .B1(_01610_ ), .B2(_01613_ ), .ZN(_01614_ ) );
OAI21_X1 _17257_ ( .A(_01600_ ), .B1(_01608_ ), .B2(_01614_ ), .ZN(_01615_ ) );
BUF_X4 _17258_ ( .A(_07646_ ), .Z(_01616_ ) );
BUF_X4 _17259_ ( .A(_07885_ ), .Z(_01617_ ) );
NAND2_X1 _17260_ ( .A1(_01617_ ), .A2(\ICACHE.cache_reg[0][31] ), .ZN(_01618_ ) );
BUF_X4 _17261_ ( .A(_01603_ ), .Z(_01619_ ) );
BUF_X4 _17262_ ( .A(_01605_ ), .Z(_01620_ ) );
NAND3_X1 _17263_ ( .A1(_01619_ ), .A2(_01620_ ), .A3(\ICACHE.cache_reg[1][31] ), .ZN(_01621_ ) );
AOI21_X1 _17264_ ( .A(_01616_ ), .B1(_01618_ ), .B2(_01621_ ), .ZN(_01622_ ) );
BUF_X4 _17265_ ( .A(_07645_ ), .Z(_01623_ ) );
BUF_X4 _17266_ ( .A(_07693_ ), .Z(_01624_ ) );
NAND2_X1 _17267_ ( .A1(_01624_ ), .A2(\ICACHE.cache_reg[2][31] ), .ZN(_01625_ ) );
BUF_X4 _17268_ ( .A(_01603_ ), .Z(_01626_ ) );
BUF_X4 _17269_ ( .A(_01605_ ), .Z(_01627_ ) );
NAND3_X1 _17270_ ( .A1(_01626_ ), .A2(_01627_ ), .A3(\ICACHE.cache_reg[3][31] ), .ZN(_01628_ ) );
AOI21_X1 _17271_ ( .A(_01623_ ), .B1(_01625_ ), .B2(_01628_ ), .ZN(_01629_ ) );
OAI21_X1 _17272_ ( .A(_07837_ ), .B1(_01622_ ), .B2(_01629_ ), .ZN(_01630_ ) );
AOI21_X1 _17273_ ( .A(_01599_ ), .B1(_01615_ ), .B2(_01630_ ), .ZN(_01631_ ) );
NAND3_X1 _17274_ ( .A1(_01596_ ), .A2(_01597_ ), .A3(_01631_ ), .ZN(_01632_ ) );
OAI21_X1 _17275_ ( .A(_01632_ ), .B1(_03926_ ), .B2(\IFU.updata ), .ZN(_00743_ ) );
BUF_X4 _17276_ ( .A(_07652_ ), .Z(_01633_ ) );
BUF_X4 _17277_ ( .A(_07646_ ), .Z(_01634_ ) );
BUF_X4 _17278_ ( .A(_07885_ ), .Z(_01635_ ) );
NAND2_X1 _17279_ ( .A1(_01635_ ), .A2(\ICACHE.cache_reg[4][30] ), .ZN(_01636_ ) );
NAND3_X1 _17280_ ( .A1(_01604_ ), .A2(_01606_ ), .A3(\ICACHE.cache_reg[5][30] ), .ZN(_01637_ ) );
AOI21_X1 _17281_ ( .A(_01634_ ), .B1(_01636_ ), .B2(_01637_ ), .ZN(_01638_ ) );
BUF_X4 _17282_ ( .A(_07645_ ), .Z(_01639_ ) );
BUF_X4 _17283_ ( .A(_07693_ ), .Z(_01640_ ) );
NAND2_X1 _17284_ ( .A1(_01640_ ), .A2(\ICACHE.cache_reg[6][30] ), .ZN(_01641_ ) );
NAND3_X1 _17285_ ( .A1(_01611_ ), .A2(_01612_ ), .A3(\ICACHE.cache_reg[7][30] ), .ZN(_01642_ ) );
AOI21_X1 _17286_ ( .A(_01639_ ), .B1(_01641_ ), .B2(_01642_ ), .ZN(_01643_ ) );
OAI21_X1 _17287_ ( .A(_01633_ ), .B1(_01638_ ), .B2(_01643_ ), .ZN(_01644_ ) );
BUF_X4 _17288_ ( .A(_07836_ ), .Z(_01645_ ) );
BUF_X4 _17289_ ( .A(_07646_ ), .Z(_01646_ ) );
BUF_X4 _17290_ ( .A(_07885_ ), .Z(_01647_ ) );
NAND2_X1 _17291_ ( .A1(_01647_ ), .A2(\ICACHE.cache_reg[0][30] ), .ZN(_01648_ ) );
NAND3_X1 _17292_ ( .A1(_01619_ ), .A2(_01620_ ), .A3(\ICACHE.cache_reg[1][30] ), .ZN(_01649_ ) );
AOI21_X1 _17293_ ( .A(_01646_ ), .B1(_01648_ ), .B2(_01649_ ), .ZN(_01650_ ) );
BUF_X4 _17294_ ( .A(_07645_ ), .Z(_01651_ ) );
BUF_X4 _17295_ ( .A(_07693_ ), .Z(_01652_ ) );
NAND2_X1 _17296_ ( .A1(_01652_ ), .A2(\ICACHE.cache_reg[2][30] ), .ZN(_01653_ ) );
NAND3_X1 _17297_ ( .A1(_01626_ ), .A2(_01627_ ), .A3(\ICACHE.cache_reg[3][30] ), .ZN(_01654_ ) );
AOI21_X1 _17298_ ( .A(_01651_ ), .B1(_01653_ ), .B2(_01654_ ), .ZN(_01655_ ) );
OAI21_X1 _17299_ ( .A(_01645_ ), .B1(_01650_ ), .B2(_01655_ ), .ZN(_01656_ ) );
AOI21_X1 _17300_ ( .A(_01599_ ), .B1(_01644_ ), .B2(_01656_ ), .ZN(_01657_ ) );
BUF_X4 _17301_ ( .A(_01595_ ), .Z(_01658_ ) );
MUX2_X1 _17302_ ( .A(\IDU.funct7 [5] ), .B(_01657_ ), .S(_01658_ ), .Z(_00744_ ) );
BUF_X4 _17303_ ( .A(_01598_ ), .Z(_01659_ ) );
NAND2_X1 _17304_ ( .A1(_01635_ ), .A2(\ICACHE.cache_reg[4][21] ), .ZN(_01660_ ) );
BUF_X4 _17305_ ( .A(_01603_ ), .Z(_01661_ ) );
BUF_X4 _17306_ ( .A(_01605_ ), .Z(_01662_ ) );
NAND3_X1 _17307_ ( .A1(_01661_ ), .A2(_01662_ ), .A3(\ICACHE.cache_reg[5][21] ), .ZN(_01663_ ) );
AOI21_X1 _17308_ ( .A(_01634_ ), .B1(_01660_ ), .B2(_01663_ ), .ZN(_01664_ ) );
NAND2_X1 _17309_ ( .A1(_01640_ ), .A2(\ICACHE.cache_reg[6][21] ), .ZN(_01665_ ) );
BUF_X4 _17310_ ( .A(_01603_ ), .Z(_01666_ ) );
BUF_X4 _17311_ ( .A(_01605_ ), .Z(_01667_ ) );
NAND3_X1 _17312_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(\ICACHE.cache_reg[7][21] ), .ZN(_01668_ ) );
AOI21_X1 _17313_ ( .A(_01639_ ), .B1(_01665_ ), .B2(_01668_ ), .ZN(_01669_ ) );
OAI21_X1 _17314_ ( .A(_01633_ ), .B1(_01664_ ), .B2(_01669_ ), .ZN(_01670_ ) );
NAND2_X1 _17315_ ( .A1(_01647_ ), .A2(\ICACHE.cache_reg[0][21] ), .ZN(_01671_ ) );
BUF_X4 _17316_ ( .A(_01603_ ), .Z(_01672_ ) );
BUF_X4 _17317_ ( .A(_01605_ ), .Z(_01673_ ) );
NAND3_X1 _17318_ ( .A1(_01672_ ), .A2(_01673_ ), .A3(\ICACHE.cache_reg[1][21] ), .ZN(_01674_ ) );
AOI21_X1 _17319_ ( .A(_01646_ ), .B1(_01671_ ), .B2(_01674_ ), .ZN(_01675_ ) );
NAND2_X1 _17320_ ( .A1(_01652_ ), .A2(\ICACHE.cache_reg[2][21] ), .ZN(_01676_ ) );
BUF_X4 _17321_ ( .A(_07548_ ), .Z(_01677_ ) );
BUF_X4 _17322_ ( .A(_07550_ ), .Z(_01678_ ) );
NAND3_X1 _17323_ ( .A1(_01677_ ), .A2(_01678_ ), .A3(\ICACHE.cache_reg[3][21] ), .ZN(_01679_ ) );
AOI21_X1 _17324_ ( .A(_01651_ ), .B1(_01676_ ), .B2(_01679_ ), .ZN(_01680_ ) );
OAI21_X1 _17325_ ( .A(_01645_ ), .B1(_01675_ ), .B2(_01680_ ), .ZN(_01681_ ) );
AOI21_X1 _17326_ ( .A(_01659_ ), .B1(_01670_ ), .B2(_01681_ ), .ZN(_01682_ ) );
MUX2_X1 _17327_ ( .A(\IDU.immI [1] ), .B(_01682_ ), .S(_01658_ ), .Z(_00745_ ) );
NAND2_X1 _17328_ ( .A1(_01635_ ), .A2(\ICACHE.cache_reg[4][20] ), .ZN(_01683_ ) );
NAND3_X1 _17329_ ( .A1(_01661_ ), .A2(_01662_ ), .A3(\ICACHE.cache_reg[5][20] ), .ZN(_01684_ ) );
AOI21_X1 _17330_ ( .A(_01634_ ), .B1(_01683_ ), .B2(_01684_ ), .ZN(_01685_ ) );
NAND2_X1 _17331_ ( .A1(_01640_ ), .A2(\ICACHE.cache_reg[6][20] ), .ZN(_01686_ ) );
NAND3_X1 _17332_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(\ICACHE.cache_reg[7][20] ), .ZN(_01687_ ) );
AOI21_X1 _17333_ ( .A(_01639_ ), .B1(_01686_ ), .B2(_01687_ ), .ZN(_01688_ ) );
OAI21_X1 _17334_ ( .A(_01633_ ), .B1(_01685_ ), .B2(_01688_ ), .ZN(_01689_ ) );
NAND2_X1 _17335_ ( .A1(_01647_ ), .A2(\ICACHE.cache_reg[0][20] ), .ZN(_01690_ ) );
NAND3_X1 _17336_ ( .A1(_01672_ ), .A2(_01673_ ), .A3(\ICACHE.cache_reg[1][20] ), .ZN(_01691_ ) );
AOI21_X1 _17337_ ( .A(_01646_ ), .B1(_01690_ ), .B2(_01691_ ), .ZN(_01692_ ) );
NAND2_X1 _17338_ ( .A1(_01652_ ), .A2(\ICACHE.cache_reg[2][20] ), .ZN(_01693_ ) );
NAND3_X1 _17339_ ( .A1(_01677_ ), .A2(_01678_ ), .A3(\ICACHE.cache_reg[3][20] ), .ZN(_01694_ ) );
AOI21_X1 _17340_ ( .A(_01651_ ), .B1(_01693_ ), .B2(_01694_ ), .ZN(_01695_ ) );
OAI21_X1 _17341_ ( .A(_01645_ ), .B1(_01692_ ), .B2(_01695_ ), .ZN(_01696_ ) );
AOI21_X1 _17342_ ( .A(_01659_ ), .B1(_01689_ ), .B2(_01696_ ), .ZN(_01697_ ) );
MUX2_X1 _17343_ ( .A(\IDU.immI [0] ), .B(_01697_ ), .S(_01658_ ), .Z(_00746_ ) );
NAND2_X1 _17344_ ( .A1(_01635_ ), .A2(\ICACHE.cache_reg[4][19] ), .ZN(_01698_ ) );
NAND3_X1 _17345_ ( .A1(_01661_ ), .A2(_01662_ ), .A3(\ICACHE.cache_reg[5][19] ), .ZN(_01699_ ) );
AOI21_X1 _17346_ ( .A(_01634_ ), .B1(_01698_ ), .B2(_01699_ ), .ZN(_01700_ ) );
NAND2_X1 _17347_ ( .A1(_01640_ ), .A2(\ICACHE.cache_reg[6][19] ), .ZN(_01701_ ) );
NAND3_X1 _17348_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(\ICACHE.cache_reg[7][19] ), .ZN(_01702_ ) );
AOI21_X1 _17349_ ( .A(_01639_ ), .B1(_01701_ ), .B2(_01702_ ), .ZN(_01703_ ) );
OAI21_X1 _17350_ ( .A(_01633_ ), .B1(_01700_ ), .B2(_01703_ ), .ZN(_01704_ ) );
NAND2_X1 _17351_ ( .A1(_01647_ ), .A2(\ICACHE.cache_reg[0][19] ), .ZN(_01705_ ) );
NAND3_X1 _17352_ ( .A1(_01672_ ), .A2(_01673_ ), .A3(\ICACHE.cache_reg[1][19] ), .ZN(_01706_ ) );
AOI21_X1 _17353_ ( .A(_01646_ ), .B1(_01705_ ), .B2(_01706_ ), .ZN(_01707_ ) );
NAND2_X1 _17354_ ( .A1(_01652_ ), .A2(\ICACHE.cache_reg[2][19] ), .ZN(_01708_ ) );
NAND3_X1 _17355_ ( .A1(_01677_ ), .A2(_01678_ ), .A3(\ICACHE.cache_reg[3][19] ), .ZN(_01709_ ) );
AOI21_X1 _17356_ ( .A(_01651_ ), .B1(_01708_ ), .B2(_01709_ ), .ZN(_01710_ ) );
OAI21_X1 _17357_ ( .A(_01645_ ), .B1(_01707_ ), .B2(_01710_ ), .ZN(_01711_ ) );
AOI21_X1 _17358_ ( .A(_01659_ ), .B1(_01704_ ), .B2(_01711_ ), .ZN(_01712_ ) );
MUX2_X1 _17359_ ( .A(\IDU.immJ [19] ), .B(_01712_ ), .S(_01658_ ), .Z(_00747_ ) );
NAND2_X1 _17360_ ( .A1(_07886_ ), .A2(\ICACHE.cache_reg[4][18] ), .ZN(_01713_ ) );
NAND3_X1 _17361_ ( .A1(_01604_ ), .A2(_01606_ ), .A3(\ICACHE.cache_reg[5][18] ), .ZN(_01714_ ) );
AOI21_X1 _17362_ ( .A(_01601_ ), .B1(_01713_ ), .B2(_01714_ ), .ZN(_01715_ ) );
NAND2_X1 _17363_ ( .A1(_01609_ ), .A2(\ICACHE.cache_reg[6][18] ), .ZN(_01716_ ) );
NAND3_X1 _17364_ ( .A1(_01611_ ), .A2(_01612_ ), .A3(\ICACHE.cache_reg[7][18] ), .ZN(_01717_ ) );
AOI21_X1 _17365_ ( .A(_07841_ ), .B1(_01716_ ), .B2(_01717_ ), .ZN(_01718_ ) );
OAI21_X1 _17366_ ( .A(_01600_ ), .B1(_01715_ ), .B2(_01718_ ), .ZN(_01719_ ) );
NAND2_X1 _17367_ ( .A1(_01617_ ), .A2(\ICACHE.cache_reg[0][18] ), .ZN(_01720_ ) );
NAND3_X1 _17368_ ( .A1(_01619_ ), .A2(_01620_ ), .A3(\ICACHE.cache_reg[1][18] ), .ZN(_01721_ ) );
AOI21_X1 _17369_ ( .A(_01616_ ), .B1(_01720_ ), .B2(_01721_ ), .ZN(_01722_ ) );
NAND2_X1 _17370_ ( .A1(_01624_ ), .A2(\ICACHE.cache_reg[2][18] ), .ZN(_01723_ ) );
NAND3_X1 _17371_ ( .A1(_01626_ ), .A2(_01627_ ), .A3(\ICACHE.cache_reg[3][18] ), .ZN(_01724_ ) );
AOI21_X1 _17372_ ( .A(_01623_ ), .B1(_01723_ ), .B2(_01724_ ), .ZN(_01725_ ) );
OAI21_X1 _17373_ ( .A(_07837_ ), .B1(_01722_ ), .B2(_01725_ ), .ZN(_01726_ ) );
AOI21_X1 _17374_ ( .A(_01599_ ), .B1(_01719_ ), .B2(_01726_ ), .ZN(_01727_ ) );
NAND3_X1 _17375_ ( .A1(_01596_ ), .A2(_01597_ ), .A3(_01727_ ), .ZN(_01728_ ) );
OAI21_X1 _17376_ ( .A(_01728_ ), .B1(_05497_ ), .B2(\IFU.updata ), .ZN(_00748_ ) );
NAND2_X1 _17377_ ( .A1(_07886_ ), .A2(\ICACHE.cache_reg[4][17] ), .ZN(_01729_ ) );
NAND3_X1 _17378_ ( .A1(_01604_ ), .A2(_01606_ ), .A3(\ICACHE.cache_reg[5][17] ), .ZN(_01730_ ) );
AOI21_X1 _17379_ ( .A(_01601_ ), .B1(_01729_ ), .B2(_01730_ ), .ZN(_01731_ ) );
NAND2_X1 _17380_ ( .A1(_01609_ ), .A2(\ICACHE.cache_reg[6][17] ), .ZN(_01732_ ) );
NAND3_X1 _17381_ ( .A1(_01611_ ), .A2(_01612_ ), .A3(\ICACHE.cache_reg[7][17] ), .ZN(_01733_ ) );
AOI21_X1 _17382_ ( .A(_07841_ ), .B1(_01732_ ), .B2(_01733_ ), .ZN(_01734_ ) );
OAI21_X1 _17383_ ( .A(_01600_ ), .B1(_01731_ ), .B2(_01734_ ), .ZN(_01735_ ) );
NAND2_X1 _17384_ ( .A1(_01617_ ), .A2(\ICACHE.cache_reg[0][17] ), .ZN(_01736_ ) );
NAND3_X1 _17385_ ( .A1(_01619_ ), .A2(_01620_ ), .A3(\ICACHE.cache_reg[1][17] ), .ZN(_01737_ ) );
AOI21_X1 _17386_ ( .A(_01616_ ), .B1(_01736_ ), .B2(_01737_ ), .ZN(_01738_ ) );
NAND2_X1 _17387_ ( .A1(_01624_ ), .A2(\ICACHE.cache_reg[2][17] ), .ZN(_01739_ ) );
NAND3_X1 _17388_ ( .A1(_01626_ ), .A2(_01627_ ), .A3(\ICACHE.cache_reg[3][17] ), .ZN(_01740_ ) );
AOI21_X1 _17389_ ( .A(_01623_ ), .B1(_01739_ ), .B2(_01740_ ), .ZN(_01741_ ) );
OAI21_X1 _17390_ ( .A(_07837_ ), .B1(_01738_ ), .B2(_01741_ ), .ZN(_01742_ ) );
AOI21_X1 _17391_ ( .A(_01599_ ), .B1(_01735_ ), .B2(_01742_ ), .ZN(_01743_ ) );
NAND3_X1 _17392_ ( .A1(_01596_ ), .A2(_01597_ ), .A3(_01743_ ), .ZN(_01744_ ) );
OAI21_X1 _17393_ ( .A(_01744_ ), .B1(_05502_ ), .B2(\IFU.updata ), .ZN(_00749_ ) );
NAND2_X1 _17394_ ( .A1(_07886_ ), .A2(\ICACHE.cache_reg[4][16] ), .ZN(_01745_ ) );
NAND3_X1 _17395_ ( .A1(_01604_ ), .A2(_01606_ ), .A3(\ICACHE.cache_reg[5][16] ), .ZN(_01746_ ) );
AOI21_X1 _17396_ ( .A(_01601_ ), .B1(_01745_ ), .B2(_01746_ ), .ZN(_01747_ ) );
NAND2_X1 _17397_ ( .A1(_01609_ ), .A2(\ICACHE.cache_reg[6][16] ), .ZN(_01748_ ) );
NAND3_X1 _17398_ ( .A1(_01611_ ), .A2(_01612_ ), .A3(\ICACHE.cache_reg[7][16] ), .ZN(_01749_ ) );
AOI21_X1 _17399_ ( .A(_07841_ ), .B1(_01748_ ), .B2(_01749_ ), .ZN(_01750_ ) );
OAI21_X1 _17400_ ( .A(_01600_ ), .B1(_01747_ ), .B2(_01750_ ), .ZN(_01751_ ) );
NAND2_X1 _17401_ ( .A1(_01617_ ), .A2(\ICACHE.cache_reg[0][16] ), .ZN(_01752_ ) );
NAND3_X1 _17402_ ( .A1(_01619_ ), .A2(_01620_ ), .A3(\ICACHE.cache_reg[1][16] ), .ZN(_01753_ ) );
AOI21_X1 _17403_ ( .A(_01616_ ), .B1(_01752_ ), .B2(_01753_ ), .ZN(_01754_ ) );
NAND2_X1 _17404_ ( .A1(_01624_ ), .A2(\ICACHE.cache_reg[2][16] ), .ZN(_01755_ ) );
NAND3_X1 _17405_ ( .A1(_01626_ ), .A2(_01627_ ), .A3(\ICACHE.cache_reg[3][16] ), .ZN(_01756_ ) );
AOI21_X1 _17406_ ( .A(_01623_ ), .B1(_01755_ ), .B2(_01756_ ), .ZN(_01757_ ) );
OAI21_X1 _17407_ ( .A(_07837_ ), .B1(_01754_ ), .B2(_01757_ ), .ZN(_01758_ ) );
AOI21_X1 _17408_ ( .A(_01599_ ), .B1(_01751_ ), .B2(_01758_ ), .ZN(_01759_ ) );
NAND3_X1 _17409_ ( .A1(_01596_ ), .A2(_01597_ ), .A3(_01759_ ), .ZN(_01760_ ) );
OAI21_X1 _17410_ ( .A(_01760_ ), .B1(_05505_ ), .B2(\IFU.updata ), .ZN(_00750_ ) );
NAND2_X1 _17411_ ( .A1(_07886_ ), .A2(\ICACHE.cache_reg[4][15] ), .ZN(_01761_ ) );
NAND3_X1 _17412_ ( .A1(_01604_ ), .A2(_01606_ ), .A3(\ICACHE.cache_reg[5][15] ), .ZN(_01762_ ) );
AOI21_X1 _17413_ ( .A(_01601_ ), .B1(_01761_ ), .B2(_01762_ ), .ZN(_01763_ ) );
NAND2_X1 _17414_ ( .A1(_01609_ ), .A2(\ICACHE.cache_reg[6][15] ), .ZN(_01764_ ) );
NAND3_X1 _17415_ ( .A1(_01611_ ), .A2(_01612_ ), .A3(\ICACHE.cache_reg[7][15] ), .ZN(_01765_ ) );
AOI21_X1 _17416_ ( .A(_07841_ ), .B1(_01764_ ), .B2(_01765_ ), .ZN(_01766_ ) );
OAI21_X1 _17417_ ( .A(_01600_ ), .B1(_01763_ ), .B2(_01766_ ), .ZN(_01767_ ) );
NAND2_X1 _17418_ ( .A1(_01617_ ), .A2(\ICACHE.cache_reg[0][15] ), .ZN(_01768_ ) );
NAND3_X1 _17419_ ( .A1(_01619_ ), .A2(_01620_ ), .A3(\ICACHE.cache_reg[1][15] ), .ZN(_01769_ ) );
AOI21_X1 _17420_ ( .A(_01616_ ), .B1(_01768_ ), .B2(_01769_ ), .ZN(_01770_ ) );
NAND2_X1 _17421_ ( .A1(_01624_ ), .A2(\ICACHE.cache_reg[2][15] ), .ZN(_01771_ ) );
NAND3_X1 _17422_ ( .A1(_01626_ ), .A2(_01627_ ), .A3(\ICACHE.cache_reg[3][15] ), .ZN(_01772_ ) );
AOI21_X1 _17423_ ( .A(_01623_ ), .B1(_01771_ ), .B2(_01772_ ), .ZN(_01773_ ) );
OAI21_X1 _17424_ ( .A(_07837_ ), .B1(_01770_ ), .B2(_01773_ ), .ZN(_01774_ ) );
AOI21_X1 _17425_ ( .A(_01599_ ), .B1(_01767_ ), .B2(_01774_ ), .ZN(_01775_ ) );
NAND3_X1 _17426_ ( .A1(_01596_ ), .A2(_01597_ ), .A3(_01775_ ), .ZN(_01776_ ) );
OAI21_X1 _17427_ ( .A(_01776_ ), .B1(_03949_ ), .B2(\IFU.updata ), .ZN(_00751_ ) );
NAND2_X1 _17428_ ( .A1(_01635_ ), .A2(\ICACHE.cache_reg[4][14] ), .ZN(_01777_ ) );
NAND3_X1 _17429_ ( .A1(_01661_ ), .A2(_01662_ ), .A3(\ICACHE.cache_reg[5][14] ), .ZN(_01778_ ) );
AOI21_X1 _17430_ ( .A(_01634_ ), .B1(_01777_ ), .B2(_01778_ ), .ZN(_01779_ ) );
NAND2_X1 _17431_ ( .A1(_01640_ ), .A2(\ICACHE.cache_reg[6][14] ), .ZN(_01780_ ) );
NAND3_X1 _17432_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(\ICACHE.cache_reg[7][14] ), .ZN(_01781_ ) );
AOI21_X1 _17433_ ( .A(_01639_ ), .B1(_01780_ ), .B2(_01781_ ), .ZN(_01782_ ) );
OAI21_X1 _17434_ ( .A(_01633_ ), .B1(_01779_ ), .B2(_01782_ ), .ZN(_01783_ ) );
NAND2_X1 _17435_ ( .A1(_01647_ ), .A2(\ICACHE.cache_reg[0][14] ), .ZN(_01784_ ) );
NAND3_X1 _17436_ ( .A1(_01672_ ), .A2(_01673_ ), .A3(\ICACHE.cache_reg[1][14] ), .ZN(_01785_ ) );
AOI21_X1 _17437_ ( .A(_01646_ ), .B1(_01784_ ), .B2(_01785_ ), .ZN(_01786_ ) );
NAND2_X1 _17438_ ( .A1(_01652_ ), .A2(\ICACHE.cache_reg[2][14] ), .ZN(_01787_ ) );
NAND3_X1 _17439_ ( .A1(_01677_ ), .A2(_01678_ ), .A3(\ICACHE.cache_reg[3][14] ), .ZN(_01788_ ) );
AOI21_X1 _17440_ ( .A(_01651_ ), .B1(_01787_ ), .B2(_01788_ ), .ZN(_01789_ ) );
OAI21_X1 _17441_ ( .A(_01645_ ), .B1(_01786_ ), .B2(_01789_ ), .ZN(_01790_ ) );
AOI21_X1 _17442_ ( .A(_01659_ ), .B1(_01783_ ), .B2(_01790_ ), .ZN(_01791_ ) );
MUX2_X1 _17443_ ( .A(\IDU.funct3 [2] ), .B(_01791_ ), .S(_01658_ ), .Z(_00752_ ) );
NAND2_X1 _17444_ ( .A1(_01635_ ), .A2(\ICACHE.cache_reg[4][13] ), .ZN(_01792_ ) );
NAND3_X1 _17445_ ( .A1(_01661_ ), .A2(_01662_ ), .A3(\ICACHE.cache_reg[5][13] ), .ZN(_01793_ ) );
AOI21_X1 _17446_ ( .A(_01634_ ), .B1(_01792_ ), .B2(_01793_ ), .ZN(_01794_ ) );
NAND2_X1 _17447_ ( .A1(_01640_ ), .A2(\ICACHE.cache_reg[6][13] ), .ZN(_01795_ ) );
NAND3_X1 _17448_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(\ICACHE.cache_reg[7][13] ), .ZN(_01796_ ) );
AOI21_X1 _17449_ ( .A(_01639_ ), .B1(_01795_ ), .B2(_01796_ ), .ZN(_01797_ ) );
OAI21_X1 _17450_ ( .A(_01633_ ), .B1(_01794_ ), .B2(_01797_ ), .ZN(_01798_ ) );
NAND2_X1 _17451_ ( .A1(_01647_ ), .A2(\ICACHE.cache_reg[0][13] ), .ZN(_01799_ ) );
NAND3_X1 _17452_ ( .A1(_01672_ ), .A2(_01673_ ), .A3(\ICACHE.cache_reg[1][13] ), .ZN(_01800_ ) );
AOI21_X1 _17453_ ( .A(_01646_ ), .B1(_01799_ ), .B2(_01800_ ), .ZN(_01801_ ) );
NAND2_X1 _17454_ ( .A1(_01652_ ), .A2(\ICACHE.cache_reg[2][13] ), .ZN(_01802_ ) );
NAND3_X1 _17455_ ( .A1(_01677_ ), .A2(_01678_ ), .A3(\ICACHE.cache_reg[3][13] ), .ZN(_01803_ ) );
AOI21_X1 _17456_ ( .A(_01651_ ), .B1(_01802_ ), .B2(_01803_ ), .ZN(_01804_ ) );
OAI21_X1 _17457_ ( .A(_01645_ ), .B1(_01801_ ), .B2(_01804_ ), .ZN(_01805_ ) );
AOI21_X1 _17458_ ( .A(_01659_ ), .B1(_01798_ ), .B2(_01805_ ), .ZN(_01806_ ) );
MUX2_X1 _17459_ ( .A(\IDU.funct3 [1] ), .B(_01806_ ), .S(_01658_ ), .Z(_00753_ ) );
NAND2_X1 _17460_ ( .A1(_01635_ ), .A2(\ICACHE.cache_reg[4][12] ), .ZN(_01807_ ) );
NAND3_X1 _17461_ ( .A1(_01661_ ), .A2(_01662_ ), .A3(\ICACHE.cache_reg[5][12] ), .ZN(_01808_ ) );
AOI21_X1 _17462_ ( .A(_01634_ ), .B1(_01807_ ), .B2(_01808_ ), .ZN(_01809_ ) );
NAND2_X1 _17463_ ( .A1(_01640_ ), .A2(\ICACHE.cache_reg[6][12] ), .ZN(_01810_ ) );
NAND3_X1 _17464_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(\ICACHE.cache_reg[7][12] ), .ZN(_01811_ ) );
AOI21_X1 _17465_ ( .A(_01639_ ), .B1(_01810_ ), .B2(_01811_ ), .ZN(_01812_ ) );
OAI21_X1 _17466_ ( .A(_01633_ ), .B1(_01809_ ), .B2(_01812_ ), .ZN(_01813_ ) );
NAND2_X1 _17467_ ( .A1(_01647_ ), .A2(\ICACHE.cache_reg[0][12] ), .ZN(_01814_ ) );
NAND3_X1 _17468_ ( .A1(_01672_ ), .A2(_01673_ ), .A3(\ICACHE.cache_reg[1][12] ), .ZN(_01815_ ) );
AOI21_X1 _17469_ ( .A(_01646_ ), .B1(_01814_ ), .B2(_01815_ ), .ZN(_01816_ ) );
NAND2_X1 _17470_ ( .A1(_01652_ ), .A2(\ICACHE.cache_reg[2][12] ), .ZN(_01817_ ) );
NAND3_X1 _17471_ ( .A1(_01677_ ), .A2(_01678_ ), .A3(\ICACHE.cache_reg[3][12] ), .ZN(_01818_ ) );
AOI21_X1 _17472_ ( .A(_01651_ ), .B1(_01817_ ), .B2(_01818_ ), .ZN(_01819_ ) );
OAI21_X1 _17473_ ( .A(_01645_ ), .B1(_01816_ ), .B2(_01819_ ), .ZN(_01820_ ) );
AOI21_X1 _17474_ ( .A(_01659_ ), .B1(_01813_ ), .B2(_01820_ ), .ZN(_01821_ ) );
MUX2_X1 _17475_ ( .A(\IDU.funct3 [0] ), .B(_01821_ ), .S(_01658_ ), .Z(_00754_ ) );
BUF_X4 _17476_ ( .A(_07885_ ), .Z(_01822_ ) );
NAND2_X1 _17477_ ( .A1(_01822_ ), .A2(\ICACHE.cache_reg[4][29] ), .ZN(_01823_ ) );
NAND3_X1 _17478_ ( .A1(_01661_ ), .A2(_01662_ ), .A3(\ICACHE.cache_reg[5][29] ), .ZN(_01824_ ) );
AOI21_X1 _17479_ ( .A(_01634_ ), .B1(_01823_ ), .B2(_01824_ ), .ZN(_01825_ ) );
BUF_X4 _17480_ ( .A(_07693_ ), .Z(_01826_ ) );
NAND2_X1 _17481_ ( .A1(_01826_ ), .A2(\ICACHE.cache_reg[6][29] ), .ZN(_01827_ ) );
NAND3_X1 _17482_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(\ICACHE.cache_reg[7][29] ), .ZN(_01828_ ) );
AOI21_X1 _17483_ ( .A(_01639_ ), .B1(_01827_ ), .B2(_01828_ ), .ZN(_01829_ ) );
OAI21_X1 _17484_ ( .A(_01633_ ), .B1(_01825_ ), .B2(_01829_ ), .ZN(_01830_ ) );
BUF_X4 _17485_ ( .A(_07885_ ), .Z(_01831_ ) );
NAND2_X1 _17486_ ( .A1(_01831_ ), .A2(\ICACHE.cache_reg[0][29] ), .ZN(_01832_ ) );
NAND3_X1 _17487_ ( .A1(_01672_ ), .A2(_01673_ ), .A3(\ICACHE.cache_reg[1][29] ), .ZN(_01833_ ) );
AOI21_X1 _17488_ ( .A(_01646_ ), .B1(_01832_ ), .B2(_01833_ ), .ZN(_01834_ ) );
BUF_X4 _17489_ ( .A(_07693_ ), .Z(_01835_ ) );
NAND2_X1 _17490_ ( .A1(_01835_ ), .A2(\ICACHE.cache_reg[2][29] ), .ZN(_01836_ ) );
NAND3_X1 _17491_ ( .A1(_01677_ ), .A2(_01678_ ), .A3(\ICACHE.cache_reg[3][29] ), .ZN(_01837_ ) );
AOI21_X1 _17492_ ( .A(_01651_ ), .B1(_01836_ ), .B2(_01837_ ), .ZN(_01838_ ) );
OAI21_X1 _17493_ ( .A(_01645_ ), .B1(_01834_ ), .B2(_01838_ ), .ZN(_01839_ ) );
AOI21_X1 _17494_ ( .A(_01659_ ), .B1(_01830_ ), .B2(_01839_ ), .ZN(_01840_ ) );
BUF_X4 _17495_ ( .A(_01595_ ), .Z(_01841_ ) );
MUX2_X1 _17496_ ( .A(\IDU.funct7 [4] ), .B(_01840_ ), .S(_01841_ ), .Z(_00755_ ) );
NAND2_X1 _17497_ ( .A1(_01822_ ), .A2(\ICACHE.cache_reg[4][11] ), .ZN(_01842_ ) );
NAND3_X1 _17498_ ( .A1(_01661_ ), .A2(_01662_ ), .A3(\ICACHE.cache_reg[5][11] ), .ZN(_01843_ ) );
AOI21_X1 _17499_ ( .A(_01634_ ), .B1(_01842_ ), .B2(_01843_ ), .ZN(_01844_ ) );
NAND2_X1 _17500_ ( .A1(_01826_ ), .A2(\ICACHE.cache_reg[6][11] ), .ZN(_01845_ ) );
NAND3_X1 _17501_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(\ICACHE.cache_reg[7][11] ), .ZN(_01846_ ) );
AOI21_X1 _17502_ ( .A(_01639_ ), .B1(_01845_ ), .B2(_01846_ ), .ZN(_01847_ ) );
OAI21_X1 _17503_ ( .A(_01633_ ), .B1(_01844_ ), .B2(_01847_ ), .ZN(_01848_ ) );
NAND2_X1 _17504_ ( .A1(_01831_ ), .A2(\ICACHE.cache_reg[0][11] ), .ZN(_01849_ ) );
NAND3_X1 _17505_ ( .A1(_01672_ ), .A2(_01673_ ), .A3(\ICACHE.cache_reg[1][11] ), .ZN(_01850_ ) );
AOI21_X1 _17506_ ( .A(_01646_ ), .B1(_01849_ ), .B2(_01850_ ), .ZN(_01851_ ) );
NAND2_X1 _17507_ ( .A1(_01835_ ), .A2(\ICACHE.cache_reg[2][11] ), .ZN(_01852_ ) );
NAND3_X1 _17508_ ( .A1(_01677_ ), .A2(_01678_ ), .A3(\ICACHE.cache_reg[3][11] ), .ZN(_01853_ ) );
AOI21_X1 _17509_ ( .A(_01651_ ), .B1(_01852_ ), .B2(_01853_ ), .ZN(_01854_ ) );
OAI21_X1 _17510_ ( .A(_01645_ ), .B1(_01851_ ), .B2(_01854_ ), .ZN(_01855_ ) );
AOI21_X1 _17511_ ( .A(_01659_ ), .B1(_01848_ ), .B2(_01855_ ), .ZN(_01856_ ) );
MUX2_X1 _17512_ ( .A(\IDU.immB [4] ), .B(_01856_ ), .S(_01841_ ), .Z(_00756_ ) );
NAND2_X1 _17513_ ( .A1(_01822_ ), .A2(\ICACHE.cache_reg[4][10] ), .ZN(_01857_ ) );
NAND3_X1 _17514_ ( .A1(_01661_ ), .A2(_01662_ ), .A3(\ICACHE.cache_reg[5][10] ), .ZN(_01858_ ) );
AOI21_X1 _17515_ ( .A(_01634_ ), .B1(_01857_ ), .B2(_01858_ ), .ZN(_01859_ ) );
NAND2_X1 _17516_ ( .A1(_01826_ ), .A2(\ICACHE.cache_reg[6][10] ), .ZN(_01860_ ) );
NAND3_X1 _17517_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(\ICACHE.cache_reg[7][10] ), .ZN(_01861_ ) );
AOI21_X1 _17518_ ( .A(_01639_ ), .B1(_01860_ ), .B2(_01861_ ), .ZN(_01862_ ) );
OAI21_X1 _17519_ ( .A(_01633_ ), .B1(_01859_ ), .B2(_01862_ ), .ZN(_01863_ ) );
NAND2_X1 _17520_ ( .A1(_01831_ ), .A2(\ICACHE.cache_reg[0][10] ), .ZN(_01864_ ) );
NAND3_X1 _17521_ ( .A1(_01672_ ), .A2(_01673_ ), .A3(\ICACHE.cache_reg[1][10] ), .ZN(_01865_ ) );
AOI21_X1 _17522_ ( .A(_01646_ ), .B1(_01864_ ), .B2(_01865_ ), .ZN(_01866_ ) );
NAND2_X1 _17523_ ( .A1(_01835_ ), .A2(\ICACHE.cache_reg[2][10] ), .ZN(_01867_ ) );
NAND3_X1 _17524_ ( .A1(_01677_ ), .A2(_01678_ ), .A3(\ICACHE.cache_reg[3][10] ), .ZN(_01868_ ) );
AOI21_X1 _17525_ ( .A(_01651_ ), .B1(_01867_ ), .B2(_01868_ ), .ZN(_01869_ ) );
OAI21_X1 _17526_ ( .A(_01645_ ), .B1(_01866_ ), .B2(_01869_ ), .ZN(_01870_ ) );
AOI21_X1 _17527_ ( .A(_01659_ ), .B1(_01863_ ), .B2(_01870_ ), .ZN(_01871_ ) );
MUX2_X1 _17528_ ( .A(\IDU.immB [3] ), .B(_01871_ ), .S(_01841_ ), .Z(_00757_ ) );
BUF_X4 _17529_ ( .A(_07652_ ), .Z(_01872_ ) );
BUF_X4 _17530_ ( .A(_07646_ ), .Z(_01873_ ) );
NAND2_X1 _17531_ ( .A1(_01822_ ), .A2(\ICACHE.cache_reg[4][9] ), .ZN(_01874_ ) );
NAND3_X1 _17532_ ( .A1(_01661_ ), .A2(_01662_ ), .A3(\ICACHE.cache_reg[5][9] ), .ZN(_01875_ ) );
AOI21_X1 _17533_ ( .A(_01873_ ), .B1(_01874_ ), .B2(_01875_ ), .ZN(_01876_ ) );
BUF_X4 _17534_ ( .A(_07645_ ), .Z(_01877_ ) );
NAND2_X1 _17535_ ( .A1(_01826_ ), .A2(\ICACHE.cache_reg[6][9] ), .ZN(_01878_ ) );
NAND3_X1 _17536_ ( .A1(_01666_ ), .A2(_01667_ ), .A3(\ICACHE.cache_reg[7][9] ), .ZN(_01879_ ) );
AOI21_X1 _17537_ ( .A(_01877_ ), .B1(_01878_ ), .B2(_01879_ ), .ZN(_01880_ ) );
OAI21_X1 _17538_ ( .A(_01872_ ), .B1(_01876_ ), .B2(_01880_ ), .ZN(_01881_ ) );
BUF_X4 _17539_ ( .A(_07836_ ), .Z(_01882_ ) );
BUF_X4 _17540_ ( .A(_07646_ ), .Z(_01883_ ) );
NAND2_X1 _17541_ ( .A1(_01831_ ), .A2(\ICACHE.cache_reg[0][9] ), .ZN(_01884_ ) );
NAND3_X1 _17542_ ( .A1(_01672_ ), .A2(_01673_ ), .A3(\ICACHE.cache_reg[1][9] ), .ZN(_01885_ ) );
AOI21_X1 _17543_ ( .A(_01883_ ), .B1(_01884_ ), .B2(_01885_ ), .ZN(_01886_ ) );
BUF_X4 _17544_ ( .A(_07645_ ), .Z(_01887_ ) );
NAND2_X1 _17545_ ( .A1(_01835_ ), .A2(\ICACHE.cache_reg[2][9] ), .ZN(_01888_ ) );
NAND3_X1 _17546_ ( .A1(_01677_ ), .A2(_01678_ ), .A3(\ICACHE.cache_reg[3][9] ), .ZN(_01889_ ) );
AOI21_X1 _17547_ ( .A(_01887_ ), .B1(_01888_ ), .B2(_01889_ ), .ZN(_01890_ ) );
OAI21_X1 _17548_ ( .A(_01882_ ), .B1(_01886_ ), .B2(_01890_ ), .ZN(_01891_ ) );
AOI21_X1 _17549_ ( .A(_01659_ ), .B1(_01881_ ), .B2(_01891_ ), .ZN(_01892_ ) );
MUX2_X1 _17550_ ( .A(\IDU.immB [2] ), .B(_01892_ ), .S(_01841_ ), .Z(_00758_ ) );
BUF_X4 _17551_ ( .A(_01598_ ), .Z(_01893_ ) );
NAND2_X1 _17552_ ( .A1(_01822_ ), .A2(\ICACHE.cache_reg[4][8] ), .ZN(_01894_ ) );
BUF_X4 _17553_ ( .A(_01603_ ), .Z(_01895_ ) );
BUF_X4 _17554_ ( .A(_01605_ ), .Z(_01896_ ) );
NAND3_X1 _17555_ ( .A1(_01895_ ), .A2(_01896_ ), .A3(\ICACHE.cache_reg[5][8] ), .ZN(_01897_ ) );
AOI21_X1 _17556_ ( .A(_01873_ ), .B1(_01894_ ), .B2(_01897_ ), .ZN(_01898_ ) );
NAND2_X1 _17557_ ( .A1(_01826_ ), .A2(\ICACHE.cache_reg[6][8] ), .ZN(_01899_ ) );
BUF_X4 _17558_ ( .A(_01603_ ), .Z(_01900_ ) );
BUF_X4 _17559_ ( .A(_01605_ ), .Z(_01901_ ) );
NAND3_X1 _17560_ ( .A1(_01900_ ), .A2(_01901_ ), .A3(\ICACHE.cache_reg[7][8] ), .ZN(_01902_ ) );
AOI21_X1 _17561_ ( .A(_01877_ ), .B1(_01899_ ), .B2(_01902_ ), .ZN(_01903_ ) );
OAI21_X1 _17562_ ( .A(_01872_ ), .B1(_01898_ ), .B2(_01903_ ), .ZN(_01904_ ) );
NAND2_X1 _17563_ ( .A1(_01831_ ), .A2(\ICACHE.cache_reg[0][8] ), .ZN(_01905_ ) );
BUF_X4 _17564_ ( .A(_01603_ ), .Z(_01906_ ) );
BUF_X4 _17565_ ( .A(_01605_ ), .Z(_01907_ ) );
NAND3_X1 _17566_ ( .A1(_01906_ ), .A2(_01907_ ), .A3(\ICACHE.cache_reg[1][8] ), .ZN(_01908_ ) );
AOI21_X1 _17567_ ( .A(_01883_ ), .B1(_01905_ ), .B2(_01908_ ), .ZN(_01909_ ) );
NAND2_X1 _17568_ ( .A1(_01835_ ), .A2(\ICACHE.cache_reg[2][8] ), .ZN(_01910_ ) );
BUF_X4 _17569_ ( .A(_07548_ ), .Z(_01911_ ) );
BUF_X4 _17570_ ( .A(_07550_ ), .Z(_01912_ ) );
NAND3_X1 _17571_ ( .A1(_01911_ ), .A2(_01912_ ), .A3(\ICACHE.cache_reg[3][8] ), .ZN(_01913_ ) );
AOI21_X1 _17572_ ( .A(_01887_ ), .B1(_01910_ ), .B2(_01913_ ), .ZN(_01914_ ) );
OAI21_X1 _17573_ ( .A(_01882_ ), .B1(_01909_ ), .B2(_01914_ ), .ZN(_01915_ ) );
AOI21_X1 _17574_ ( .A(_01893_ ), .B1(_01904_ ), .B2(_01915_ ), .ZN(_01916_ ) );
MUX2_X1 _17575_ ( .A(\IDU.immB [1] ), .B(_01916_ ), .S(_01841_ ), .Z(_00759_ ) );
NAND2_X1 _17576_ ( .A1(_01822_ ), .A2(\ICACHE.cache_reg[4][7] ), .ZN(_01917_ ) );
NAND3_X1 _17577_ ( .A1(_01895_ ), .A2(_01896_ ), .A3(\ICACHE.cache_reg[5][7] ), .ZN(_01918_ ) );
AOI21_X1 _17578_ ( .A(_01873_ ), .B1(_01917_ ), .B2(_01918_ ), .ZN(_01919_ ) );
NAND2_X1 _17579_ ( .A1(_01826_ ), .A2(\ICACHE.cache_reg[6][7] ), .ZN(_01920_ ) );
NAND3_X1 _17580_ ( .A1(_01900_ ), .A2(_01901_ ), .A3(\ICACHE.cache_reg[7][7] ), .ZN(_01921_ ) );
AOI21_X1 _17581_ ( .A(_01877_ ), .B1(_01920_ ), .B2(_01921_ ), .ZN(_01922_ ) );
OAI21_X1 _17582_ ( .A(_01872_ ), .B1(_01919_ ), .B2(_01922_ ), .ZN(_01923_ ) );
NAND2_X1 _17583_ ( .A1(_01831_ ), .A2(\ICACHE.cache_reg[0][7] ), .ZN(_01924_ ) );
NAND3_X1 _17584_ ( .A1(_01906_ ), .A2(_01907_ ), .A3(\ICACHE.cache_reg[1][7] ), .ZN(_01925_ ) );
AOI21_X1 _17585_ ( .A(_01883_ ), .B1(_01924_ ), .B2(_01925_ ), .ZN(_01926_ ) );
NAND2_X1 _17586_ ( .A1(_01835_ ), .A2(\ICACHE.cache_reg[2][7] ), .ZN(_01927_ ) );
NAND3_X1 _17587_ ( .A1(_01911_ ), .A2(_01912_ ), .A3(\ICACHE.cache_reg[3][7] ), .ZN(_01928_ ) );
AOI21_X1 _17588_ ( .A(_01887_ ), .B1(_01927_ ), .B2(_01928_ ), .ZN(_01929_ ) );
OAI21_X1 _17589_ ( .A(_01882_ ), .B1(_01926_ ), .B2(_01929_ ), .ZN(_01930_ ) );
AOI21_X1 _17590_ ( .A(_01893_ ), .B1(_01923_ ), .B2(_01930_ ), .ZN(_01931_ ) );
MUX2_X1 _17591_ ( .A(\IDU.immB [11] ), .B(_01931_ ), .S(_01841_ ), .Z(_00760_ ) );
NAND2_X1 _17592_ ( .A1(_07886_ ), .A2(\ICACHE.cache_reg[4][6] ), .ZN(_01932_ ) );
NAND3_X1 _17593_ ( .A1(_01604_ ), .A2(_01606_ ), .A3(\ICACHE.cache_reg[5][6] ), .ZN(_01933_ ) );
AOI21_X1 _17594_ ( .A(_01601_ ), .B1(_01932_ ), .B2(_01933_ ), .ZN(_01934_ ) );
NAND2_X1 _17595_ ( .A1(_01609_ ), .A2(\ICACHE.cache_reg[6][6] ), .ZN(_01935_ ) );
NAND3_X1 _17596_ ( .A1(_01611_ ), .A2(_01612_ ), .A3(\ICACHE.cache_reg[7][6] ), .ZN(_01936_ ) );
AOI21_X1 _17597_ ( .A(_07841_ ), .B1(_01935_ ), .B2(_01936_ ), .ZN(_01937_ ) );
OAI21_X1 _17598_ ( .A(_01600_ ), .B1(_01934_ ), .B2(_01937_ ), .ZN(_01938_ ) );
NAND2_X1 _17599_ ( .A1(_01617_ ), .A2(\ICACHE.cache_reg[0][6] ), .ZN(_01939_ ) );
NAND3_X1 _17600_ ( .A1(_01619_ ), .A2(_01620_ ), .A3(\ICACHE.cache_reg[1][6] ), .ZN(_01940_ ) );
AOI21_X1 _17601_ ( .A(_01616_ ), .B1(_01939_ ), .B2(_01940_ ), .ZN(_01941_ ) );
NAND2_X1 _17602_ ( .A1(_01624_ ), .A2(\ICACHE.cache_reg[2][6] ), .ZN(_01942_ ) );
NAND3_X1 _17603_ ( .A1(_01626_ ), .A2(_01627_ ), .A3(\ICACHE.cache_reg[3][6] ), .ZN(_01943_ ) );
AOI21_X1 _17604_ ( .A(_01623_ ), .B1(_01942_ ), .B2(_01943_ ), .ZN(_01944_ ) );
OAI21_X1 _17605_ ( .A(_07837_ ), .B1(_01941_ ), .B2(_01944_ ), .ZN(_01945_ ) );
AOI21_X1 _17606_ ( .A(_01599_ ), .B1(_01938_ ), .B2(_01945_ ), .ZN(_01946_ ) );
NAND3_X1 _17607_ ( .A1(_01596_ ), .A2(_01597_ ), .A3(_01946_ ), .ZN(_01947_ ) );
OAI21_X1 _17608_ ( .A(_01947_ ), .B1(_03732_ ), .B2(\IFU.updata ), .ZN(_00761_ ) );
NAND2_X1 _17609_ ( .A1(_01635_ ), .A2(\ICACHE.cache_reg[4][5] ), .ZN(_01948_ ) );
NAND3_X1 _17610_ ( .A1(_01604_ ), .A2(_01606_ ), .A3(\ICACHE.cache_reg[5][5] ), .ZN(_01949_ ) );
AOI21_X1 _17611_ ( .A(_01601_ ), .B1(_01948_ ), .B2(_01949_ ), .ZN(_01950_ ) );
NAND2_X1 _17612_ ( .A1(_01640_ ), .A2(\ICACHE.cache_reg[6][5] ), .ZN(_01951_ ) );
NAND3_X1 _17613_ ( .A1(_01611_ ), .A2(_01612_ ), .A3(\ICACHE.cache_reg[7][5] ), .ZN(_01952_ ) );
AOI21_X1 _17614_ ( .A(_07841_ ), .B1(_01951_ ), .B2(_01952_ ), .ZN(_01953_ ) );
OAI21_X1 _17615_ ( .A(_01600_ ), .B1(_01950_ ), .B2(_01953_ ), .ZN(_01954_ ) );
NAND2_X1 _17616_ ( .A1(_01647_ ), .A2(\ICACHE.cache_reg[0][5] ), .ZN(_01955_ ) );
NAND3_X1 _17617_ ( .A1(_01619_ ), .A2(_01620_ ), .A3(\ICACHE.cache_reg[1][5] ), .ZN(_01956_ ) );
AOI21_X1 _17618_ ( .A(_01616_ ), .B1(_01955_ ), .B2(_01956_ ), .ZN(_01957_ ) );
NAND2_X1 _17619_ ( .A1(_01652_ ), .A2(\ICACHE.cache_reg[2][5] ), .ZN(_01958_ ) );
NAND3_X1 _17620_ ( .A1(_01626_ ), .A2(_01627_ ), .A3(\ICACHE.cache_reg[3][5] ), .ZN(_01959_ ) );
AOI21_X1 _17621_ ( .A(_01623_ ), .B1(_01958_ ), .B2(_01959_ ), .ZN(_01960_ ) );
OAI21_X1 _17622_ ( .A(_07837_ ), .B1(_01957_ ), .B2(_01960_ ), .ZN(_01961_ ) );
AOI21_X1 _17623_ ( .A(_01599_ ), .B1(_01954_ ), .B2(_01961_ ), .ZN(_01962_ ) );
NAND3_X1 _17624_ ( .A1(_01596_ ), .A2(_01597_ ), .A3(_01962_ ), .ZN(_01963_ ) );
OAI21_X1 _17625_ ( .A(_01963_ ), .B1(_03733_ ), .B2(\IFU.updata ), .ZN(_00762_ ) );
NAND2_X1 _17626_ ( .A1(_01635_ ), .A2(\ICACHE.cache_reg[4][4] ), .ZN(_01964_ ) );
NAND3_X1 _17627_ ( .A1(_01604_ ), .A2(_01606_ ), .A3(\ICACHE.cache_reg[5][4] ), .ZN(_01965_ ) );
AOI21_X1 _17628_ ( .A(_01601_ ), .B1(_01964_ ), .B2(_01965_ ), .ZN(_01966_ ) );
NAND2_X1 _17629_ ( .A1(_01640_ ), .A2(\ICACHE.cache_reg[6][4] ), .ZN(_01967_ ) );
NAND3_X1 _17630_ ( .A1(_01611_ ), .A2(_01612_ ), .A3(\ICACHE.cache_reg[7][4] ), .ZN(_01968_ ) );
AOI21_X1 _17631_ ( .A(_07841_ ), .B1(_01967_ ), .B2(_01968_ ), .ZN(_01969_ ) );
OAI21_X1 _17632_ ( .A(_01600_ ), .B1(_01966_ ), .B2(_01969_ ), .ZN(_01970_ ) );
NAND2_X1 _17633_ ( .A1(_01647_ ), .A2(\ICACHE.cache_reg[0][4] ), .ZN(_01971_ ) );
NAND3_X1 _17634_ ( .A1(_01619_ ), .A2(_01620_ ), .A3(\ICACHE.cache_reg[1][4] ), .ZN(_01972_ ) );
AOI21_X1 _17635_ ( .A(_01616_ ), .B1(_01971_ ), .B2(_01972_ ), .ZN(_01973_ ) );
NAND2_X1 _17636_ ( .A1(_01652_ ), .A2(\ICACHE.cache_reg[2][4] ), .ZN(_01974_ ) );
NAND3_X1 _17637_ ( .A1(_01626_ ), .A2(_01627_ ), .A3(\ICACHE.cache_reg[3][4] ), .ZN(_01975_ ) );
AOI21_X1 _17638_ ( .A(_01623_ ), .B1(_01974_ ), .B2(_01975_ ), .ZN(_01976_ ) );
OAI21_X1 _17639_ ( .A(_07837_ ), .B1(_01973_ ), .B2(_01976_ ), .ZN(_01977_ ) );
AOI21_X1 _17640_ ( .A(_01599_ ), .B1(_01970_ ), .B2(_01977_ ), .ZN(_01978_ ) );
NAND3_X1 _17641_ ( .A1(_01596_ ), .A2(_01597_ ), .A3(_01978_ ), .ZN(_01979_ ) );
OAI21_X1 _17642_ ( .A(_01979_ ), .B1(_03722_ ), .B2(_01658_ ), .ZN(_00763_ ) );
NAND2_X1 _17643_ ( .A1(_01822_ ), .A2(\ICACHE.cache_reg[4][3] ), .ZN(_01980_ ) );
NAND3_X1 _17644_ ( .A1(_01895_ ), .A2(_01896_ ), .A3(\ICACHE.cache_reg[5][3] ), .ZN(_01981_ ) );
AOI21_X1 _17645_ ( .A(_01873_ ), .B1(_01980_ ), .B2(_01981_ ), .ZN(_01982_ ) );
NAND2_X1 _17646_ ( .A1(_01826_ ), .A2(\ICACHE.cache_reg[6][3] ), .ZN(_01983_ ) );
NAND3_X1 _17647_ ( .A1(_01900_ ), .A2(_01901_ ), .A3(\ICACHE.cache_reg[7][3] ), .ZN(_01984_ ) );
AOI21_X1 _17648_ ( .A(_01877_ ), .B1(_01983_ ), .B2(_01984_ ), .ZN(_01985_ ) );
OAI21_X1 _17649_ ( .A(_01872_ ), .B1(_01982_ ), .B2(_01985_ ), .ZN(_01986_ ) );
NAND2_X1 _17650_ ( .A1(_01831_ ), .A2(\ICACHE.cache_reg[0][3] ), .ZN(_01987_ ) );
NAND3_X1 _17651_ ( .A1(_01906_ ), .A2(_01907_ ), .A3(\ICACHE.cache_reg[1][3] ), .ZN(_01988_ ) );
AOI21_X1 _17652_ ( .A(_01883_ ), .B1(_01987_ ), .B2(_01988_ ), .ZN(_01989_ ) );
NAND2_X1 _17653_ ( .A1(_01835_ ), .A2(\ICACHE.cache_reg[2][3] ), .ZN(_01990_ ) );
NAND3_X1 _17654_ ( .A1(_01911_ ), .A2(_01912_ ), .A3(\ICACHE.cache_reg[3][3] ), .ZN(_01991_ ) );
AOI21_X1 _17655_ ( .A(_01887_ ), .B1(_01990_ ), .B2(_01991_ ), .ZN(_01992_ ) );
OAI21_X1 _17656_ ( .A(_01882_ ), .B1(_01989_ ), .B2(_01992_ ), .ZN(_01993_ ) );
AOI21_X1 _17657_ ( .A(_01893_ ), .B1(_01986_ ), .B2(_01993_ ), .ZN(_01994_ ) );
MUX2_X1 _17658_ ( .A(\IDU.inst_i [3] ), .B(_01994_ ), .S(_01841_ ), .Z(_00764_ ) );
NAND2_X1 _17659_ ( .A1(_01635_ ), .A2(\ICACHE.cache_reg[4][2] ), .ZN(_01995_ ) );
NAND3_X1 _17660_ ( .A1(_01604_ ), .A2(_01606_ ), .A3(\ICACHE.cache_reg[5][2] ), .ZN(_01996_ ) );
AOI21_X1 _17661_ ( .A(_01601_ ), .B1(_01995_ ), .B2(_01996_ ), .ZN(_01997_ ) );
NAND2_X1 _17662_ ( .A1(_01640_ ), .A2(\ICACHE.cache_reg[6][2] ), .ZN(_01998_ ) );
NAND3_X1 _17663_ ( .A1(_01611_ ), .A2(_01612_ ), .A3(\ICACHE.cache_reg[7][2] ), .ZN(_01999_ ) );
AOI21_X1 _17664_ ( .A(_07841_ ), .B1(_01998_ ), .B2(_01999_ ), .ZN(_02000_ ) );
OAI21_X1 _17665_ ( .A(_01600_ ), .B1(_01997_ ), .B2(_02000_ ), .ZN(_02001_ ) );
NAND2_X1 _17666_ ( .A1(_01647_ ), .A2(\ICACHE.cache_reg[0][2] ), .ZN(_02002_ ) );
NAND3_X1 _17667_ ( .A1(_01619_ ), .A2(_01620_ ), .A3(\ICACHE.cache_reg[1][2] ), .ZN(_02003_ ) );
AOI21_X1 _17668_ ( .A(_01616_ ), .B1(_02002_ ), .B2(_02003_ ), .ZN(_02004_ ) );
NAND2_X1 _17669_ ( .A1(_01652_ ), .A2(\ICACHE.cache_reg[2][2] ), .ZN(_02005_ ) );
NAND3_X1 _17670_ ( .A1(_01626_ ), .A2(_01627_ ), .A3(\ICACHE.cache_reg[3][2] ), .ZN(_02006_ ) );
AOI21_X1 _17671_ ( .A(_01623_ ), .B1(_02005_ ), .B2(_02006_ ), .ZN(_02007_ ) );
OAI21_X1 _17672_ ( .A(_07837_ ), .B1(_02004_ ), .B2(_02007_ ), .ZN(_02008_ ) );
AOI21_X1 _17673_ ( .A(_01599_ ), .B1(_02001_ ), .B2(_02008_ ), .ZN(_02009_ ) );
NAND3_X1 _17674_ ( .A1(_01596_ ), .A2(_01597_ ), .A3(_02009_ ), .ZN(_02010_ ) );
OAI21_X1 _17675_ ( .A(_02010_ ), .B1(_03729_ ), .B2(_01658_ ), .ZN(_00765_ ) );
NAND2_X1 _17676_ ( .A1(_01822_ ), .A2(\ICACHE.cache_reg[4][28] ), .ZN(_02011_ ) );
NAND3_X1 _17677_ ( .A1(_01895_ ), .A2(_01896_ ), .A3(\ICACHE.cache_reg[5][28] ), .ZN(_02012_ ) );
AOI21_X1 _17678_ ( .A(_01873_ ), .B1(_02011_ ), .B2(_02012_ ), .ZN(_02013_ ) );
NAND2_X1 _17679_ ( .A1(_01826_ ), .A2(\ICACHE.cache_reg[6][28] ), .ZN(_02014_ ) );
NAND3_X1 _17680_ ( .A1(_01900_ ), .A2(_01901_ ), .A3(\ICACHE.cache_reg[7][28] ), .ZN(_02015_ ) );
AOI21_X1 _17681_ ( .A(_01877_ ), .B1(_02014_ ), .B2(_02015_ ), .ZN(_02016_ ) );
OAI21_X1 _17682_ ( .A(_01872_ ), .B1(_02013_ ), .B2(_02016_ ), .ZN(_02017_ ) );
NAND2_X1 _17683_ ( .A1(_01831_ ), .A2(\ICACHE.cache_reg[0][28] ), .ZN(_02018_ ) );
NAND3_X1 _17684_ ( .A1(_01906_ ), .A2(_01907_ ), .A3(\ICACHE.cache_reg[1][28] ), .ZN(_02019_ ) );
AOI21_X1 _17685_ ( .A(_01883_ ), .B1(_02018_ ), .B2(_02019_ ), .ZN(_02020_ ) );
NAND2_X1 _17686_ ( .A1(_01835_ ), .A2(\ICACHE.cache_reg[2][28] ), .ZN(_02021_ ) );
NAND3_X1 _17687_ ( .A1(_01911_ ), .A2(_01912_ ), .A3(\ICACHE.cache_reg[3][28] ), .ZN(_02022_ ) );
AOI21_X1 _17688_ ( .A(_01887_ ), .B1(_02021_ ), .B2(_02022_ ), .ZN(_02023_ ) );
OAI21_X1 _17689_ ( .A(_01882_ ), .B1(_02020_ ), .B2(_02023_ ), .ZN(_02024_ ) );
AOI21_X1 _17690_ ( .A(_01893_ ), .B1(_02017_ ), .B2(_02024_ ), .ZN(_02025_ ) );
MUX2_X1 _17691_ ( .A(\IDU.funct7 [3] ), .B(_02025_ ), .S(_01841_ ), .Z(_00766_ ) );
NAND2_X1 _17692_ ( .A1(_01822_ ), .A2(\ICACHE.cache_reg[4][27] ), .ZN(_02026_ ) );
NAND3_X1 _17693_ ( .A1(_01895_ ), .A2(_01896_ ), .A3(\ICACHE.cache_reg[5][27] ), .ZN(_02027_ ) );
AOI21_X1 _17694_ ( .A(_01873_ ), .B1(_02026_ ), .B2(_02027_ ), .ZN(_02028_ ) );
NAND2_X1 _17695_ ( .A1(_01826_ ), .A2(\ICACHE.cache_reg[6][27] ), .ZN(_02029_ ) );
NAND3_X1 _17696_ ( .A1(_01900_ ), .A2(_01901_ ), .A3(\ICACHE.cache_reg[7][27] ), .ZN(_02030_ ) );
AOI21_X1 _17697_ ( .A(_01877_ ), .B1(_02029_ ), .B2(_02030_ ), .ZN(_02031_ ) );
OAI21_X1 _17698_ ( .A(_01872_ ), .B1(_02028_ ), .B2(_02031_ ), .ZN(_02032_ ) );
NAND2_X1 _17699_ ( .A1(_01831_ ), .A2(\ICACHE.cache_reg[0][27] ), .ZN(_02033_ ) );
NAND3_X1 _17700_ ( .A1(_01906_ ), .A2(_01907_ ), .A3(\ICACHE.cache_reg[1][27] ), .ZN(_02034_ ) );
AOI21_X1 _17701_ ( .A(_01883_ ), .B1(_02033_ ), .B2(_02034_ ), .ZN(_02035_ ) );
NAND2_X1 _17702_ ( .A1(_01835_ ), .A2(\ICACHE.cache_reg[2][27] ), .ZN(_02036_ ) );
NAND3_X1 _17703_ ( .A1(_01911_ ), .A2(_01912_ ), .A3(\ICACHE.cache_reg[3][27] ), .ZN(_02037_ ) );
AOI21_X1 _17704_ ( .A(_01887_ ), .B1(_02036_ ), .B2(_02037_ ), .ZN(_02038_ ) );
OAI21_X1 _17705_ ( .A(_01882_ ), .B1(_02035_ ), .B2(_02038_ ), .ZN(_02039_ ) );
AOI21_X1 _17706_ ( .A(_01893_ ), .B1(_02032_ ), .B2(_02039_ ), .ZN(_02040_ ) );
MUX2_X1 _17707_ ( .A(\IDU.funct7 [2] ), .B(_02040_ ), .S(_01841_ ), .Z(_00767_ ) );
NAND2_X1 _17708_ ( .A1(_01822_ ), .A2(\ICACHE.cache_reg[4][26] ), .ZN(_02041_ ) );
NAND3_X1 _17709_ ( .A1(_01895_ ), .A2(_01896_ ), .A3(\ICACHE.cache_reg[5][26] ), .ZN(_02042_ ) );
AOI21_X1 _17710_ ( .A(_01873_ ), .B1(_02041_ ), .B2(_02042_ ), .ZN(_02043_ ) );
NAND2_X1 _17711_ ( .A1(_01826_ ), .A2(\ICACHE.cache_reg[6][26] ), .ZN(_02044_ ) );
NAND3_X1 _17712_ ( .A1(_01900_ ), .A2(_01901_ ), .A3(\ICACHE.cache_reg[7][26] ), .ZN(_02045_ ) );
AOI21_X1 _17713_ ( .A(_01877_ ), .B1(_02044_ ), .B2(_02045_ ), .ZN(_02046_ ) );
OAI21_X1 _17714_ ( .A(_01872_ ), .B1(_02043_ ), .B2(_02046_ ), .ZN(_02047_ ) );
NAND2_X1 _17715_ ( .A1(_01831_ ), .A2(\ICACHE.cache_reg[0][26] ), .ZN(_02048_ ) );
NAND3_X1 _17716_ ( .A1(_01906_ ), .A2(_01907_ ), .A3(\ICACHE.cache_reg[1][26] ), .ZN(_02049_ ) );
AOI21_X1 _17717_ ( .A(_01883_ ), .B1(_02048_ ), .B2(_02049_ ), .ZN(_02050_ ) );
NAND2_X1 _17718_ ( .A1(_01835_ ), .A2(\ICACHE.cache_reg[2][26] ), .ZN(_02051_ ) );
NAND3_X1 _17719_ ( .A1(_01911_ ), .A2(_01912_ ), .A3(\ICACHE.cache_reg[3][26] ), .ZN(_02052_ ) );
AOI21_X1 _17720_ ( .A(_01887_ ), .B1(_02051_ ), .B2(_02052_ ), .ZN(_02053_ ) );
OAI21_X1 _17721_ ( .A(_01882_ ), .B1(_02050_ ), .B2(_02053_ ), .ZN(_02054_ ) );
AOI21_X1 _17722_ ( .A(_01893_ ), .B1(_02047_ ), .B2(_02054_ ), .ZN(_02055_ ) );
MUX2_X1 _17723_ ( .A(\IDU.funct7 [1] ), .B(_02055_ ), .S(_01841_ ), .Z(_00768_ ) );
NAND2_X1 _17724_ ( .A1(_01617_ ), .A2(\ICACHE.cache_reg[4][25] ), .ZN(_02056_ ) );
NAND3_X1 _17725_ ( .A1(_01895_ ), .A2(_01896_ ), .A3(\ICACHE.cache_reg[5][25] ), .ZN(_02057_ ) );
AOI21_X1 _17726_ ( .A(_01873_ ), .B1(_02056_ ), .B2(_02057_ ), .ZN(_02058_ ) );
NAND2_X1 _17727_ ( .A1(_01624_ ), .A2(\ICACHE.cache_reg[6][25] ), .ZN(_02059_ ) );
NAND3_X1 _17728_ ( .A1(_01900_ ), .A2(_01901_ ), .A3(\ICACHE.cache_reg[7][25] ), .ZN(_02060_ ) );
AOI21_X1 _17729_ ( .A(_01877_ ), .B1(_02059_ ), .B2(_02060_ ), .ZN(_02061_ ) );
OAI21_X1 _17730_ ( .A(_01872_ ), .B1(_02058_ ), .B2(_02061_ ), .ZN(_02062_ ) );
NAND2_X1 _17731_ ( .A1(_01609_ ), .A2(\ICACHE.cache_reg[0][25] ), .ZN(_02063_ ) );
NAND3_X1 _17732_ ( .A1(_01906_ ), .A2(_01907_ ), .A3(\ICACHE.cache_reg[1][25] ), .ZN(_02064_ ) );
AOI21_X1 _17733_ ( .A(_01883_ ), .B1(_02063_ ), .B2(_02064_ ), .ZN(_02065_ ) );
NAND2_X1 _17734_ ( .A1(_07885_ ), .A2(\ICACHE.cache_reg[2][25] ), .ZN(_02066_ ) );
NAND3_X1 _17735_ ( .A1(_01911_ ), .A2(_01912_ ), .A3(\ICACHE.cache_reg[3][25] ), .ZN(_02067_ ) );
AOI21_X1 _17736_ ( .A(_01887_ ), .B1(_02066_ ), .B2(_02067_ ), .ZN(_02068_ ) );
OAI21_X1 _17737_ ( .A(_01882_ ), .B1(_02065_ ), .B2(_02068_ ), .ZN(_02069_ ) );
AOI21_X1 _17738_ ( .A(_01893_ ), .B1(_02062_ ), .B2(_02069_ ), .ZN(_02070_ ) );
BUF_X4 _17739_ ( .A(_01595_ ), .Z(_02071_ ) );
MUX2_X1 _17740_ ( .A(\IDU.funct7 [0] ), .B(_02070_ ), .S(_02071_ ), .Z(_00769_ ) );
NAND2_X1 _17741_ ( .A1(_01617_ ), .A2(\ICACHE.cache_reg[4][24] ), .ZN(_02072_ ) );
NAND3_X1 _17742_ ( .A1(_01895_ ), .A2(_01896_ ), .A3(\ICACHE.cache_reg[5][24] ), .ZN(_02073_ ) );
AOI21_X1 _17743_ ( .A(_01873_ ), .B1(_02072_ ), .B2(_02073_ ), .ZN(_02074_ ) );
NAND2_X1 _17744_ ( .A1(_01624_ ), .A2(\ICACHE.cache_reg[6][24] ), .ZN(_02075_ ) );
NAND3_X1 _17745_ ( .A1(_01900_ ), .A2(_01901_ ), .A3(\ICACHE.cache_reg[7][24] ), .ZN(_02076_ ) );
AOI21_X1 _17746_ ( .A(_01877_ ), .B1(_02075_ ), .B2(_02076_ ), .ZN(_02077_ ) );
OAI21_X1 _17747_ ( .A(_01872_ ), .B1(_02074_ ), .B2(_02077_ ), .ZN(_02078_ ) );
NAND2_X1 _17748_ ( .A1(_01609_ ), .A2(\ICACHE.cache_reg[0][24] ), .ZN(_02079_ ) );
NAND3_X1 _17749_ ( .A1(_01906_ ), .A2(_01907_ ), .A3(\ICACHE.cache_reg[1][24] ), .ZN(_02080_ ) );
AOI21_X1 _17750_ ( .A(_01883_ ), .B1(_02079_ ), .B2(_02080_ ), .ZN(_02081_ ) );
NAND2_X1 _17751_ ( .A1(_07885_ ), .A2(\ICACHE.cache_reg[2][24] ), .ZN(_02082_ ) );
NAND3_X1 _17752_ ( .A1(_01911_ ), .A2(_01912_ ), .A3(\ICACHE.cache_reg[3][24] ), .ZN(_02083_ ) );
AOI21_X1 _17753_ ( .A(_01887_ ), .B1(_02082_ ), .B2(_02083_ ), .ZN(_02084_ ) );
OAI21_X1 _17754_ ( .A(_01882_ ), .B1(_02081_ ), .B2(_02084_ ), .ZN(_02085_ ) );
AOI21_X1 _17755_ ( .A(_01893_ ), .B1(_02078_ ), .B2(_02085_ ), .ZN(_02086_ ) );
MUX2_X1 _17756_ ( .A(\IDU.immI [4] ), .B(_02086_ ), .S(_02071_ ), .Z(_00770_ ) );
NAND2_X1 _17757_ ( .A1(_01617_ ), .A2(\ICACHE.cache_reg[4][23] ), .ZN(_02087_ ) );
NAND3_X1 _17758_ ( .A1(_01895_ ), .A2(_01896_ ), .A3(\ICACHE.cache_reg[5][23] ), .ZN(_02088_ ) );
AOI21_X1 _17759_ ( .A(_01873_ ), .B1(_02087_ ), .B2(_02088_ ), .ZN(_02089_ ) );
NAND2_X1 _17760_ ( .A1(_01624_ ), .A2(\ICACHE.cache_reg[6][23] ), .ZN(_02090_ ) );
NAND3_X1 _17761_ ( .A1(_01900_ ), .A2(_01901_ ), .A3(\ICACHE.cache_reg[7][23] ), .ZN(_02091_ ) );
AOI21_X1 _17762_ ( .A(_01877_ ), .B1(_02090_ ), .B2(_02091_ ), .ZN(_02092_ ) );
OAI21_X1 _17763_ ( .A(_01872_ ), .B1(_02089_ ), .B2(_02092_ ), .ZN(_02093_ ) );
NAND2_X1 _17764_ ( .A1(_01609_ ), .A2(\ICACHE.cache_reg[0][23] ), .ZN(_02094_ ) );
NAND3_X1 _17765_ ( .A1(_01906_ ), .A2(_01907_ ), .A3(\ICACHE.cache_reg[1][23] ), .ZN(_02095_ ) );
AOI21_X1 _17766_ ( .A(_01883_ ), .B1(_02094_ ), .B2(_02095_ ), .ZN(_02096_ ) );
NAND2_X1 _17767_ ( .A1(_07885_ ), .A2(\ICACHE.cache_reg[2][23] ), .ZN(_02097_ ) );
NAND3_X1 _17768_ ( .A1(_01911_ ), .A2(_01912_ ), .A3(\ICACHE.cache_reg[3][23] ), .ZN(_02098_ ) );
AOI21_X1 _17769_ ( .A(_01887_ ), .B1(_02097_ ), .B2(_02098_ ), .ZN(_02099_ ) );
OAI21_X1 _17770_ ( .A(_01882_ ), .B1(_02096_ ), .B2(_02099_ ), .ZN(_02100_ ) );
AOI21_X1 _17771_ ( .A(_01893_ ), .B1(_02093_ ), .B2(_02100_ ), .ZN(_02101_ ) );
MUX2_X1 _17772_ ( .A(\IDU.immI [3] ), .B(_02101_ ), .S(_02071_ ), .Z(_00771_ ) );
NAND2_X1 _17773_ ( .A1(_01617_ ), .A2(\ICACHE.cache_reg[4][22] ), .ZN(_02102_ ) );
NAND3_X1 _17774_ ( .A1(_01895_ ), .A2(_01896_ ), .A3(\ICACHE.cache_reg[5][22] ), .ZN(_02103_ ) );
AOI21_X1 _17775_ ( .A(_01616_ ), .B1(_02102_ ), .B2(_02103_ ), .ZN(_02104_ ) );
NAND2_X1 _17776_ ( .A1(_01624_ ), .A2(\ICACHE.cache_reg[6][22] ), .ZN(_02105_ ) );
NAND3_X1 _17777_ ( .A1(_01900_ ), .A2(_01901_ ), .A3(\ICACHE.cache_reg[7][22] ), .ZN(_02106_ ) );
AOI21_X1 _17778_ ( .A(_01623_ ), .B1(_02105_ ), .B2(_02106_ ), .ZN(_02107_ ) );
OAI21_X1 _17779_ ( .A(_07652_ ), .B1(_02104_ ), .B2(_02107_ ), .ZN(_02108_ ) );
NAND2_X1 _17780_ ( .A1(_01609_ ), .A2(\ICACHE.cache_reg[0][22] ), .ZN(_02109_ ) );
NAND3_X1 _17781_ ( .A1(_01906_ ), .A2(_01907_ ), .A3(\ICACHE.cache_reg[1][22] ), .ZN(_02110_ ) );
AOI21_X1 _17782_ ( .A(_07646_ ), .B1(_02109_ ), .B2(_02110_ ), .ZN(_02111_ ) );
NAND2_X1 _17783_ ( .A1(_07885_ ), .A2(\ICACHE.cache_reg[2][22] ), .ZN(_02112_ ) );
NAND3_X1 _17784_ ( .A1(_01911_ ), .A2(_01912_ ), .A3(\ICACHE.cache_reg[3][22] ), .ZN(_02113_ ) );
AOI21_X1 _17785_ ( .A(_07645_ ), .B1(_02112_ ), .B2(_02113_ ), .ZN(_02114_ ) );
OAI21_X1 _17786_ ( .A(_07836_ ), .B1(_02111_ ), .B2(_02114_ ), .ZN(_02115_ ) );
AOI21_X1 _17787_ ( .A(_01893_ ), .B1(_02108_ ), .B2(_02115_ ), .ZN(_02116_ ) );
MUX2_X1 _17788_ ( .A(\IDU.immI [2] ), .B(_02116_ ), .S(_02071_ ), .Z(_00772_ ) );
MUX2_X1 _17789_ ( .A(\BTB.btag_reg[0][0] ), .B(\BTB.btag_reg[1][0] ), .S(fanout_net_9 ), .Z(_02117_ ) );
XNOR2_X1 _17790_ ( .A(_02117_ ), .B(\ICACHE.state_$_MUX__S_A ), .ZN(_02118_ ) );
INV_X1 _17791_ ( .A(_02118_ ), .ZN(_02119_ ) );
MUX2_X1 _17792_ ( .A(\BTB.btag_reg[0][3] ), .B(\BTB.btag_reg[1][3] ), .S(fanout_net_9 ), .Z(_02120_ ) );
NAND2_X1 _17793_ ( .A1(_02120_ ), .A2(_07553_ ), .ZN(_02121_ ) );
OR2_X1 _17794_ ( .A1(_02120_ ), .A2(_07553_ ), .ZN(_02122_ ) );
MUX2_X1 _17795_ ( .A(\BTB.btag_reg[0][1] ), .B(\BTB.btag_reg[1][1] ), .S(fanout_net_9 ), .Z(_02123_ ) );
XNOR2_X1 _17796_ ( .A(_02123_ ), .B(\BTB.btag [1] ), .ZN(_02124_ ) );
AND4_X1 _17797_ ( .A1(_02119_ ), .A2(_02121_ ), .A3(_02122_ ), .A4(_02124_ ), .ZN(_02125_ ) );
MUX2_X1 _17798_ ( .A(\BTB.btag_reg[0][6] ), .B(\BTB.btag_reg[1][6] ), .S(fanout_net_9 ), .Z(_02126_ ) );
NAND2_X1 _17799_ ( .A1(_02126_ ), .A2(_07624_ ), .ZN(_02127_ ) );
OR2_X1 _17800_ ( .A1(_02126_ ), .A2(_07624_ ), .ZN(_02128_ ) );
MUX2_X1 _17801_ ( .A(\BTB.btag_reg[0][5] ), .B(\BTB.btag_reg[1][5] ), .S(fanout_net_9 ), .Z(_02129_ ) );
OR2_X1 _17802_ ( .A1(_02129_ ), .A2(_07560_ ), .ZN(_02130_ ) );
NAND2_X1 _17803_ ( .A1(_02129_ ), .A2(_07560_ ), .ZN(_02131_ ) );
AND4_X1 _17804_ ( .A1(_02127_ ), .A2(_02128_ ), .A3(_02130_ ), .A4(_02131_ ), .ZN(_02132_ ) );
MUX2_X1 _17805_ ( .A(\BTB.btag_reg[0][2] ), .B(\BTB.btag_reg[1][2] ), .S(fanout_net_9 ), .Z(_02133_ ) );
OR2_X1 _17806_ ( .A1(_02133_ ), .A2(_07603_ ), .ZN(_02134_ ) );
MUX2_X1 _17807_ ( .A(\BTB.btag_reg[0][7] ), .B(\BTB.btag_reg[1][7] ), .S(fanout_net_9 ), .Z(_02135_ ) );
OR2_X1 _17808_ ( .A1(_02135_ ), .A2(_07575_ ), .ZN(_02136_ ) );
NAND2_X1 _17809_ ( .A1(_02135_ ), .A2(_07575_ ), .ZN(_02137_ ) );
NAND2_X1 _17810_ ( .A1(_02133_ ), .A2(_07603_ ), .ZN(_02138_ ) );
AND4_X1 _17811_ ( .A1(_02134_ ), .A2(_02136_ ), .A3(_02137_ ), .A4(_02138_ ), .ZN(_02139_ ) );
AND3_X1 _17812_ ( .A1(_02125_ ), .A2(_02132_ ), .A3(_02139_ ), .ZN(_02140_ ) );
MUX2_X1 _17813_ ( .A(\BTB.btag_reg[0][9] ), .B(\BTB.btag_reg[1][9] ), .S(fanout_net_9 ), .Z(_02141_ ) );
XNOR2_X1 _17814_ ( .A(_02141_ ), .B(\BTB.btag [9] ), .ZN(_02142_ ) );
MUX2_X1 _17815_ ( .A(\BTB.btag_reg[0][8] ), .B(\BTB.btag_reg[1][8] ), .S(fanout_net_9 ), .Z(_02143_ ) );
OR2_X1 _17816_ ( .A1(_02143_ ), .A2(_07616_ ), .ZN(_02144_ ) );
NAND2_X1 _17817_ ( .A1(_02143_ ), .A2(_07616_ ), .ZN(_02145_ ) );
AND3_X1 _17818_ ( .A1(_02142_ ), .A2(_02144_ ), .A3(_02145_ ), .ZN(_02146_ ) );
MUX2_X1 _17819_ ( .A(\BTB.btag_reg[0][11] ), .B(\BTB.btag_reg[1][11] ), .S(fanout_net_9 ), .Z(_02147_ ) );
XNOR2_X1 _17820_ ( .A(_02147_ ), .B(\BTB.btag [11] ), .ZN(_02148_ ) );
MUX2_X1 _17821_ ( .A(\BTB.btag_reg[0][10] ), .B(\BTB.btag_reg[1][10] ), .S(fanout_net_9 ), .Z(_02149_ ) );
NAND2_X1 _17822_ ( .A1(_02149_ ), .A2(_07591_ ), .ZN(_02150_ ) );
OR2_X1 _17823_ ( .A1(_02149_ ), .A2(_07591_ ), .ZN(_02151_ ) );
AND3_X1 _17824_ ( .A1(_02148_ ), .A2(_02150_ ), .A3(_02151_ ), .ZN(_02152_ ) );
MUX2_X1 _17825_ ( .A(\BTB.btag_reg[0][12] ), .B(\BTB.btag_reg[1][12] ), .S(fanout_net_9 ), .Z(_02153_ ) );
XNOR2_X1 _17826_ ( .A(_02153_ ), .B(\BTB.btag [12] ), .ZN(_02154_ ) );
MUX2_X1 _17827_ ( .A(\BTB.btag_reg[0][4] ), .B(\BTB.btag_reg[1][4] ), .S(fanout_net_9 ), .Z(_02155_ ) );
INV_X1 _17828_ ( .A(\BTB.btag [4] ), .ZN(_02156_ ) );
NAND2_X1 _17829_ ( .A1(_02155_ ), .A2(_02156_ ), .ZN(_02157_ ) );
OR2_X1 _17830_ ( .A1(_02155_ ), .A2(_02156_ ), .ZN(_02158_ ) );
AND3_X1 _17831_ ( .A1(_02154_ ), .A2(_02157_ ), .A3(_02158_ ), .ZN(_02159_ ) );
AND3_X1 _17832_ ( .A1(_02146_ ), .A2(_02152_ ), .A3(_02159_ ), .ZN(_02160_ ) );
AND2_X1 _17833_ ( .A1(_02140_ ), .A2(_02160_ ), .ZN(_02161_ ) );
MUX2_X1 _17834_ ( .A(\BTB.jtag_reg[0][6] ), .B(\BTB.jtag_reg[1][6] ), .S(fanout_net_9 ), .Z(_02162_ ) );
OR2_X1 _17835_ ( .A1(_02162_ ), .A2(_07624_ ), .ZN(_02163_ ) );
MUX2_X1 _17836_ ( .A(\BTB.jtag_reg[0][5] ), .B(\BTB.jtag_reg[1][5] ), .S(fanout_net_9 ), .Z(_02164_ ) );
OR2_X1 _17837_ ( .A1(_02164_ ), .A2(_07560_ ), .ZN(_02165_ ) );
NAND2_X1 _17838_ ( .A1(_02162_ ), .A2(_07624_ ), .ZN(_02166_ ) );
NAND2_X1 _17839_ ( .A1(_02164_ ), .A2(_07560_ ), .ZN(_02167_ ) );
NAND4_X1 _17840_ ( .A1(_02163_ ), .A2(_02165_ ), .A3(_02166_ ), .A4(_02167_ ), .ZN(_02168_ ) );
MUX2_X1 _17841_ ( .A(\BTB.jtag_reg[0][2] ), .B(\BTB.jtag_reg[1][2] ), .S(fanout_net_9 ), .Z(_02169_ ) );
OR2_X1 _17842_ ( .A1(_02169_ ), .A2(_07603_ ), .ZN(_02170_ ) );
MUX2_X1 _17843_ ( .A(\BTB.jtag_reg[0][7] ), .B(\BTB.jtag_reg[1][7] ), .S(fanout_net_9 ), .Z(_02171_ ) );
OR2_X1 _17844_ ( .A1(_02171_ ), .A2(_07575_ ), .ZN(_02172_ ) );
NAND2_X1 _17845_ ( .A1(_02171_ ), .A2(_07575_ ), .ZN(_02173_ ) );
NAND2_X1 _17846_ ( .A1(_02169_ ), .A2(_07603_ ), .ZN(_02174_ ) );
NAND4_X1 _17847_ ( .A1(_02170_ ), .A2(_02172_ ), .A3(_02173_ ), .A4(_02174_ ), .ZN(_02175_ ) );
NOR2_X1 _17848_ ( .A1(_02168_ ), .A2(_02175_ ), .ZN(_02176_ ) );
MUX2_X1 _17849_ ( .A(\BTB.jtag_reg[0][0] ), .B(\BTB.jtag_reg[1][0] ), .S(fanout_net_9 ), .Z(_02177_ ) );
XNOR2_X1 _17850_ ( .A(_02177_ ), .B(\ICACHE.state_$_MUX__S_A ), .ZN(_02178_ ) );
INV_X1 _17851_ ( .A(_02178_ ), .ZN(_02179_ ) );
MUX2_X1 _17852_ ( .A(\BTB.jtag_reg[0][1] ), .B(\BTB.jtag_reg[1][1] ), .S(fanout_net_9 ), .Z(_02180_ ) );
OR2_X1 _17853_ ( .A1(_02180_ ), .A2(_07547_ ), .ZN(_02181_ ) );
MUX2_X1 _17854_ ( .A(\BTB.jtag_reg[0][3] ), .B(\BTB.jtag_reg[1][3] ), .S(fanout_net_9 ), .Z(_02182_ ) );
OR2_X1 _17855_ ( .A1(_02182_ ), .A2(_07553_ ), .ZN(_02183_ ) );
NAND2_X1 _17856_ ( .A1(_02182_ ), .A2(_07553_ ), .ZN(_02184_ ) );
NAND2_X1 _17857_ ( .A1(_02180_ ), .A2(_07547_ ), .ZN(_02185_ ) );
AND4_X1 _17858_ ( .A1(_02181_ ), .A2(_02183_ ), .A3(_02184_ ), .A4(_02185_ ), .ZN(_02186_ ) );
AND3_X1 _17859_ ( .A1(_02176_ ), .A2(_02179_ ), .A3(_02186_ ), .ZN(_02187_ ) );
MUX2_X1 _17860_ ( .A(\BTB.jtag_reg[0][9] ), .B(\BTB.jtag_reg[1][9] ), .S(fanout_net_9 ), .Z(_02188_ ) );
XNOR2_X1 _17861_ ( .A(_02188_ ), .B(\BTB.btag [9] ), .ZN(_02189_ ) );
MUX2_X1 _17862_ ( .A(\BTB.jtag_reg[0][8] ), .B(\BTB.jtag_reg[1][8] ), .S(fanout_net_9 ), .Z(_02190_ ) );
OR2_X1 _17863_ ( .A1(_02190_ ), .A2(_07616_ ), .ZN(_02191_ ) );
NAND2_X1 _17864_ ( .A1(_02190_ ), .A2(_07616_ ), .ZN(_02192_ ) );
AND3_X1 _17865_ ( .A1(_02189_ ), .A2(_02191_ ), .A3(_02192_ ), .ZN(_02193_ ) );
MUX2_X1 _17866_ ( .A(\BTB.jtag_reg[0][10] ), .B(\BTB.jtag_reg[1][10] ), .S(fanout_net_9 ), .Z(_02194_ ) );
XNOR2_X1 _17867_ ( .A(_02194_ ), .B(\BTB.btag [10] ), .ZN(_02195_ ) );
MUX2_X1 _17868_ ( .A(\BTB.jtag_reg[0][11] ), .B(\BTB.jtag_reg[1][11] ), .S(fanout_net_9 ), .Z(_02196_ ) );
OR2_X1 _17869_ ( .A1(_02196_ ), .A2(_07582_ ), .ZN(_02197_ ) );
NAND2_X1 _17870_ ( .A1(_02196_ ), .A2(_07582_ ), .ZN(_02198_ ) );
AND3_X1 _17871_ ( .A1(_02195_ ), .A2(_02197_ ), .A3(_02198_ ), .ZN(_02199_ ) );
MUX2_X1 _17872_ ( .A(\BTB.jtag_reg[0][12] ), .B(\BTB.jtag_reg[1][12] ), .S(fanout_net_9 ), .Z(_02200_ ) );
XNOR2_X1 _17873_ ( .A(_02200_ ), .B(\BTB.btag [12] ), .ZN(_02201_ ) );
MUX2_X1 _17874_ ( .A(\BTB.jtag_reg[0][4] ), .B(\BTB.jtag_reg[1][4] ), .S(fanout_net_9 ), .Z(_02202_ ) );
NAND2_X1 _17875_ ( .A1(_02202_ ), .A2(_02156_ ), .ZN(_02203_ ) );
OR2_X1 _17876_ ( .A1(_02202_ ), .A2(_02156_ ), .ZN(_02204_ ) );
AND3_X1 _17877_ ( .A1(_02201_ ), .A2(_02203_ ), .A3(_02204_ ), .ZN(_02205_ ) );
AND3_X1 _17878_ ( .A1(_02193_ ), .A2(_02199_ ), .A3(_02205_ ), .ZN(_02206_ ) );
AND2_X2 _17879_ ( .A1(_02187_ ), .A2(_02206_ ), .ZN(_02207_ ) );
NOR2_X1 _17880_ ( .A1(_02161_ ), .A2(_02207_ ), .ZN(_02208_ ) );
INV_X1 _17881_ ( .A(_02208_ ), .ZN(_02209_ ) );
AND3_X1 _17882_ ( .A1(_01594_ ), .A2(_05080_ ), .A3(_02209_ ), .ZN(_02210_ ) );
NOR2_X1 _17883_ ( .A1(_01594_ ), .A2(_05086_ ), .ZN(_02211_ ) );
NOR2_X1 _17884_ ( .A1(_02210_ ), .A2(_02211_ ), .ZN(_02212_ ) );
INV_X1 _17885_ ( .A(_02212_ ), .ZN(_02213_ ) );
NAND4_X1 _17886_ ( .A1(_02179_ ), .A2(_02201_ ), .A3(_02166_ ), .A4(_02172_ ), .ZN(_02214_ ) );
NAND4_X1 _17887_ ( .A1(_02181_ ), .A2(_02183_ ), .A3(_02184_ ), .A4(_02198_ ), .ZN(_02215_ ) );
NAND4_X1 _17888_ ( .A1(_02163_ ), .A2(_02165_ ), .A3(_02167_ ), .A4(_02185_ ), .ZN(_02216_ ) );
NOR3_X1 _17889_ ( .A1(_02214_ ), .A2(_02215_ ), .A3(_02216_ ), .ZN(_02217_ ) );
AND4_X1 _17890_ ( .A1(_02170_ ), .A2(_02191_ ), .A3(_02173_ ), .A4(_02203_ ), .ZN(_02218_ ) );
OR2_X1 _17891_ ( .A1(_02188_ ), .A2(_07610_ ), .ZN(_02219_ ) );
AND4_X1 _17892_ ( .A1(_02219_ ), .A2(_02204_ ), .A3(_02192_ ), .A4(_02174_ ), .ZN(_02220_ ) );
NAND2_X1 _17893_ ( .A1(_02194_ ), .A2(_07591_ ), .ZN(_02221_ ) );
AND2_X1 _17894_ ( .A1(_02197_ ), .A2(_02221_ ), .ZN(_02222_ ) );
NOR2_X1 _17895_ ( .A1(_02194_ ), .A2(_07591_ ), .ZN(_02223_ ) );
AOI21_X1 _17896_ ( .A(_02223_ ), .B1(_07610_ ), .B2(_02188_ ), .ZN(_02224_ ) );
AND4_X1 _17897_ ( .A1(_02218_ ), .A2(_02220_ ), .A3(_02222_ ), .A4(_02224_ ), .ZN(_02225_ ) );
AND2_X1 _17898_ ( .A1(_02217_ ), .A2(_02225_ ), .ZN(_02226_ ) );
NAND4_X1 _17899_ ( .A1(_02119_ ), .A2(_02154_ ), .A3(_02127_ ), .A4(_02136_ ), .ZN(_02227_ ) );
OR2_X1 _17900_ ( .A1(_02123_ ), .A2(_07547_ ), .ZN(_02228_ ) );
NAND2_X1 _17901_ ( .A1(_02147_ ), .A2(_07582_ ), .ZN(_02229_ ) );
NAND4_X1 _17902_ ( .A1(_02228_ ), .A2(_02122_ ), .A3(_02121_ ), .A4(_02229_ ), .ZN(_02230_ ) );
NAND2_X1 _17903_ ( .A1(_02123_ ), .A2(_07547_ ), .ZN(_02231_ ) );
NAND4_X1 _17904_ ( .A1(_02128_ ), .A2(_02130_ ), .A3(_02131_ ), .A4(_02231_ ), .ZN(_02232_ ) );
NOR3_X1 _17905_ ( .A1(_02227_ ), .A2(_02230_ ), .A3(_02232_ ), .ZN(_02233_ ) );
AND4_X1 _17906_ ( .A1(_02134_ ), .A2(_02144_ ), .A3(_02137_ ), .A4(_02157_ ), .ZN(_02234_ ) );
OR2_X1 _17907_ ( .A1(_02141_ ), .A2(_07610_ ), .ZN(_02235_ ) );
AND4_X1 _17908_ ( .A1(_02235_ ), .A2(_02158_ ), .A3(_02145_ ), .A4(_02138_ ), .ZN(_02236_ ) );
OR2_X1 _17909_ ( .A1(_02147_ ), .A2(_07582_ ), .ZN(_02237_ ) );
NAND2_X1 _17910_ ( .A1(_02141_ ), .A2(_07610_ ), .ZN(_02238_ ) );
AND4_X1 _17911_ ( .A1(_02237_ ), .A2(_02151_ ), .A3(_02150_ ), .A4(_02238_ ), .ZN(_02239_ ) );
AND3_X1 _17912_ ( .A1(_02234_ ), .A2(_02236_ ), .A3(_02239_ ), .ZN(_02240_ ) );
AND2_X1 _17913_ ( .A1(_02233_ ), .A2(_02240_ ), .ZN(_02241_ ) );
NOR2_X1 _17914_ ( .A1(_02226_ ), .A2(_02241_ ), .ZN(_02242_ ) );
INV_X1 _17915_ ( .A(_02242_ ), .ZN(_02243_ ) );
NAND3_X1 _17916_ ( .A1(\BTB.btag [1] ), .A2(\BTB.btag [0] ), .A3(\BTB.bindex ), .ZN(_02244_ ) );
OR3_X1 _17917_ ( .A1(_02244_ ), .A2(_07553_ ), .A3(_07603_ ), .ZN(_02245_ ) );
NOR3_X1 _17918_ ( .A1(_02245_ ), .A2(_07560_ ), .A3(_02156_ ), .ZN(_02246_ ) );
AND3_X1 _17919_ ( .A1(_02246_ ), .A2(\BTB.btag [7] ), .A3(\BTB.btag [6] ), .ZN(_02247_ ) );
AND2_X1 _17920_ ( .A1(_02247_ ), .A2(\BTB.btag [8] ), .ZN(_02248_ ) );
AND2_X1 _17921_ ( .A1(_02248_ ), .A2(\BTB.btag [9] ), .ZN(_02249_ ) );
AND2_X1 _17922_ ( .A1(_02249_ ), .A2(\BTB.btag [10] ), .ZN(_02250_ ) );
AND2_X1 _17923_ ( .A1(_02250_ ), .A2(\BTB.btag [11] ), .ZN(_02251_ ) );
AND2_X1 _17924_ ( .A1(_02251_ ), .A2(\BTB.btag [12] ), .ZN(_02252_ ) );
AND2_X1 _17925_ ( .A1(_02252_ ), .A2(\BTB.pc_i [16] ), .ZN(_02253_ ) );
AND2_X1 _17926_ ( .A1(_02253_ ), .A2(\BTB.pc_i [17] ), .ZN(_02254_ ) );
AND2_X1 _17927_ ( .A1(_02254_ ), .A2(\BTB.pc_i [18] ), .ZN(_02255_ ) );
AND2_X1 _17928_ ( .A1(_02255_ ), .A2(\BTB.pc_i [19] ), .ZN(_02256_ ) );
AND2_X1 _17929_ ( .A1(\BTB.pc_i [23] ), .A2(\BTB.pc_i [22] ), .ZN(_02257_ ) );
AND2_X1 _17930_ ( .A1(\BTB.pc_i [25] ), .A2(\BTB.pc_i [24] ), .ZN(_02258_ ) );
AND3_X1 _17931_ ( .A1(_02258_ ), .A2(\BTB.pc_i [21] ), .A3(\BTB.pc_i [20] ), .ZN(_02259_ ) );
AND3_X1 _17932_ ( .A1(_02256_ ), .A2(_02257_ ), .A3(_02259_ ), .ZN(_02260_ ) );
AND3_X1 _17933_ ( .A1(_02260_ ), .A2(\BTB.pc_i [27] ), .A3(\BTB.pc_i [26] ), .ZN(_02261_ ) );
AND3_X1 _17934_ ( .A1(_02261_ ), .A2(\BTB.pc_i [29] ), .A3(\BTB.pc_i [28] ), .ZN(_02262_ ) );
AOI21_X1 _17935_ ( .A(_02243_ ), .B1(_02262_ ), .B2(\BTB.pc_i [30] ), .ZN(_02263_ ) );
AND3_X1 _17936_ ( .A1(_01595_ ), .A2(_05080_ ), .A3(_02263_ ), .ZN(_02264_ ) );
OAI21_X1 _17937_ ( .A(\BTB.pc_i [31] ), .B1(_02213_ ), .B2(_02264_ ), .ZN(_02265_ ) );
INV_X1 _17938_ ( .A(_02262_ ), .ZN(_02266_ ) );
NOR4_X1 _17939_ ( .A1(_02266_ ), .A2(\BTB.pc_i [31] ), .A3(_07838_ ), .A4(_02243_ ), .ZN(_02267_ ) );
NAND4_X1 _17940_ ( .A1(_01596_ ), .A2(_05252_ ), .A3(_01597_ ), .A4(_02267_ ), .ZN(_02268_ ) );
AND2_X1 _17941_ ( .A1(_04331_ ), .A2(_03805_ ), .ZN(_02269_ ) );
INV_X1 _17942_ ( .A(_02269_ ), .ZN(_02270_ ) );
BUF_X4 _17943_ ( .A(_02270_ ), .Z(_02271_ ) );
OAI211_X1 _17944_ ( .A(_02265_ ), .B(_02268_ ), .C1(_05085_ ), .C2(_02271_ ), .ZN(_00773_ ) );
AND2_X1 _17945_ ( .A1(_01594_ ), .A2(_05080_ ), .ZN(_02272_ ) );
BUF_X4 _17946_ ( .A(_02272_ ), .Z(_02273_ ) );
BUF_X4 _17947_ ( .A(_02209_ ), .Z(_02274_ ) );
AND4_X1 _17948_ ( .A1(\BTB.pc_i [19] ), .A2(\BTB.pc_i [18] ), .A3(\BTB.pc_i [23] ), .A4(\BTB.pc_i [22] ), .ZN(_02275_ ) );
AND3_X1 _17949_ ( .A1(_02254_ ), .A2(_02259_ ), .A3(_02275_ ), .ZN(_02276_ ) );
AND3_X1 _17950_ ( .A1(_02276_ ), .A2(\BTB.pc_i [27] ), .A3(\BTB.pc_i [26] ), .ZN(_02277_ ) );
AND3_X1 _17951_ ( .A1(_02277_ ), .A2(\BTB.pc_i [29] ), .A3(\BTB.pc_i [28] ), .ZN(_02278_ ) );
AOI21_X1 _17952_ ( .A(_02274_ ), .B1(_02278_ ), .B2(\BTB.pc_i [30] ), .ZN(_02279_ ) );
OAI211_X1 _17953_ ( .A(_02273_ ), .B(_02279_ ), .C1(\BTB.pc_i [30] ), .C2(_02278_ ), .ZN(_02280_ ) );
BUF_X4 _17954_ ( .A(_02270_ ), .Z(_02281_ ) );
OAI221_X1 _17955_ ( .A(_02280_ ), .B1(_05107_ ), .B2(_02281_ ), .C1(_02212_ ), .C2(_07838_ ), .ZN(_00774_ ) );
BUF_X4 _17956_ ( .A(_02273_ ), .Z(_02282_ ) );
INV_X1 _17957_ ( .A(\BTB.pc_i [21] ), .ZN(_02283_ ) );
AND2_X2 _17958_ ( .A1(_02246_ ), .A2(\BTB.btag [6] ), .ZN(_02284_ ) );
AND2_X1 _17959_ ( .A1(\BTB.pc_i [19] ), .A2(\BTB.pc_i [18] ), .ZN(_02285_ ) );
AND4_X1 _17960_ ( .A1(\BTB.pc_i [17] ), .A2(\BTB.pc_i [16] ), .A3(\BTB.btag [12] ), .A4(\BTB.btag [11] ), .ZN(_02286_ ) );
AND2_X1 _17961_ ( .A1(\BTB.btag [8] ), .A2(\BTB.btag [7] ), .ZN(_02287_ ) );
AND4_X1 _17962_ ( .A1(\BTB.btag [10] ), .A2(_02286_ ), .A3(\BTB.btag [9] ), .A4(_02287_ ), .ZN(_02288_ ) );
AND3_X1 _17963_ ( .A1(_02284_ ), .A2(_02285_ ), .A3(_02288_ ), .ZN(_02289_ ) );
INV_X1 _17964_ ( .A(_02289_ ), .ZN(_02290_ ) );
INV_X1 _17965_ ( .A(\BTB.pc_i [20] ), .ZN(_02291_ ) );
OAI21_X1 _17966_ ( .A(_02283_ ), .B1(_02290_ ), .B2(_02291_ ), .ZN(_02292_ ) );
AND3_X1 _17967_ ( .A1(_02255_ ), .A2(\BTB.pc_i [20] ), .A3(\BTB.pc_i [19] ), .ZN(_02293_ ) );
AND2_X1 _17968_ ( .A1(_02293_ ), .A2(\BTB.pc_i [21] ), .ZN(_02294_ ) );
INV_X1 _17969_ ( .A(_02294_ ), .ZN(_02295_ ) );
NAND4_X1 _17970_ ( .A1(_02282_ ), .A2(_02208_ ), .A3(_02292_ ), .A4(_02295_ ), .ZN(_02296_ ) );
OAI221_X1 _17971_ ( .A(_02296_ ), .B1(_04251_ ), .B2(_02281_ ), .C1(_02212_ ), .C2(_02283_ ), .ZN(_00775_ ) );
AND3_X1 _17972_ ( .A1(_02253_ ), .A2(\BTB.pc_i [17] ), .A3(_02285_ ), .ZN(_02297_ ) );
AOI21_X1 _17973_ ( .A(_02209_ ), .B1(_02297_ ), .B2(\BTB.pc_i [20] ), .ZN(_02298_ ) );
OAI211_X1 _17974_ ( .A(_02273_ ), .B(_02298_ ), .C1(\BTB.pc_i [20] ), .C2(_02256_ ), .ZN(_02299_ ) );
OAI221_X1 _17975_ ( .A(_02299_ ), .B1(_04252_ ), .B2(_02281_ ), .C1(_02212_ ), .C2(_02291_ ), .ZN(_00776_ ) );
BUF_X4 _17976_ ( .A(_02209_ ), .Z(_02300_ ) );
NOR2_X1 _17977_ ( .A1(_02297_ ), .A2(_02300_ ), .ZN(_02301_ ) );
OAI211_X1 _17978_ ( .A(_02282_ ), .B(_02301_ ), .C1(\BTB.pc_i [19] ), .C2(_02255_ ), .ZN(_02302_ ) );
BUF_X4 _17979_ ( .A(_05080_ ), .Z(_02303_ ) );
BUF_X4 _17980_ ( .A(_02303_ ), .Z(_02304_ ) );
INV_X1 _17981_ ( .A(_01594_ ), .ZN(_02305_ ) );
BUF_X4 _17982_ ( .A(_02305_ ), .Z(_02306_ ) );
OAI211_X1 _17983_ ( .A(\BTB.pc_i [19] ), .B(_02304_ ), .C1(_02306_ ), .C2(_02300_ ), .ZN(_02307_ ) );
OAI211_X1 _17984_ ( .A(_02302_ ), .B(_02307_ ), .C1(_05156_ ), .C2(_02271_ ), .ZN(_00777_ ) );
AOI21_X1 _17985_ ( .A(_02274_ ), .B1(_02254_ ), .B2(\BTB.pc_i [18] ), .ZN(_02308_ ) );
OAI211_X1 _17986_ ( .A(_02282_ ), .B(_02308_ ), .C1(\BTB.pc_i [18] ), .C2(_02254_ ), .ZN(_02309_ ) );
OAI211_X1 _17987_ ( .A(\BTB.pc_i [18] ), .B(_02304_ ), .C1(_02306_ ), .C2(_02300_ ), .ZN(_02310_ ) );
OAI211_X1 _17988_ ( .A(_02309_ ), .B(_02310_ ), .C1(_05165_ ), .C2(_02271_ ), .ZN(_00778_ ) );
AOI21_X1 _17989_ ( .A(_02274_ ), .B1(_02253_ ), .B2(\BTB.pc_i [17] ), .ZN(_02311_ ) );
OAI211_X1 _17990_ ( .A(_02282_ ), .B(_02311_ ), .C1(\BTB.pc_i [17] ), .C2(_02253_ ), .ZN(_02312_ ) );
OAI211_X1 _17991_ ( .A(\BTB.pc_i [17] ), .B(_02304_ ), .C1(_02306_ ), .C2(_02300_ ), .ZN(_02313_ ) );
OAI211_X1 _17992_ ( .A(_02312_ ), .B(_02313_ ), .C1(_04242_ ), .C2(_02271_ ), .ZN(_00779_ ) );
AOI21_X1 _17993_ ( .A(_02274_ ), .B1(_02252_ ), .B2(\BTB.pc_i [16] ), .ZN(_02314_ ) );
OAI211_X1 _17994_ ( .A(_02282_ ), .B(_02314_ ), .C1(\BTB.pc_i [16] ), .C2(_02252_ ), .ZN(_02315_ ) );
OAI211_X1 _17995_ ( .A(\BTB.pc_i [16] ), .B(_02304_ ), .C1(_02306_ ), .C2(_02300_ ), .ZN(_02316_ ) );
OAI211_X1 _17996_ ( .A(_02315_ ), .B(_02316_ ), .C1(_04243_ ), .C2(_02271_ ), .ZN(_00780_ ) );
BUF_X4 _17997_ ( .A(_01595_ ), .Z(_02317_ ) );
INV_X1 _17998_ ( .A(_02251_ ), .ZN(_02318_ ) );
OAI21_X1 _17999_ ( .A(_02242_ ), .B1(_02318_ ), .B2(_07632_ ), .ZN(_02319_ ) );
AND3_X1 _18000_ ( .A1(_02287_ ), .A2(\BTB.btag [10] ), .A3(\BTB.btag [9] ), .ZN(_02320_ ) );
NAND3_X1 _18001_ ( .A1(_02284_ ), .A2(\BTB.btag [11] ), .A3(_02320_ ), .ZN(_02321_ ) );
AOI21_X1 _18002_ ( .A(_02319_ ), .B1(_07632_ ), .B2(_02321_ ), .ZN(_02322_ ) );
NAND4_X1 _18003_ ( .A1(_02172_ ), .A2(_02163_ ), .A3(_02173_ ), .A4(_02166_ ), .ZN(_02323_ ) );
NAND4_X1 _18004_ ( .A1(_02204_ ), .A2(_02165_ ), .A3(_02203_ ), .A4(_02167_ ), .ZN(_02324_ ) );
NOR2_X1 _18005_ ( .A1(_02323_ ), .A2(_02324_ ), .ZN(_02325_ ) );
XNOR2_X1 _18006_ ( .A(_02180_ ), .B(\BTB.btag [1] ), .ZN(_02326_ ) );
AND4_X1 _18007_ ( .A1(_02170_ ), .A2(_02183_ ), .A3(_02174_ ), .A4(_02184_ ), .ZN(_02327_ ) );
AND4_X1 _18008_ ( .A1(_02179_ ), .A2(_02325_ ), .A3(_02326_ ), .A4(_02327_ ), .ZN(_02328_ ) );
AND3_X1 _18009_ ( .A1(_02193_ ), .A2(_02199_ ), .A3(_02201_ ), .ZN(_02329_ ) );
NAND2_X2 _18010_ ( .A1(_02328_ ), .A2(_02329_ ), .ZN(_02330_ ) );
MUX2_X1 _18011_ ( .A(_03960_ ), .B(_04005_ ), .S(fanout_net_9 ), .Z(_02331_ ) );
NOR2_X1 _18012_ ( .A1(_02330_ ), .A2(_02331_ ), .ZN(_02332_ ) );
OAI211_X1 _18013_ ( .A(_02317_ ), .B(_02303_ ), .C1(_02322_ ), .C2(_02332_ ), .ZN(_02333_ ) );
INV_X1 _18014_ ( .A(_02241_ ), .ZN(_02334_ ) );
NOR2_X1 _18015_ ( .A1(_02334_ ), .A2(_02226_ ), .ZN(_02335_ ) );
INV_X1 _18016_ ( .A(_02335_ ), .ZN(_02336_ ) );
NAND4_X1 _18017_ ( .A1(_07877_ ), .A2(_02303_ ), .A3(_01592_ ), .A4(_02336_ ), .ZN(_02337_ ) );
NAND2_X1 _18018_ ( .A1(_02337_ ), .A2(_02303_ ), .ZN(_02338_ ) );
OAI221_X1 _18019_ ( .A(_02333_ ), .B1(_05207_ ), .B2(_02281_ ), .C1(_02338_ ), .C2(_07632_ ), .ZN(_00781_ ) );
INV_X1 _18020_ ( .A(_02250_ ), .ZN(_02339_ ) );
OAI21_X1 _18021_ ( .A(_02242_ ), .B1(_02339_ ), .B2(_07582_ ), .ZN(_02340_ ) );
NAND2_X1 _18022_ ( .A1(_02284_ ), .A2(_02320_ ), .ZN(_02341_ ) );
AOI21_X1 _18023_ ( .A(_02340_ ), .B1(_07582_ ), .B2(_02341_ ), .ZN(_02342_ ) );
MUX2_X1 _18024_ ( .A(_03966_ ), .B(_04008_ ), .S(fanout_net_9 ), .Z(_02343_ ) );
NOR2_X1 _18025_ ( .A1(_02330_ ), .A2(_02343_ ), .ZN(_02344_ ) );
OAI211_X1 _18026_ ( .A(_02317_ ), .B(_02303_ ), .C1(_02342_ ), .C2(_02344_ ), .ZN(_02345_ ) );
OAI221_X1 _18027_ ( .A(_02345_ ), .B1(_05218_ ), .B2(_02281_ ), .C1(_02338_ ), .C2(_07582_ ), .ZN(_00782_ ) );
NAND2_X1 _18028_ ( .A1(_02242_ ), .A2(_02339_ ), .ZN(_02346_ ) );
NAND3_X1 _18029_ ( .A1(_02284_ ), .A2(\BTB.btag [9] ), .A3(_02287_ ), .ZN(_02347_ ) );
AOI21_X1 _18030_ ( .A(_02346_ ), .B1(_07591_ ), .B2(_02347_ ), .ZN(_02348_ ) );
MUX2_X1 _18031_ ( .A(_03981_ ), .B(_04017_ ), .S(fanout_net_9 ), .Z(_02349_ ) );
NOR2_X1 _18032_ ( .A1(_02330_ ), .A2(_02349_ ), .ZN(_02350_ ) );
OAI211_X1 _18033_ ( .A(_02317_ ), .B(_02303_ ), .C1(_02348_ ), .C2(_02350_ ), .ZN(_02351_ ) );
OAI221_X1 _18034_ ( .A(_02351_ ), .B1(_04226_ ), .B2(_02281_ ), .C1(_02338_ ), .C2(_07591_ ), .ZN(_00783_ ) );
INV_X1 _18035_ ( .A(_02226_ ), .ZN(_02352_ ) );
INV_X1 _18036_ ( .A(_02249_ ), .ZN(_02353_ ) );
NAND3_X1 _18037_ ( .A1(_02352_ ), .A2(_02334_ ), .A3(_02353_ ), .ZN(_02354_ ) );
INV_X1 _18038_ ( .A(_02248_ ), .ZN(_02355_ ) );
AOI21_X1 _18039_ ( .A(_02354_ ), .B1(_07610_ ), .B2(_02355_ ), .ZN(_02356_ ) );
MUX2_X1 _18040_ ( .A(_03984_ ), .B(_04018_ ), .S(fanout_net_9 ), .Z(_02357_ ) );
NOR2_X1 _18041_ ( .A1(_02330_ ), .A2(_02357_ ), .ZN(_02358_ ) );
OAI211_X1 _18042_ ( .A(_02317_ ), .B(_02303_ ), .C1(_02356_ ), .C2(_02358_ ), .ZN(_02359_ ) );
OAI221_X1 _18043_ ( .A(_02359_ ), .B1(_04227_ ), .B2(_02281_ ), .C1(_02338_ ), .C2(_07610_ ), .ZN(_00784_ ) );
AND2_X1 _18044_ ( .A1(_02272_ ), .A2(_02242_ ), .ZN(_02360_ ) );
AND2_X1 _18045_ ( .A1(_02261_ ), .A2(\BTB.pc_i [28] ), .ZN(_02361_ ) );
XOR2_X1 _18046_ ( .A(_02361_ ), .B(\BTB.pc_i [29] ), .Z(_02362_ ) );
AOI22_X1 _18047_ ( .A1(_02360_ ), .A2(_02362_ ), .B1(\EXU.dnpc_o [29] ), .B2(_02269_ ), .ZN(_02363_ ) );
OAI21_X1 _18048_ ( .A(_02363_ ), .B1(_02273_ ), .B2(_02269_ ), .ZN(_02364_ ) );
MUX2_X1 _18049_ ( .A(\BTB.pc_i [29] ), .B(_02364_ ), .S(_02212_ ), .Z(_00785_ ) );
NAND3_X1 _18050_ ( .A1(_02352_ ), .A2(_02334_ ), .A3(_02355_ ), .ZN(_02365_ ) );
INV_X1 _18051_ ( .A(_02247_ ), .ZN(_02366_ ) );
AOI21_X1 _18052_ ( .A(_02365_ ), .B1(_07616_ ), .B2(_02366_ ), .ZN(_02367_ ) );
MUX2_X1 _18053_ ( .A(_03988_ ), .B(_04019_ ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02368_ ) );
NOR2_X1 _18054_ ( .A1(_02330_ ), .A2(_02368_ ), .ZN(_02369_ ) );
OAI211_X1 _18055_ ( .A(_01595_ ), .B(_02303_ ), .C1(_02367_ ), .C2(_02369_ ), .ZN(_02370_ ) );
BUF_X4 _18056_ ( .A(_02270_ ), .Z(_02371_ ) );
OAI221_X1 _18057_ ( .A(_02370_ ), .B1(_05268_ ), .B2(_02371_ ), .C1(_02338_ ), .C2(_07616_ ), .ZN(_00786_ ) );
MUX2_X1 _18058_ ( .A(_03991_ ), .B(_04020_ ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02372_ ) );
OR2_X1 _18059_ ( .A1(_02330_ ), .A2(_02372_ ), .ZN(_02373_ ) );
XNOR2_X1 _18060_ ( .A(_02284_ ), .B(\BTB.btag [7] ), .ZN(_02374_ ) );
OAI21_X1 _18061_ ( .A(_02373_ ), .B1(_02243_ ), .B2(_02374_ ), .ZN(_02375_ ) );
NAND4_X1 _18062_ ( .A1(_07877_ ), .A2(_05252_ ), .A3(_01592_ ), .A4(_02375_ ), .ZN(_02376_ ) );
OAI221_X1 _18063_ ( .A(_02376_ ), .B1(_05276_ ), .B2(_02371_ ), .C1(_02338_ ), .C2(_07575_ ), .ZN(_00787_ ) );
MUX2_X1 _18064_ ( .A(_03995_ ), .B(_04021_ ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02377_ ) );
OR2_X1 _18065_ ( .A1(_02330_ ), .A2(_02377_ ), .ZN(_02378_ ) );
XNOR2_X1 _18066_ ( .A(_02246_ ), .B(\BTB.btag [6] ), .ZN(_02379_ ) );
OAI21_X1 _18067_ ( .A(_02378_ ), .B1(_02243_ ), .B2(_02379_ ), .ZN(_02380_ ) );
NAND4_X1 _18068_ ( .A1(_07877_ ), .A2(_05252_ ), .A3(_01592_ ), .A4(_02380_ ), .ZN(_02381_ ) );
OAI221_X1 _18069_ ( .A(_02381_ ), .B1(_05288_ ), .B2(_02371_ ), .C1(_02338_ ), .C2(_07624_ ), .ZN(_00788_ ) );
INV_X1 _18070_ ( .A(_02246_ ), .ZN(_02382_ ) );
OAI21_X1 _18071_ ( .A(_07560_ ), .B1(_02245_ ), .B2(_02156_ ), .ZN(_02383_ ) );
AND3_X1 _18072_ ( .A1(_02242_ ), .A2(_02382_ ), .A3(_02383_ ), .ZN(_02384_ ) );
MUX2_X1 _18073_ ( .A(_03999_ ), .B(_04022_ ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02385_ ) );
NOR2_X1 _18074_ ( .A1(_02330_ ), .A2(_02385_ ), .ZN(_02386_ ) );
OAI211_X1 _18075_ ( .A(_01595_ ), .B(_02303_ ), .C1(_02384_ ), .C2(_02386_ ), .ZN(_02387_ ) );
OAI221_X1 _18076_ ( .A(_02387_ ), .B1(_05297_ ), .B2(_02371_ ), .C1(_02338_ ), .C2(_07560_ ), .ZN(_00789_ ) );
OAI211_X1 _18077_ ( .A(\BTB.pc_i [1] ), .B(_05252_ ), .C1(_02306_ ), .C2(_02208_ ), .ZN(_02388_ ) );
NOR2_X1 _18078_ ( .A1(\BTB.bsnpc_reg[0][1] ), .A2(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .ZN(_02389_ ) );
NAND4_X1 _18079_ ( .A1(_02136_ ), .A2(_02128_ ), .A3(_02137_ ), .A4(_02127_ ), .ZN(_02390_ ) );
NAND4_X1 _18080_ ( .A1(_02158_ ), .A2(_02130_ ), .A3(_02157_ ), .A4(_02131_ ), .ZN(_02391_ ) );
NOR2_X1 _18081_ ( .A1(_02390_ ), .A2(_02391_ ), .ZN(_02392_ ) );
AND4_X1 _18082_ ( .A1(_02134_ ), .A2(_02122_ ), .A3(_02138_ ), .A4(_02121_ ), .ZN(_02393_ ) );
AND4_X1 _18083_ ( .A1(_02119_ ), .A2(_02392_ ), .A3(_02124_ ), .A4(_02393_ ), .ZN(_02394_ ) );
AND3_X1 _18084_ ( .A1(_02146_ ), .A2(_02152_ ), .A3(_02154_ ), .ZN(_02395_ ) );
NAND2_X1 _18085_ ( .A1(_02394_ ), .A2(_02395_ ), .ZN(_02396_ ) );
AOI211_X1 _18086_ ( .A(_02389_ ), .B(_02396_ ), .C1(_03852_ ), .C2(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .ZN(_02397_ ) );
NAND2_X1 _18087_ ( .A1(_02397_ ), .A2(_02330_ ), .ZN(_02398_ ) );
AND2_X1 _18088_ ( .A1(_02328_ ), .A2(_02329_ ), .ZN(_02399_ ) );
MUX2_X1 _18089_ ( .A(\BTB.jsnpc_reg[0][1] ), .B(\BTB.jsnpc_reg[1][1] ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02400_ ) );
NAND2_X1 _18090_ ( .A1(_02399_ ), .A2(_02400_ ), .ZN(_02401_ ) );
NAND2_X1 _18091_ ( .A1(_02398_ ), .A2(_02401_ ), .ZN(_02402_ ) );
NAND4_X1 _18092_ ( .A1(_07877_ ), .A2(_05252_ ), .A3(_01592_ ), .A4(_02402_ ), .ZN(_02403_ ) );
OAI211_X1 _18093_ ( .A(_02388_ ), .B(_02403_ ), .C1(_04232_ ), .C2(_02271_ ), .ZN(_00790_ ) );
OAI211_X1 _18094_ ( .A(\BTB.pc_i [0] ), .B(_05252_ ), .C1(_02306_ ), .C2(_02208_ ), .ZN(_02404_ ) );
NOR2_X1 _18095_ ( .A1(\BTB.bsnpc_reg[0][0] ), .A2(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .ZN(_02405_ ) );
AOI211_X1 _18096_ ( .A(_02405_ ), .B(_02396_ ), .C1(_03854_ ), .C2(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .ZN(_02406_ ) );
NAND2_X1 _18097_ ( .A1(_02406_ ), .A2(_02330_ ), .ZN(_02407_ ) );
MUX2_X1 _18098_ ( .A(\BTB.jsnpc_reg[0][0] ), .B(\BTB.jsnpc_reg[1][0] ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02408_ ) );
NAND2_X1 _18099_ ( .A1(_02399_ ), .A2(_02408_ ), .ZN(_02409_ ) );
NAND2_X1 _18100_ ( .A1(_02407_ ), .A2(_02409_ ), .ZN(_02410_ ) );
NAND4_X1 _18101_ ( .A1(_07877_ ), .A2(_05252_ ), .A3(_01592_ ), .A4(_02410_ ), .ZN(_02411_ ) );
OAI211_X1 _18102_ ( .A(_02404_ ), .B(_02411_ ), .C1(_04233_ ), .C2(_02271_ ), .ZN(_00791_ ) );
MUX2_X1 _18103_ ( .A(\BTB.bsnpc_reg[0]_$_NOT__A_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ), .B(\BTB.bsnpc_reg[0]_$_NOT__A_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02412_ ) );
NAND3_X1 _18104_ ( .A1(_02328_ ), .A2(_02329_ ), .A3(_02412_ ), .ZN(_02413_ ) );
MUX2_X1 _18105_ ( .A(\BTB.bsnpc_reg[0]_$_NOT__A_Y ), .B(\BTB.bsnpc_reg[1]_$_NOT__A_Y ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02414_ ) );
AND3_X1 _18106_ ( .A1(_02394_ ), .A2(_02395_ ), .A3(_02414_ ), .ZN(_02415_ ) );
XNOR2_X1 _18107_ ( .A(_02245_ ), .B(_02156_ ), .ZN(_02416_ ) );
AOI21_X1 _18108_ ( .A(_02415_ ), .B1(_02396_ ), .B2(_02416_ ), .ZN(_02417_ ) );
OAI211_X1 _18109_ ( .A(_02273_ ), .B(_02413_ ), .C1(_02207_ ), .C2(_02417_ ), .ZN(_02418_ ) );
INV_X1 _18110_ ( .A(_02211_ ), .ZN(_02419_ ) );
OAI221_X1 _18111_ ( .A(_02418_ ), .B1(_04235_ ), .B2(_02371_ ), .C1(_02419_ ), .C2(_02156_ ), .ZN(_00792_ ) );
MUX2_X1 _18112_ ( .A(\BTB.bsnpc_reg[0]_$_NOT__A_1_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ), .B(\BTB.bsnpc_reg[0]_$_NOT__A_1_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02420_ ) );
NAND2_X1 _18113_ ( .A1(_02399_ ), .A2(_02420_ ), .ZN(_02421_ ) );
AND2_X1 _18114_ ( .A1(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .A2(\BTB.bsnpc_reg[1]_$_NOT__A_1_Y ), .ZN(_02422_ ) );
INV_X1 _18115_ ( .A(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .ZN(_02423_ ) );
AOI21_X1 _18116_ ( .A(_02422_ ), .B1(_02423_ ), .B2(\BTB.bsnpc_reg[0]_$_NOT__A_1_Y ), .ZN(_02424_ ) );
NAND3_X1 _18117_ ( .A1(_02233_ ), .A2(_02240_ ), .A3(_02424_ ), .ZN(_02425_ ) );
NOR2_X1 _18118_ ( .A1(_02244_ ), .A2(_07603_ ), .ZN(_02426_ ) );
XNOR2_X1 _18119_ ( .A(_02426_ ), .B(\BTB.btag [3] ), .ZN(_02427_ ) );
OAI21_X1 _18120_ ( .A(_02425_ ), .B1(_02241_ ), .B2(_02427_ ), .ZN(_02428_ ) );
OAI211_X1 _18121_ ( .A(_02273_ ), .B(_02421_ ), .C1(_02207_ ), .C2(_02428_ ), .ZN(_02429_ ) );
OAI221_X1 _18122_ ( .A(_02429_ ), .B1(_04236_ ), .B2(_02371_ ), .C1(_07553_ ), .C2(_02419_ ), .ZN(_00793_ ) );
MUX2_X1 _18123_ ( .A(\BTB.bsnpc_reg[0]_$_NOT__A_2_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ), .B(\BTB.bsnpc_reg[0]_$_NOT__A_2_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02430_ ) );
NAND3_X1 _18124_ ( .A1(_02328_ ), .A2(_02329_ ), .A3(_02430_ ), .ZN(_02431_ ) );
MUX2_X1 _18125_ ( .A(\BTB.bsnpc_reg[0]_$_NOT__A_2_Y ), .B(\BTB.bsnpc_reg[1]_$_NOT__A_2_Y ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02432_ ) );
AND3_X1 _18126_ ( .A1(_02394_ ), .A2(_02395_ ), .A3(_02432_ ), .ZN(_02433_ ) );
XNOR2_X1 _18127_ ( .A(_02244_ ), .B(_07603_ ), .ZN(_02434_ ) );
AOI21_X1 _18128_ ( .A(_02433_ ), .B1(_02396_ ), .B2(_02434_ ), .ZN(_02435_ ) );
OAI211_X1 _18129_ ( .A(_02273_ ), .B(_02431_ ), .C1(_02207_ ), .C2(_02435_ ), .ZN(_02436_ ) );
OAI221_X1 _18130_ ( .A(_02436_ ), .B1(_04237_ ), .B2(_02371_ ), .C1(_02419_ ), .C2(_07603_ ), .ZN(_00794_ ) );
INV_X1 _18131_ ( .A(_02207_ ), .ZN(_02437_ ) );
AND2_X1 _18132_ ( .A1(_02394_ ), .A2(_02395_ ), .ZN(_02438_ ) );
INV_X1 _18133_ ( .A(\BTB.btag [0] ), .ZN(_02439_ ) );
INV_X1 _18134_ ( .A(\BTB.bindex ), .ZN(_02440_ ) );
OAI21_X1 _18135_ ( .A(_07547_ ), .B1(_02439_ ), .B2(_02440_ ), .ZN(_02441_ ) );
AOI21_X1 _18136_ ( .A(_02438_ ), .B1(_02244_ ), .B2(_02441_ ), .ZN(_02442_ ) );
MUX2_X1 _18137_ ( .A(\BTB.bsnpc_reg[0]_$_NOT__A_3_Y ), .B(\BTB.bsnpc_reg[1]_$_NOT__A_3_Y ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02443_ ) );
AND3_X1 _18138_ ( .A1(_02394_ ), .A2(_02395_ ), .A3(_02443_ ), .ZN(_02444_ ) );
OAI21_X1 _18139_ ( .A(_02437_ ), .B1(_02442_ ), .B2(_02444_ ), .ZN(_02445_ ) );
MUX2_X1 _18140_ ( .A(\BTB.bsnpc_reg[0]_$_NOT__A_3_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ), .B(\BTB.bsnpc_reg[0]_$_NOT__A_3_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02446_ ) );
NAND2_X1 _18141_ ( .A1(_02399_ ), .A2(_02446_ ), .ZN(_02447_ ) );
NAND4_X1 _18142_ ( .A1(_01658_ ), .A2(_02304_ ), .A3(_02445_ ), .A4(_02447_ ), .ZN(_02448_ ) );
OAI221_X1 _18143_ ( .A(_02448_ ), .B1(_04238_ ), .B2(_02371_ ), .C1(_02419_ ), .C2(_07547_ ), .ZN(_00795_ ) );
AND2_X1 _18144_ ( .A1(_02284_ ), .A2(_02288_ ), .ZN(_02449_ ) );
AND4_X1 _18145_ ( .A1(\BTB.pc_i [21] ), .A2(\BTB.pc_i [20] ), .A3(\BTB.pc_i [19] ), .A4(\BTB.pc_i [18] ), .ZN(_02450_ ) );
AND3_X1 _18146_ ( .A1(_02450_ ), .A2(_02257_ ), .A3(_02258_ ), .ZN(_02451_ ) );
AND2_X1 _18147_ ( .A1(_02449_ ), .A2(_02451_ ), .ZN(_02452_ ) );
NAND3_X1 _18148_ ( .A1(_02452_ ), .A2(\BTB.pc_i [27] ), .A3(\BTB.pc_i [26] ), .ZN(_02453_ ) );
XNOR2_X1 _18149_ ( .A(_02453_ ), .B(\BTB.pc_i [28] ), .ZN(_02454_ ) );
AOI22_X1 _18150_ ( .A1(_02360_ ), .A2(_02454_ ), .B1(\EXU.dnpc_o [28] ), .B2(_02269_ ), .ZN(_02455_ ) );
OAI21_X1 _18151_ ( .A(_02455_ ), .B1(_02273_ ), .B2(_02269_ ), .ZN(_02456_ ) );
MUX2_X1 _18152_ ( .A(\BTB.pc_i [28] ), .B(_02456_ ), .S(_02212_ ), .Z(_00796_ ) );
MUX2_X1 _18153_ ( .A(\BTB.bsnpc_reg[0]_$_NOT__A_4_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ), .B(\BTB.bsnpc_reg[0]_$_NOT__A_4_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02457_ ) );
NAND2_X1 _18154_ ( .A1(_02399_ ), .A2(_02457_ ), .ZN(_02458_ ) );
AND2_X1 _18155_ ( .A1(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .A2(\BTB.bsnpc_reg[1]_$_NOT__A_4_Y ), .ZN(_02459_ ) );
AOI21_X1 _18156_ ( .A(_02459_ ), .B1(_02423_ ), .B2(\BTB.bsnpc_reg[0]_$_NOT__A_4_Y ), .ZN(_02460_ ) );
NAND3_X1 _18157_ ( .A1(_02233_ ), .A2(_02240_ ), .A3(_02460_ ), .ZN(_02461_ ) );
XNOR2_X1 _18158_ ( .A(\BTB.btag [0] ), .B(\BTB.bindex ), .ZN(_02462_ ) );
OAI21_X1 _18159_ ( .A(_02461_ ), .B1(_02241_ ), .B2(_02462_ ), .ZN(_02463_ ) );
OAI211_X1 _18160_ ( .A(_02273_ ), .B(_02458_ ), .C1(_02207_ ), .C2(_02463_ ), .ZN(_02464_ ) );
OAI221_X1 _18161_ ( .A(_02464_ ), .B1(_04230_ ), .B2(_02371_ ), .C1(_02439_ ), .C2(_02419_ ), .ZN(_00797_ ) );
MUX2_X1 _18162_ ( .A(\BTB.bsnpc_reg[0]_$_NOT__A_5_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ), .B(\BTB.bsnpc_reg[0]_$_NOT__A_5_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02465_ ) );
AND3_X1 _18163_ ( .A1(_02217_ ), .A2(_02225_ ), .A3(_02465_ ), .ZN(_02466_ ) );
MUX2_X1 _18164_ ( .A(\BTB.bsnpc_reg[0]_$_NOT__A_5_Y ), .B(\BTB.bsnpc_reg[1]_$_NOT__A_5_Y ), .S(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(_02467_ ) );
AOI221_X4 _18165_ ( .A(_02466_ ), .B1(_02242_ ), .B2(\BTB.bindex ), .C1(_02335_ ), .C2(_02467_ ), .ZN(_02468_ ) );
NAND4_X1 _18166_ ( .A1(_07877_ ), .A2(_02304_ ), .A3(_01592_ ), .A4(_02468_ ), .ZN(_02469_ ) );
OAI221_X1 _18167_ ( .A(_02469_ ), .B1(_04231_ ), .B2(_02371_ ), .C1(_02419_ ), .C2(_02440_ ), .ZN(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y ) );
NOR2_X1 _18168_ ( .A1(_02277_ ), .A2(_02274_ ), .ZN(_02470_ ) );
AND2_X1 _18169_ ( .A1(_02260_ ), .A2(\BTB.pc_i [26] ), .ZN(_02471_ ) );
OAI211_X1 _18170_ ( .A(_02282_ ), .B(_02470_ ), .C1(\BTB.pc_i [27] ), .C2(_02471_ ), .ZN(_02472_ ) );
OAI211_X1 _18171_ ( .A(\BTB.pc_i [27] ), .B(_02304_ ), .C1(_02306_ ), .C2(_02300_ ), .ZN(_02473_ ) );
OAI211_X1 _18172_ ( .A(_02472_ ), .B(_02473_ ), .C1(_04246_ ), .C2(_02271_ ), .ZN(_00798_ ) );
AOI21_X1 _18173_ ( .A(_02274_ ), .B1(_02276_ ), .B2(\BTB.pc_i [26] ), .ZN(_02474_ ) );
OAI211_X1 _18174_ ( .A(_02282_ ), .B(_02474_ ), .C1(\BTB.pc_i [26] ), .C2(_02260_ ), .ZN(_02475_ ) );
OAI211_X1 _18175_ ( .A(\BTB.pc_i [26] ), .B(_02304_ ), .C1(_02306_ ), .C2(_02300_ ), .ZN(_02476_ ) );
OAI211_X1 _18176_ ( .A(_02475_ ), .B(_02476_ ), .C1(_04247_ ), .C2(_02271_ ), .ZN(_00799_ ) );
OAI21_X1 _18177_ ( .A(\BTB.pc_i [25] ), .B1(_02210_ ), .B2(_02211_ ), .ZN(_02477_ ) );
NOR2_X1 _18178_ ( .A1(_02276_ ), .A2(_02274_ ), .ZN(_02478_ ) );
AND3_X1 _18179_ ( .A1(_02293_ ), .A2(\BTB.pc_i [21] ), .A3(_02257_ ), .ZN(_02479_ ) );
AND2_X1 _18180_ ( .A1(_02479_ ), .A2(\BTB.pc_i [24] ), .ZN(_02480_ ) );
OAI211_X1 _18181_ ( .A(_02273_ ), .B(_02478_ ), .C1(\BTB.pc_i [25] ), .C2(_02480_ ), .ZN(_02481_ ) );
OAI211_X1 _18182_ ( .A(_02477_ ), .B(_02481_ ), .C1(_04248_ ), .C2(_02271_ ), .ZN(_00800_ ) );
AND2_X1 _18183_ ( .A1(_02297_ ), .A2(\BTB.pc_i [20] ), .ZN(_02482_ ) );
AND3_X1 _18184_ ( .A1(_02482_ ), .A2(\BTB.pc_i [21] ), .A3(_02257_ ), .ZN(_02483_ ) );
AOI21_X1 _18185_ ( .A(_02274_ ), .B1(_02483_ ), .B2(\BTB.pc_i [24] ), .ZN(_02484_ ) );
OAI211_X1 _18186_ ( .A(_02282_ ), .B(_02484_ ), .C1(\BTB.pc_i [24] ), .C2(_02479_ ), .ZN(_02485_ ) );
OAI211_X1 _18187_ ( .A(\BTB.pc_i [24] ), .B(_02304_ ), .C1(_02306_ ), .C2(_02300_ ), .ZN(_02486_ ) );
OAI211_X1 _18188_ ( .A(_02485_ ), .B(_02486_ ), .C1(_04249_ ), .C2(_02281_ ), .ZN(_00801_ ) );
NAND2_X1 _18189_ ( .A1(_02297_ ), .A2(\BTB.pc_i [20] ), .ZN(_02487_ ) );
NOR2_X1 _18190_ ( .A1(_02487_ ), .A2(_02283_ ), .ZN(_02488_ ) );
AOI21_X1 _18191_ ( .A(_02274_ ), .B1(_02488_ ), .B2(_02257_ ), .ZN(_02489_ ) );
AND3_X1 _18192_ ( .A1(_02293_ ), .A2(\BTB.pc_i [21] ), .A3(\BTB.pc_i [22] ), .ZN(_02490_ ) );
OAI211_X1 _18193_ ( .A(_02282_ ), .B(_02489_ ), .C1(\BTB.pc_i [23] ), .C2(_02490_ ), .ZN(_02491_ ) );
OAI211_X1 _18194_ ( .A(\BTB.pc_i [23] ), .B(_02304_ ), .C1(_02305_ ), .C2(_02300_ ), .ZN(_02492_ ) );
OAI211_X1 _18195_ ( .A(_02491_ ), .B(_02492_ ), .C1(_04253_ ), .C2(_02281_ ), .ZN(_00802_ ) );
AOI21_X1 _18196_ ( .A(_02274_ ), .B1(_02488_ ), .B2(\BTB.pc_i [22] ), .ZN(_02493_ ) );
OAI211_X1 _18197_ ( .A(_02282_ ), .B(_02493_ ), .C1(\BTB.pc_i [22] ), .C2(_02294_ ), .ZN(_02494_ ) );
OAI211_X1 _18198_ ( .A(\BTB.pc_i [22] ), .B(_02303_ ), .C1(_02305_ ), .C2(_02300_ ), .ZN(_02495_ ) );
OAI211_X1 _18199_ ( .A(_02494_ ), .B(_02495_ ), .C1(_04254_ ), .C2(_02281_ ), .ZN(_00803_ ) );
MUX2_X1 _18200_ ( .A(\BTB.prepc_tag_i [31] ), .B(\BTB.pc_i [31] ), .S(_02071_ ), .Z(_00804_ ) );
MUX2_X1 _18201_ ( .A(\BTB.prepc_tag_i [30] ), .B(\BTB.pc_i [30] ), .S(_02071_ ), .Z(_00805_ ) );
MUX2_X1 _18202_ ( .A(\BTB.prepc_tag_i [21] ), .B(\BTB.pc_i [21] ), .S(_02071_ ), .Z(_00806_ ) );
MUX2_X1 _18203_ ( .A(\BTB.prepc_tag_i [20] ), .B(\BTB.pc_i [20] ), .S(_02071_ ), .Z(_00807_ ) );
MUX2_X1 _18204_ ( .A(\BTB.prepc_tag_i [19] ), .B(\BTB.pc_i [19] ), .S(_02071_ ), .Z(_00808_ ) );
MUX2_X1 _18205_ ( .A(\BTB.prepc_tag_i [18] ), .B(\BTB.pc_i [18] ), .S(_02071_ ), .Z(_00809_ ) );
BUF_X4 _18206_ ( .A(_01595_ ), .Z(_02496_ ) );
MUX2_X1 _18207_ ( .A(\BTB.prepc_tag_i [17] ), .B(\BTB.pc_i [17] ), .S(_02496_ ), .Z(_00810_ ) );
MUX2_X1 _18208_ ( .A(\BTB.prepc_tag_i [16] ), .B(\BTB.pc_i [16] ), .S(_02496_ ), .Z(_00811_ ) );
MUX2_X1 _18209_ ( .A(\BTB.btag_pre [12] ), .B(\BTB.btag [12] ), .S(_02496_ ), .Z(_00812_ ) );
MUX2_X1 _18210_ ( .A(\BTB.btag_pre [11] ), .B(\BTB.btag [11] ), .S(_02496_ ), .Z(_00813_ ) );
MUX2_X1 _18211_ ( .A(\BTB.btag_pre [10] ), .B(\BTB.btag [10] ), .S(_02496_ ), .Z(_00814_ ) );
MUX2_X1 _18212_ ( .A(\BTB.btag_pre [9] ), .B(\BTB.btag [9] ), .S(_02496_ ), .Z(_00815_ ) );
MUX2_X1 _18213_ ( .A(\BTB.prepc_tag_i [29] ), .B(\BTB.pc_i [29] ), .S(_02496_ ), .Z(_00816_ ) );
MUX2_X1 _18214_ ( .A(\BTB.btag_pre [8] ), .B(\BTB.btag [8] ), .S(_02496_ ), .Z(_00817_ ) );
MUX2_X1 _18215_ ( .A(\BTB.btag_pre [7] ), .B(\BTB.btag [7] ), .S(_02496_ ), .Z(_00818_ ) );
MUX2_X1 _18216_ ( .A(\BTB.btag_pre [6] ), .B(\BTB.btag [6] ), .S(_02496_ ), .Z(_00819_ ) );
BUF_X4 _18217_ ( .A(_01595_ ), .Z(_02497_ ) );
MUX2_X1 _18218_ ( .A(\BTB.btag_pre [5] ), .B(\BTB.btag [5] ), .S(_02497_ ), .Z(_00820_ ) );
MUX2_X1 _18219_ ( .A(\BTB.btag_pre [4] ), .B(\BTB.btag [4] ), .S(_02497_ ), .Z(_00821_ ) );
MUX2_X1 _18220_ ( .A(\BTB.btag_pre [3] ), .B(\BTB.btag [3] ), .S(_02497_ ), .Z(_00822_ ) );
MUX2_X1 _18221_ ( .A(\BTB.btag_pre [2] ), .B(\BTB.btag [2] ), .S(_02497_ ), .Z(_00823_ ) );
MUX2_X1 _18222_ ( .A(\BTB.btag_pre [1] ), .B(\BTB.btag [1] ), .S(_02497_ ), .Z(_00824_ ) );
MUX2_X1 _18223_ ( .A(\BTB.btag_pre [0] ), .B(\BTB.btag [0] ), .S(_02497_ ), .Z(_00825_ ) );
MUX2_X1 _18224_ ( .A(\BTB.bindex_pre ), .B(\BTB.bindex ), .S(_02497_ ), .Z(_00826_ ) );
MUX2_X1 _18225_ ( .A(\BTB.prepc_tag_i [28] ), .B(\BTB.pc_i [28] ), .S(_02497_ ), .Z(_00827_ ) );
MUX2_X1 _18226_ ( .A(\BTB.prepc_tag_i [1] ), .B(\BTB.pc_i [1] ), .S(_02497_ ), .Z(_00828_ ) );
MUX2_X1 _18227_ ( .A(\BTB.prepc_tag_i [0] ), .B(\BTB.pc_i [0] ), .S(_02497_ ), .Z(_00829_ ) );
MUX2_X1 _18228_ ( .A(\BTB.prepc_tag_i [27] ), .B(\BTB.pc_i [27] ), .S(_02317_ ), .Z(_00830_ ) );
MUX2_X1 _18229_ ( .A(\BTB.prepc_tag_i [26] ), .B(\BTB.pc_i [26] ), .S(_02317_ ), .Z(_00831_ ) );
MUX2_X1 _18230_ ( .A(\BTB.prepc_tag_i [25] ), .B(\BTB.pc_i [25] ), .S(_02317_ ), .Z(_00832_ ) );
MUX2_X1 _18231_ ( .A(\BTB.prepc_tag_i [24] ), .B(\BTB.pc_i [24] ), .S(_02317_ ), .Z(_00833_ ) );
MUX2_X1 _18232_ ( .A(\BTB.prepc_tag_i [23] ), .B(\BTB.pc_i [23] ), .S(_02317_ ), .Z(_00834_ ) );
MUX2_X1 _18233_ ( .A(\BTB.prepc_tag_i [22] ), .B(\BTB.pc_i [22] ), .S(_02317_ ), .Z(_00835_ ) );
INV_X1 _18234_ ( .A(\LSU.axi_state [2] ), .ZN(_02498_ ) );
CLKBUF_X2 _18235_ ( .A(_02498_ ), .Z(_02499_ ) );
INV_X1 _18236_ ( .A(_04390_ ), .ZN(_02500_ ) );
BUF_X4 _18237_ ( .A(_02500_ ), .Z(_02501_ ) );
AND3_X1 _18238_ ( .A1(_04653_ ), .A2(_02499_ ), .A3(_02501_ ), .ZN(_02502_ ) );
INV_X1 _18239_ ( .A(\LSU.ls_axi_arvalid_$_SDFFE_PP0P__Q_D ), .ZN(_02503_ ) );
OAI21_X1 _18240_ ( .A(\LSU.ls_axi_rready ), .B1(_04055_ ), .B2(\Xbar.state [2] ), .ZN(_02504_ ) );
OAI21_X1 _18241_ ( .A(_02503_ ), .B1(_07542_ ), .B2(_02504_ ), .ZN(_02505_ ) );
AOI21_X1 _18242_ ( .A(_07929_ ), .B1(_04287_ ), .B2(_04330_ ), .ZN(_02506_ ) );
AND2_X1 _18243_ ( .A1(_02506_ ), .A2(_06006_ ), .ZN(_02507_ ) );
MUX2_X1 _18244_ ( .A(\LSU.axi_state [2] ), .B(_02507_ ), .S(\LSU.axi_state [0] ), .Z(_02508_ ) );
AND2_X1 _18245_ ( .A1(_02508_ ), .A2(_03805_ ), .ZN(_02509_ ) );
AND2_X2 _18246_ ( .A1(_02505_ ), .A2(_02509_ ), .ZN(_02510_ ) );
BUF_X4 _18247_ ( .A(_02510_ ), .Z(_02511_ ) );
MUX2_X1 _18248_ ( .A(\LSU.ls_axi_araddr [31] ), .B(_02502_ ), .S(_02511_ ), .Z(_00837_ ) );
AND3_X1 _18249_ ( .A1(_05089_ ), .A2(_02499_ ), .A3(_02501_ ), .ZN(_02512_ ) );
MUX2_X1 _18250_ ( .A(\LSU.ls_axi_araddr [30] ), .B(_02512_ ), .S(_02511_ ), .Z(_00838_ ) );
AND3_X1 _18251_ ( .A1(_05114_ ), .A2(_02499_ ), .A3(_02501_ ), .ZN(_02513_ ) );
MUX2_X1 _18252_ ( .A(\LSU.ls_axi_araddr [21] ), .B(_02513_ ), .S(_02511_ ), .Z(_00839_ ) );
AND3_X1 _18253_ ( .A1(_05133_ ), .A2(_02499_ ), .A3(_02501_ ), .ZN(_02514_ ) );
MUX2_X1 _18254_ ( .A(\LSU.ls_axi_araddr [20] ), .B(_02514_ ), .S(_02511_ ), .Z(_00840_ ) );
AND3_X1 _18255_ ( .A1(_05147_ ), .A2(_02499_ ), .A3(_02501_ ), .ZN(_02515_ ) );
MUX2_X1 _18256_ ( .A(\LSU.ls_axi_araddr [19] ), .B(_02515_ ), .S(_02511_ ), .Z(_00841_ ) );
AND3_X1 _18257_ ( .A1(_05157_ ), .A2(_02499_ ), .A3(_02501_ ), .ZN(_02516_ ) );
MUX2_X1 _18258_ ( .A(\LSU.ls_axi_araddr [18] ), .B(_02516_ ), .S(_02511_ ), .Z(_00842_ ) );
AND3_X1 _18259_ ( .A1(_05178_ ), .A2(_02499_ ), .A3(_02501_ ), .ZN(_02517_ ) );
MUX2_X1 _18260_ ( .A(\LSU.ls_axi_araddr [17] ), .B(_02517_ ), .S(_02511_ ), .Z(_00843_ ) );
CLKBUF_X2 _18261_ ( .A(_02500_ ), .Z(_02518_ ) );
AND3_X1 _18262_ ( .A1(_05187_ ), .A2(_02499_ ), .A3(_02518_ ), .ZN(_02519_ ) );
MUX2_X1 _18263_ ( .A(\LSU.ls_axi_araddr [16] ), .B(_02519_ ), .S(_02511_ ), .Z(_00844_ ) );
AND3_X1 _18264_ ( .A1(_05198_ ), .A2(_02499_ ), .A3(_02518_ ), .ZN(_02520_ ) );
MUX2_X1 _18265_ ( .A(\LSU.ls_axi_araddr [15] ), .B(_02520_ ), .S(_02511_ ), .Z(_00845_ ) );
AND3_X1 _18266_ ( .A1(_05209_ ), .A2(_02499_ ), .A3(_02518_ ), .ZN(_02521_ ) );
MUX2_X1 _18267_ ( .A(\LSU.ls_axi_araddr [14] ), .B(_02521_ ), .S(_02511_ ), .Z(_00846_ ) );
CLKBUF_X2 _18268_ ( .A(_02498_ ), .Z(_02522_ ) );
AND3_X1 _18269_ ( .A1(_05228_ ), .A2(_02522_ ), .A3(_02518_ ), .ZN(_02523_ ) );
BUF_X4 _18270_ ( .A(_02510_ ), .Z(_02524_ ) );
MUX2_X1 _18271_ ( .A(\LSU.ls_axi_araddr [13] ), .B(_02523_ ), .S(_02524_ ), .Z(_00847_ ) );
AND3_X1 _18272_ ( .A1(_05236_ ), .A2(_02522_ ), .A3(_02518_ ), .ZN(_02525_ ) );
MUX2_X1 _18273_ ( .A(\LSU.ls_axi_araddr [12] ), .B(_02525_ ), .S(_02524_ ), .Z(_00848_ ) );
AND3_X1 _18274_ ( .A1(_05250_ ), .A2(_02522_ ), .A3(_02518_ ), .ZN(_02526_ ) );
MUX2_X1 _18275_ ( .A(\LSU.ls_axi_araddr [29] ), .B(_02526_ ), .S(_02524_ ), .Z(_00849_ ) );
AND3_X1 _18276_ ( .A1(_05258_ ), .A2(_02522_ ), .A3(_02518_ ), .ZN(_02527_ ) );
MUX2_X1 _18277_ ( .A(\LSU.ls_axi_araddr [11] ), .B(_02527_ ), .S(_02524_ ), .Z(_00850_ ) );
AND3_X1 _18278_ ( .A1(_05269_ ), .A2(_02522_ ), .A3(_02518_ ), .ZN(_02528_ ) );
MUX2_X1 _18279_ ( .A(\LSU.ls_axi_araddr [10] ), .B(_02528_ ), .S(_02524_ ), .Z(_00851_ ) );
AND3_X1 _18280_ ( .A1(_05280_ ), .A2(_02522_ ), .A3(_02518_ ), .ZN(_02529_ ) );
MUX2_X1 _18281_ ( .A(\LSU.ls_axi_araddr [9] ), .B(_02529_ ), .S(_02524_ ), .Z(_00852_ ) );
AND3_X1 _18282_ ( .A1(_05295_ ), .A2(_02522_ ), .A3(_02518_ ), .ZN(_02530_ ) );
MUX2_X1 _18283_ ( .A(\LSU.ls_axi_araddr [8] ), .B(_02530_ ), .S(_02524_ ), .Z(_00853_ ) );
CLKBUF_X2 _18284_ ( .A(_02500_ ), .Z(_02531_ ) );
AND3_X1 _18285_ ( .A1(_05303_ ), .A2(_02522_ ), .A3(_02531_ ), .ZN(_02532_ ) );
MUX2_X1 _18286_ ( .A(\LSU.ls_axi_araddr [7] ), .B(_02532_ ), .S(_02524_ ), .Z(_00854_ ) );
AND3_X1 _18287_ ( .A1(_05306_ ), .A2(_02522_ ), .A3(_02531_ ), .ZN(_02533_ ) );
MUX2_X1 _18288_ ( .A(\LSU.ls_axi_araddr [6] ), .B(_02533_ ), .S(_02524_ ), .Z(_00855_ ) );
AND3_X1 _18289_ ( .A1(_05313_ ), .A2(_02522_ ), .A3(_02531_ ), .ZN(_02534_ ) );
MUX2_X1 _18290_ ( .A(\LSU.ls_axi_araddr [5] ), .B(_02534_ ), .S(_02524_ ), .Z(_00856_ ) );
CLKBUF_X2 _18291_ ( .A(_02498_ ), .Z(_02535_ ) );
AND3_X1 _18292_ ( .A1(_05329_ ), .A2(_02535_ ), .A3(_02531_ ), .ZN(_02536_ ) );
BUF_X4 _18293_ ( .A(_02510_ ), .Z(_02537_ ) );
MUX2_X1 _18294_ ( .A(\LSU.ls_axi_araddr [4] ), .B(_02536_ ), .S(_02537_ ), .Z(_00857_ ) );
AND3_X1 _18295_ ( .A1(_05338_ ), .A2(_02535_ ), .A3(_02531_ ), .ZN(_02538_ ) );
MUX2_X1 _18296_ ( .A(\LSU.ls_axi_araddr [3] ), .B(_02538_ ), .S(_02537_ ), .Z(_00858_ ) );
AND3_X1 _18297_ ( .A1(_05343_ ), .A2(_02535_ ), .A3(_02531_ ), .ZN(_02539_ ) );
MUX2_X1 _18298_ ( .A(\LSU.ls_axi_araddr [2] ), .B(_02539_ ), .S(_02537_ ), .Z(_00859_ ) );
AND3_X1 _18299_ ( .A1(_05345_ ), .A2(_02535_ ), .A3(_02531_ ), .ZN(_02540_ ) );
MUX2_X1 _18300_ ( .A(\LSU.ls_axi_araddr [28] ), .B(_02540_ ), .S(_02537_ ), .Z(_00860_ ) );
AND3_X1 _18301_ ( .A1(_05353_ ), .A2(_02535_ ), .A3(_02531_ ), .ZN(_02541_ ) );
MUX2_X1 _18302_ ( .A(\LSU.ls_axi_araddr [1] ), .B(_02541_ ), .S(_02537_ ), .Z(_00861_ ) );
AND3_X1 _18303_ ( .A1(_05359_ ), .A2(_02535_ ), .A3(_02531_ ), .ZN(_02542_ ) );
MUX2_X1 _18304_ ( .A(\LSU.ls_axi_araddr [0] ), .B(_02542_ ), .S(_02537_ ), .Z(_00862_ ) );
AND3_X1 _18305_ ( .A1(_05370_ ), .A2(_02535_ ), .A3(_02531_ ), .ZN(_02543_ ) );
MUX2_X1 _18306_ ( .A(\LSU.ls_axi_araddr [27] ), .B(_02543_ ), .S(_02537_ ), .Z(_00863_ ) );
AND3_X1 _18307_ ( .A1(_05382_ ), .A2(_02535_ ), .A3(_02500_ ), .ZN(_02544_ ) );
MUX2_X1 _18308_ ( .A(\LSU.ls_axi_araddr [26] ), .B(_02544_ ), .S(_02537_ ), .Z(_00864_ ) );
BUF_X2 _18309_ ( .A(_04390_ ), .Z(_02545_ ) );
NOR3_X1 _18310_ ( .A1(_05394_ ), .A2(\LSU.axi_state [2] ), .A3(_02545_ ), .ZN(_02546_ ) );
MUX2_X1 _18311_ ( .A(\LSU.ls_axi_araddr [25] ), .B(_02546_ ), .S(_02537_ ), .Z(_00865_ ) );
AND3_X1 _18312_ ( .A1(_05396_ ), .A2(_02535_ ), .A3(_02500_ ), .ZN(_02547_ ) );
MUX2_X1 _18313_ ( .A(\LSU.ls_axi_araddr [24] ), .B(_02547_ ), .S(_02537_ ), .Z(_00866_ ) );
AND3_X1 _18314_ ( .A1(_05409_ ), .A2(_02535_ ), .A3(_02500_ ), .ZN(_02548_ ) );
MUX2_X1 _18315_ ( .A(\LSU.ls_axi_araddr [23] ), .B(_02548_ ), .S(_02510_ ), .Z(_00867_ ) );
AND3_X1 _18316_ ( .A1(_05416_ ), .A2(_02498_ ), .A3(_02500_ ), .ZN(_02549_ ) );
MUX2_X1 _18317_ ( .A(\LSU.ls_axi_araddr [22] ), .B(_02549_ ), .S(_02510_ ), .Z(_00868_ ) );
INV_X1 _18318_ ( .A(\LSU.axi_state [1] ), .ZN(_02550_ ) );
BUF_X4 _18319_ ( .A(_02550_ ), .Z(_02551_ ) );
BUF_X4 _18320_ ( .A(_02501_ ), .Z(_02552_ ) );
AND2_X1 _18321_ ( .A1(_02506_ ), .A2(_04384_ ), .ZN(_02553_ ) );
INV_X1 _18322_ ( .A(\LSU.axi_state [0] ), .ZN(_02554_ ) );
OAI21_X1 _18323_ ( .A(_03798_ ), .B1(_02553_ ), .B2(_02554_ ), .ZN(_02555_ ) );
AND3_X1 _18324_ ( .A1(io_master_bready ), .A2(\LSU.axi_state [1] ), .A3(io_master_bvalid ), .ZN(_02556_ ) );
NOR2_X1 _18325_ ( .A1(_02554_ ), .A2(\LSU.axi_state [1] ), .ZN(_02557_ ) );
NOR2_X1 _18326_ ( .A1(_02556_ ), .A2(_02557_ ), .ZN(_02558_ ) );
NOR2_X2 _18327_ ( .A1(_02555_ ), .A2(_02558_ ), .ZN(_02559_ ) );
BUF_X4 _18328_ ( .A(_02559_ ), .Z(_02560_ ) );
NAND4_X1 _18329_ ( .A1(_04653_ ), .A2(_02551_ ), .A3(_02552_ ), .A4(_02560_ ), .ZN(_02561_ ) );
INV_X1 _18330_ ( .A(\LSU.ls_axi_awaddr [31] ), .ZN(_02562_ ) );
BUF_X4 _18331_ ( .A(_02559_ ), .Z(_02563_ ) );
OAI21_X1 _18332_ ( .A(_02561_ ), .B1(_02562_ ), .B2(_02563_ ), .ZN(_00870_ ) );
NAND4_X1 _18333_ ( .A1(_05089_ ), .A2(_02551_ ), .A3(_02552_ ), .A4(_02560_ ), .ZN(_02564_ ) );
INV_X1 _18334_ ( .A(\LSU.ls_axi_awaddr [30] ), .ZN(_02565_ ) );
OAI21_X1 _18335_ ( .A(_02564_ ), .B1(_02565_ ), .B2(_02563_ ), .ZN(_00871_ ) );
NAND4_X1 _18336_ ( .A1(_05114_ ), .A2(_02551_ ), .A3(_02552_ ), .A4(_02560_ ), .ZN(_02566_ ) );
INV_X1 _18337_ ( .A(\LSU.ls_axi_awaddr [21] ), .ZN(_02567_ ) );
OAI21_X1 _18338_ ( .A(_02566_ ), .B1(_02567_ ), .B2(_02563_ ), .ZN(_00872_ ) );
NAND4_X1 _18339_ ( .A1(_05133_ ), .A2(_02551_ ), .A3(_02552_ ), .A4(_02560_ ), .ZN(_02568_ ) );
INV_X1 _18340_ ( .A(\LSU.ls_axi_awaddr [20] ), .ZN(_02569_ ) );
OAI21_X1 _18341_ ( .A(_02568_ ), .B1(_02569_ ), .B2(_02563_ ), .ZN(_00873_ ) );
NAND4_X1 _18342_ ( .A1(_05147_ ), .A2(_02551_ ), .A3(_02552_ ), .A4(_02560_ ), .ZN(_02570_ ) );
INV_X1 _18343_ ( .A(\LSU.ls_axi_awaddr [19] ), .ZN(_02571_ ) );
OAI21_X1 _18344_ ( .A(_02570_ ), .B1(_02571_ ), .B2(_02563_ ), .ZN(_00874_ ) );
NAND4_X1 _18345_ ( .A1(_05157_ ), .A2(_02551_ ), .A3(_02552_ ), .A4(_02560_ ), .ZN(_02572_ ) );
INV_X1 _18346_ ( .A(\LSU.ls_axi_awaddr [18] ), .ZN(_02573_ ) );
OAI21_X1 _18347_ ( .A(_02572_ ), .B1(_02573_ ), .B2(_02563_ ), .ZN(_00875_ ) );
NAND4_X1 _18348_ ( .A1(_05178_ ), .A2(_02551_ ), .A3(_02552_ ), .A4(_02560_ ), .ZN(_02574_ ) );
INV_X1 _18349_ ( .A(\LSU.ls_axi_awaddr [17] ), .ZN(_02575_ ) );
OAI21_X1 _18350_ ( .A(_02574_ ), .B1(_02575_ ), .B2(_02563_ ), .ZN(_00876_ ) );
NAND4_X1 _18351_ ( .A1(_05187_ ), .A2(_02551_ ), .A3(_02552_ ), .A4(_02560_ ), .ZN(_02576_ ) );
INV_X1 _18352_ ( .A(\LSU.ls_axi_awaddr [16] ), .ZN(_02577_ ) );
OAI21_X1 _18353_ ( .A(_02576_ ), .B1(_02577_ ), .B2(_02563_ ), .ZN(_00877_ ) );
BUF_X4 _18354_ ( .A(_02559_ ), .Z(_02578_ ) );
NAND4_X1 _18355_ ( .A1(_05198_ ), .A2(_02551_ ), .A3(_02552_ ), .A4(_02578_ ), .ZN(_02579_ ) );
INV_X1 _18356_ ( .A(\LSU.ls_axi_awaddr [15] ), .ZN(_02580_ ) );
OAI21_X1 _18357_ ( .A(_02579_ ), .B1(_02580_ ), .B2(_02563_ ), .ZN(_00878_ ) );
BUF_X4 _18358_ ( .A(_02501_ ), .Z(_02581_ ) );
NAND4_X1 _18359_ ( .A1(_05209_ ), .A2(_02551_ ), .A3(_02581_ ), .A4(_02578_ ), .ZN(_02582_ ) );
INV_X1 _18360_ ( .A(\LSU.ls_axi_awaddr [14] ), .ZN(_02583_ ) );
OAI21_X1 _18361_ ( .A(_02582_ ), .B1(_02583_ ), .B2(_02563_ ), .ZN(_00879_ ) );
BUF_X4 _18362_ ( .A(_02550_ ), .Z(_02584_ ) );
NAND4_X1 _18363_ ( .A1(_05228_ ), .A2(_02584_ ), .A3(_02581_ ), .A4(_02578_ ), .ZN(_02585_ ) );
INV_X1 _18364_ ( .A(\LSU.ls_axi_awaddr [13] ), .ZN(_02586_ ) );
BUF_X4 _18365_ ( .A(_02559_ ), .Z(_02587_ ) );
OAI21_X1 _18366_ ( .A(_02585_ ), .B1(_02586_ ), .B2(_02587_ ), .ZN(_00880_ ) );
NAND4_X1 _18367_ ( .A1(_05236_ ), .A2(_02584_ ), .A3(_02581_ ), .A4(_02578_ ), .ZN(_02588_ ) );
INV_X1 _18368_ ( .A(\LSU.ls_axi_awaddr [12] ), .ZN(_02589_ ) );
OAI21_X1 _18369_ ( .A(_02588_ ), .B1(_02589_ ), .B2(_02587_ ), .ZN(_00881_ ) );
NAND4_X1 _18370_ ( .A1(_05250_ ), .A2(_02584_ ), .A3(_02581_ ), .A4(_02578_ ), .ZN(_02590_ ) );
INV_X1 _18371_ ( .A(\LSU.ls_axi_awaddr [29] ), .ZN(_02591_ ) );
OAI21_X1 _18372_ ( .A(_02590_ ), .B1(_02591_ ), .B2(_02587_ ), .ZN(_00882_ ) );
NAND4_X1 _18373_ ( .A1(_05258_ ), .A2(_02584_ ), .A3(_02581_ ), .A4(_02578_ ), .ZN(_02592_ ) );
INV_X1 _18374_ ( .A(\LSU.ls_axi_awaddr [11] ), .ZN(_02593_ ) );
OAI21_X1 _18375_ ( .A(_02592_ ), .B1(_02593_ ), .B2(_02587_ ), .ZN(_00883_ ) );
NAND4_X1 _18376_ ( .A1(_05269_ ), .A2(_02584_ ), .A3(_02581_ ), .A4(_02578_ ), .ZN(_02594_ ) );
INV_X1 _18377_ ( .A(\LSU.ls_axi_awaddr [10] ), .ZN(_02595_ ) );
OAI21_X1 _18378_ ( .A(_02594_ ), .B1(_02595_ ), .B2(_02587_ ), .ZN(_00884_ ) );
NAND4_X1 _18379_ ( .A1(_05280_ ), .A2(_02584_ ), .A3(_02581_ ), .A4(_02578_ ), .ZN(_02596_ ) );
INV_X1 _18380_ ( .A(\LSU.ls_axi_awaddr [9] ), .ZN(_02597_ ) );
OAI21_X1 _18381_ ( .A(_02596_ ), .B1(_02597_ ), .B2(_02587_ ), .ZN(_00885_ ) );
NAND4_X1 _18382_ ( .A1(_05295_ ), .A2(_02584_ ), .A3(_02581_ ), .A4(_02578_ ), .ZN(_02598_ ) );
INV_X1 _18383_ ( .A(\LSU.ls_axi_awaddr [8] ), .ZN(_02599_ ) );
OAI21_X1 _18384_ ( .A(_02598_ ), .B1(_02599_ ), .B2(_02587_ ), .ZN(_00886_ ) );
NAND4_X1 _18385_ ( .A1(_05303_ ), .A2(_02584_ ), .A3(_02581_ ), .A4(_02578_ ), .ZN(_02600_ ) );
INV_X1 _18386_ ( .A(\LSU.ls_axi_awaddr [7] ), .ZN(_02601_ ) );
OAI21_X1 _18387_ ( .A(_02600_ ), .B1(_02601_ ), .B2(_02587_ ), .ZN(_00887_ ) );
BUF_X4 _18388_ ( .A(_02559_ ), .Z(_02602_ ) );
NAND4_X1 _18389_ ( .A1(_05306_ ), .A2(_02584_ ), .A3(_02581_ ), .A4(_02602_ ), .ZN(_02603_ ) );
INV_X1 _18390_ ( .A(\LSU.ls_axi_awaddr [6] ), .ZN(_02604_ ) );
OAI21_X1 _18391_ ( .A(_02603_ ), .B1(_02604_ ), .B2(_02587_ ), .ZN(_00888_ ) );
BUF_X4 _18392_ ( .A(_02501_ ), .Z(_02605_ ) );
NAND4_X1 _18393_ ( .A1(_05313_ ), .A2(_02584_ ), .A3(_02605_ ), .A4(_02602_ ), .ZN(_02606_ ) );
INV_X1 _18394_ ( .A(\LSU.ls_axi_awaddr [5] ), .ZN(_02607_ ) );
OAI21_X1 _18395_ ( .A(_02606_ ), .B1(_02607_ ), .B2(_02587_ ), .ZN(_00889_ ) );
BUF_X2 _18396_ ( .A(_02550_ ), .Z(_02608_ ) );
NAND4_X1 _18397_ ( .A1(_05329_ ), .A2(_02608_ ), .A3(_02605_ ), .A4(_02602_ ), .ZN(_02609_ ) );
INV_X1 _18398_ ( .A(\LSU.ls_axi_awaddr [4] ), .ZN(_02610_ ) );
BUF_X4 _18399_ ( .A(_02559_ ), .Z(_02611_ ) );
OAI21_X1 _18400_ ( .A(_02609_ ), .B1(_02610_ ), .B2(_02611_ ), .ZN(_00890_ ) );
NAND4_X1 _18401_ ( .A1(_05338_ ), .A2(_02608_ ), .A3(_02605_ ), .A4(_02602_ ), .ZN(_02612_ ) );
INV_X1 _18402_ ( .A(\LSU.ls_axi_awaddr [3] ), .ZN(_02613_ ) );
OAI21_X1 _18403_ ( .A(_02612_ ), .B1(_02613_ ), .B2(_02611_ ), .ZN(_00891_ ) );
NAND4_X1 _18404_ ( .A1(_05343_ ), .A2(_02608_ ), .A3(_02605_ ), .A4(_02602_ ), .ZN(_02614_ ) );
INV_X1 _18405_ ( .A(\LSU.ls_axi_awaddr [2] ), .ZN(_02615_ ) );
OAI21_X1 _18406_ ( .A(_02614_ ), .B1(_02615_ ), .B2(_02611_ ), .ZN(_00892_ ) );
NAND4_X1 _18407_ ( .A1(_05345_ ), .A2(_02608_ ), .A3(_02605_ ), .A4(_02602_ ), .ZN(_02616_ ) );
INV_X1 _18408_ ( .A(\LSU.ls_axi_awaddr [28] ), .ZN(_02617_ ) );
OAI21_X1 _18409_ ( .A(_02616_ ), .B1(_02617_ ), .B2(_02611_ ), .ZN(_00893_ ) );
AND2_X2 _18410_ ( .A1(_05352_ ), .A2(_02500_ ), .ZN(_02618_ ) );
INV_X1 _18411_ ( .A(_02618_ ), .ZN(_02619_ ) );
NAND2_X1 _18412_ ( .A1(_02559_ ), .A2(_02550_ ), .ZN(_02620_ ) );
INV_X1 _18413_ ( .A(\LSU.ls_axi_awaddr [1] ), .ZN(_02621_ ) );
OAI22_X1 _18414_ ( .A1(_02619_ ), .A2(_02620_ ), .B1(_02621_ ), .B2(_02560_ ), .ZN(_00894_ ) );
AND2_X2 _18415_ ( .A1(_05359_ ), .A2(_02500_ ), .ZN(_02622_ ) );
INV_X1 _18416_ ( .A(_02622_ ), .ZN(_02623_ ) );
INV_X1 _18417_ ( .A(\LSU.ls_axi_awaddr [0] ), .ZN(_02624_ ) );
OAI22_X1 _18418_ ( .A1(_02623_ ), .A2(_02620_ ), .B1(_02624_ ), .B2(_02560_ ), .ZN(_00895_ ) );
NAND4_X1 _18419_ ( .A1(_05370_ ), .A2(_02608_ ), .A3(_02605_ ), .A4(_02602_ ), .ZN(_02625_ ) );
INV_X1 _18420_ ( .A(\LSU.ls_axi_awaddr [27] ), .ZN(_02626_ ) );
OAI21_X1 _18421_ ( .A(_02625_ ), .B1(_02626_ ), .B2(_02611_ ), .ZN(_00896_ ) );
NAND4_X1 _18422_ ( .A1(_05382_ ), .A2(_02608_ ), .A3(_02605_ ), .A4(_02602_ ), .ZN(_02627_ ) );
INV_X1 _18423_ ( .A(\LSU.ls_axi_awaddr [26] ), .ZN(_02628_ ) );
OAI21_X1 _18424_ ( .A(_02627_ ), .B1(_02628_ ), .B2(_02611_ ), .ZN(_00897_ ) );
OR3_X1 _18425_ ( .A1(_05394_ ), .A2(_02545_ ), .A3(_02620_ ), .ZN(_02629_ ) );
INV_X1 _18426_ ( .A(\LSU.ls_axi_awaddr [25] ), .ZN(_02630_ ) );
OAI21_X1 _18427_ ( .A(_02629_ ), .B1(_02630_ ), .B2(_02611_ ), .ZN(_00898_ ) );
NAND4_X1 _18428_ ( .A1(_05396_ ), .A2(_02608_ ), .A3(_02605_ ), .A4(_02602_ ), .ZN(_02631_ ) );
INV_X1 _18429_ ( .A(\LSU.ls_axi_awaddr [24] ), .ZN(_02632_ ) );
OAI21_X1 _18430_ ( .A(_02631_ ), .B1(_02632_ ), .B2(_02611_ ), .ZN(_00899_ ) );
NAND4_X1 _18431_ ( .A1(_05409_ ), .A2(_02608_ ), .A3(_02605_ ), .A4(_02602_ ), .ZN(_02633_ ) );
INV_X1 _18432_ ( .A(\LSU.ls_axi_awaddr [23] ), .ZN(_02634_ ) );
OAI21_X1 _18433_ ( .A(_02633_ ), .B1(_02634_ ), .B2(_02611_ ), .ZN(_00900_ ) );
NAND4_X1 _18434_ ( .A1(_05416_ ), .A2(_02608_ ), .A3(_02605_ ), .A4(_02559_ ), .ZN(_02635_ ) );
INV_X1 _18435_ ( .A(\LSU.ls_axi_awaddr [22] ), .ZN(_02636_ ) );
OAI21_X1 _18436_ ( .A(_02635_ ), .B1(_02636_ ), .B2(_02611_ ), .ZN(_00901_ ) );
INV_X1 _18437_ ( .A(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ), .ZN(_02637_ ) );
AND4_X1 _18438_ ( .A1(_02637_ ), .A2(io_master_bready ), .A3(_03805_ ), .A4(io_master_bvalid ), .ZN(_02638_ ) );
NOR2_X1 _18439_ ( .A1(_04058_ ), .A2(\LSU.ls_axi_awvalid_$_NOT__A_Y ), .ZN(io_master_awvalid ) );
AND2_X1 _18440_ ( .A1(io_master_awvalid ), .A2(io_master_awready ), .ZN(_02639_ ) );
NOR2_X1 _18441_ ( .A1(_04105_ ), .A2(\LSU.ls_axi_wvalid_$_NOT__A_Y ), .ZN(io_master_wvalid ) );
AND3_X1 _18442_ ( .A1(_02639_ ), .A2(io_master_wready ), .A3(io_master_wvalid ), .ZN(_02640_ ) );
NAND3_X1 _18443_ ( .A1(_02640_ ), .A2(_02637_ ), .A3(_03806_ ), .ZN(_02641_ ) );
AOI21_X1 _18444_ ( .A(_02638_ ), .B1(_02641_ ), .B2(_04379_ ), .ZN(_00903_ ) );
NAND3_X1 _18445_ ( .A1(_07887_ ), .A2(_07543_ ), .A3(_07888_ ), .ZN(_02642_ ) );
INV_X1 _18446_ ( .A(\LSU.ls_axi_arvalid ), .ZN(_02643_ ) );
NOR4_X1 _18447_ ( .A1(_02642_ ), .A2(_02643_ ), .A3(\LSU.ls_axi_arvalid_$_SDFFE_PP0P__Q_D ), .A4(fanout_net_11 ), .ZN(_02644_ ) );
OR2_X1 _18448_ ( .A1(_02644_ ), .A2(\LSU.ls_axi_rready ), .ZN(_02645_ ) );
NOR2_X1 _18449_ ( .A1(_07542_ ), .A2(_02504_ ), .ZN(_02646_ ) );
BUF_X4 _18450_ ( .A(_02646_ ), .Z(_02647_ ) );
NAND3_X1 _18451_ ( .A1(_02647_ ), .A2(_02503_ ), .A3(_03833_ ), .ZN(_02648_ ) );
AND2_X1 _18452_ ( .A1(_02645_ ), .A2(_02648_ ), .ZN(_00904_ ) );
BUF_X4 _18453_ ( .A(_02618_ ), .Z(_02649_ ) );
BUF_X4 _18454_ ( .A(_02622_ ), .Z(_02650_ ) );
NAND3_X1 _18455_ ( .A1(_02649_ ), .A2(\EXU.r2_i [7] ), .A3(_02650_ ), .ZN(_02651_ ) );
NOR2_X1 _18456_ ( .A1(_02618_ ), .A2(_02623_ ), .ZN(_02652_ ) );
INV_X1 _18457_ ( .A(_02652_ ), .ZN(_02653_ ) );
BUF_X4 _18458_ ( .A(_02653_ ), .Z(_02654_ ) );
AND2_X1 _18459_ ( .A1(_02618_ ), .A2(_02623_ ), .ZN(_02655_ ) );
INV_X1 _18460_ ( .A(_02655_ ), .ZN(_02656_ ) );
INV_X1 _18461_ ( .A(\EXU.r2_i [15] ), .ZN(_02657_ ) );
OAI221_X1 _18462_ ( .A(_02651_ ), .B1(_02654_ ), .B2(_09429_ ), .C1(_02656_ ), .C2(_02657_ ), .ZN(_02658_ ) );
NOR2_X2 _18463_ ( .A1(_02618_ ), .A2(_02622_ ), .ZN(_02659_ ) );
BUF_X4 _18464_ ( .A(_02659_ ), .Z(_02660_ ) );
AOI21_X1 _18465_ ( .A(_02658_ ), .B1(\EXU.r2_i [31] ), .B2(_02660_ ), .ZN(_02661_ ) );
AOI21_X1 _18466_ ( .A(_02557_ ), .B1(_02640_ ), .B2(\LSU.axi_state [1] ), .ZN(_02662_ ) );
NOR2_X2 _18467_ ( .A1(_02555_ ), .A2(_02662_ ), .ZN(_02663_ ) );
NAND2_X1 _18468_ ( .A1(_02663_ ), .A2(_02550_ ), .ZN(_02664_ ) );
BUF_X4 _18469_ ( .A(_02664_ ), .Z(_02665_ ) );
INV_X1 _18470_ ( .A(\LSU.ls_axi_wdata [31] ), .ZN(_02666_ ) );
BUF_X4 _18471_ ( .A(_02663_ ), .Z(_02667_ ) );
OAI22_X1 _18472_ ( .A1(_02661_ ), .A2(_02665_ ), .B1(_02666_ ), .B2(_02667_ ), .ZN(_00905_ ) );
NAND3_X1 _18473_ ( .A1(_02649_ ), .A2(\EXU.r2_i [6] ), .A3(_02650_ ), .ZN(_02668_ ) );
OAI221_X1 _18474_ ( .A(_02668_ ), .B1(_02654_ ), .B2(_05684_ ), .C1(_02656_ ), .C2(_05663_ ), .ZN(_02669_ ) );
AOI21_X1 _18475_ ( .A(_02669_ ), .B1(\EXU.r2_i [30] ), .B2(_02660_ ), .ZN(_02670_ ) );
INV_X1 _18476_ ( .A(\LSU.ls_axi_wdata [30] ), .ZN(_02671_ ) );
OAI22_X1 _18477_ ( .A1(_02670_ ), .A2(_02665_ ), .B1(_02671_ ), .B2(_02667_ ), .ZN(_00906_ ) );
BUF_X4 _18478_ ( .A(_02656_ ), .Z(_02672_ ) );
OAI22_X1 _18479_ ( .A1(_02672_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_18_A_$_ANDNOT__Y_B ), .B1(_02654_ ), .B2(_05667_ ), .ZN(_02673_ ) );
AOI21_X1 _18480_ ( .A(_02673_ ), .B1(\EXU.r2_i [21] ), .B2(_02660_ ), .ZN(_02674_ ) );
INV_X1 _18481_ ( .A(\LSU.ls_axi_wdata [21] ), .ZN(_02675_ ) );
BUF_X4 _18482_ ( .A(_02663_ ), .Z(_02676_ ) );
OAI22_X1 _18483_ ( .A1(_02674_ ), .A2(_02665_ ), .B1(_02675_ ), .B2(_02676_ ), .ZN(_00907_ ) );
INV_X1 _18484_ ( .A(\EXU.r2_i [12] ), .ZN(_02677_ ) );
OAI22_X1 _18485_ ( .A1(_02672_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_19_A_$_ANDNOT__Y_B ), .B1(_02654_ ), .B2(_02677_ ), .ZN(_02678_ ) );
AOI21_X1 _18486_ ( .A(_02678_ ), .B1(\EXU.r2_i [20] ), .B2(_02660_ ), .ZN(_02679_ ) );
INV_X1 _18487_ ( .A(\LSU.ls_axi_wdata [20] ), .ZN(_02680_ ) );
OAI22_X1 _18488_ ( .A1(_02679_ ), .A2(_02665_ ), .B1(_02680_ ), .B2(_02676_ ), .ZN(_00908_ ) );
INV_X1 _18489_ ( .A(\EXU.r2_i [11] ), .ZN(_02681_ ) );
OAI22_X1 _18490_ ( .A1(_02672_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_20_A_$_ANDNOT__Y_B ), .B1(_02654_ ), .B2(_02681_ ), .ZN(_02682_ ) );
BUF_X4 _18491_ ( .A(_02659_ ), .Z(_02683_ ) );
AOI21_X1 _18492_ ( .A(_02682_ ), .B1(\EXU.r2_i [19] ), .B2(_02683_ ), .ZN(_02684_ ) );
INV_X1 _18493_ ( .A(\LSU.ls_axi_wdata [19] ), .ZN(_02685_ ) );
OAI22_X1 _18494_ ( .A1(_02684_ ), .A2(_02665_ ), .B1(_02685_ ), .B2(_02676_ ), .ZN(_00909_ ) );
INV_X1 _18495_ ( .A(\EXU.r2_i [10] ), .ZN(_02686_ ) );
OAI22_X1 _18496_ ( .A1(_02672_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_21_A_$_ANDNOT__Y_B ), .B1(_02654_ ), .B2(_02686_ ), .ZN(_02687_ ) );
AOI21_X1 _18497_ ( .A(_02687_ ), .B1(\EXU.r2_i [18] ), .B2(_02683_ ), .ZN(_02688_ ) );
INV_X1 _18498_ ( .A(\LSU.ls_axi_wdata [18] ), .ZN(_02689_ ) );
OAI22_X1 _18499_ ( .A1(_02688_ ), .A2(_02665_ ), .B1(_02689_ ), .B2(_02676_ ), .ZN(_00910_ ) );
OAI22_X1 _18500_ ( .A1(_02672_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_22_A_$_ANDNOT__Y_B ), .B1(_02654_ ), .B2(_05672_ ), .ZN(_02690_ ) );
AOI21_X1 _18501_ ( .A(_02690_ ), .B1(\EXU.r2_i [17] ), .B2(_02683_ ), .ZN(_02691_ ) );
INV_X1 _18502_ ( .A(\LSU.ls_axi_wdata [17] ), .ZN(_02692_ ) );
OAI22_X1 _18503_ ( .A1(_02691_ ), .A2(_02665_ ), .B1(_02692_ ), .B2(_02676_ ), .ZN(_00911_ ) );
INV_X1 _18504_ ( .A(\EXU.r2_i [8] ), .ZN(_02693_ ) );
OAI22_X1 _18505_ ( .A1(_02672_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_23_A_$_ANDNOT__Y_B ), .B1(_02654_ ), .B2(_02693_ ), .ZN(_02694_ ) );
AOI21_X1 _18506_ ( .A(_02694_ ), .B1(\EXU.r2_i [16] ), .B2(_02683_ ), .ZN(_02695_ ) );
INV_X1 _18507_ ( .A(\LSU.ls_axi_wdata [16] ), .ZN(_02696_ ) );
OAI22_X1 _18508_ ( .A1(_02695_ ), .A2(_02665_ ), .B1(_02696_ ), .B2(_02676_ ), .ZN(_00912_ ) );
NOR4_X1 _18509_ ( .A1(_05353_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_16_A_$_ANDNOT__Y_B ), .A3(_02545_ ), .A4(_05361_ ), .ZN(_02697_ ) );
BUF_X4 _18510_ ( .A(_02659_ ), .Z(_02698_ ) );
AOI21_X1 _18511_ ( .A(_02697_ ), .B1(_02698_ ), .B2(\EXU.r2_i [15] ), .ZN(_02699_ ) );
INV_X1 _18512_ ( .A(\LSU.ls_axi_wdata [15] ), .ZN(_02700_ ) );
OAI22_X1 _18513_ ( .A1(_02699_ ), .A2(_02665_ ), .B1(_02700_ ), .B2(_02676_ ), .ZN(_00913_ ) );
NOR4_X1 _18514_ ( .A1(_05353_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_17_A_$_ANDNOT__Y_B ), .A3(_02545_ ), .A4(_05361_ ), .ZN(_02701_ ) );
AOI21_X1 _18515_ ( .A(_02701_ ), .B1(_02698_ ), .B2(\EXU.r2_i [14] ), .ZN(_02702_ ) );
INV_X1 _18516_ ( .A(\LSU.ls_axi_wdata [14] ), .ZN(_02703_ ) );
OAI22_X1 _18517_ ( .A1(_02702_ ), .A2(_02665_ ), .B1(_02703_ ), .B2(_02676_ ), .ZN(_00914_ ) );
NOR4_X1 _18518_ ( .A1(_05353_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_18_A_$_ANDNOT__Y_B ), .A3(_02545_ ), .A4(_05361_ ), .ZN(_02704_ ) );
AOI21_X1 _18519_ ( .A(_02704_ ), .B1(_02698_ ), .B2(\EXU.r2_i [13] ), .ZN(_02705_ ) );
BUF_X4 _18520_ ( .A(_02664_ ), .Z(_02706_ ) );
INV_X1 _18521_ ( .A(\LSU.ls_axi_wdata [13] ), .ZN(_02707_ ) );
OAI22_X1 _18522_ ( .A1(_02705_ ), .A2(_02706_ ), .B1(_02707_ ), .B2(_02676_ ), .ZN(_00915_ ) );
NOR4_X1 _18523_ ( .A1(_05353_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_19_A_$_ANDNOT__Y_B ), .A3(_02545_ ), .A4(_05361_ ), .ZN(_02708_ ) );
AOI21_X1 _18524_ ( .A(_02708_ ), .B1(_02698_ ), .B2(\EXU.r2_i [12] ), .ZN(_02709_ ) );
INV_X1 _18525_ ( .A(\LSU.ls_axi_wdata [12] ), .ZN(_02710_ ) );
OAI22_X1 _18526_ ( .A1(_02709_ ), .A2(_02706_ ), .B1(_02710_ ), .B2(_02676_ ), .ZN(_00916_ ) );
NAND3_X1 _18527_ ( .A1(_02649_ ), .A2(\EXU.r2_i [5] ), .A3(_02650_ ), .ZN(_02711_ ) );
OAI221_X1 _18528_ ( .A(_02711_ ), .B1(_02653_ ), .B2(_05688_ ), .C1(_02656_ ), .C2(_05667_ ), .ZN(_02712_ ) );
AOI21_X1 _18529_ ( .A(_02712_ ), .B1(\EXU.r2_i [29] ), .B2(_02683_ ), .ZN(_02713_ ) );
INV_X1 _18530_ ( .A(\LSU.ls_axi_wdata [29] ), .ZN(_02714_ ) );
BUF_X4 _18531_ ( .A(_02663_ ), .Z(_02715_ ) );
OAI22_X1 _18532_ ( .A1(_02713_ ), .A2(_02706_ ), .B1(_02714_ ), .B2(_02715_ ), .ZN(_00917_ ) );
NOR4_X1 _18533_ ( .A1(_05353_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_20_A_$_ANDNOT__Y_B ), .A3(_02545_ ), .A4(_05361_ ), .ZN(_02716_ ) );
AOI21_X1 _18534_ ( .A(_02716_ ), .B1(_02698_ ), .B2(\EXU.r2_i [11] ), .ZN(_02717_ ) );
INV_X1 _18535_ ( .A(\LSU.ls_axi_wdata [11] ), .ZN(_02718_ ) );
OAI22_X1 _18536_ ( .A1(_02717_ ), .A2(_02706_ ), .B1(_02718_ ), .B2(_02715_ ), .ZN(_00918_ ) );
NOR4_X1 _18537_ ( .A1(_05353_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_21_A_$_ANDNOT__Y_B ), .A3(_02545_ ), .A4(_05361_ ), .ZN(_02719_ ) );
AOI21_X1 _18538_ ( .A(_02719_ ), .B1(_02698_ ), .B2(\EXU.r2_i [10] ), .ZN(_02720_ ) );
INV_X1 _18539_ ( .A(\LSU.ls_axi_wdata [10] ), .ZN(_02721_ ) );
OAI22_X1 _18540_ ( .A1(_02720_ ), .A2(_02706_ ), .B1(_02721_ ), .B2(_02715_ ), .ZN(_00919_ ) );
NOR4_X1 _18541_ ( .A1(_05353_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_22_A_$_ANDNOT__Y_B ), .A3(_02545_ ), .A4(_05361_ ), .ZN(_02722_ ) );
AOI21_X1 _18542_ ( .A(_02722_ ), .B1(_02698_ ), .B2(\EXU.r2_i [9] ), .ZN(_02723_ ) );
INV_X1 _18543_ ( .A(\LSU.ls_axi_wdata [9] ), .ZN(_02724_ ) );
OAI22_X1 _18544_ ( .A1(_02723_ ), .A2(_02706_ ), .B1(_02724_ ), .B2(_02715_ ), .ZN(_00920_ ) );
NOR4_X1 _18545_ ( .A1(_05353_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_23_A_$_ANDNOT__Y_B ), .A3(_02545_ ), .A4(_05361_ ), .ZN(_02725_ ) );
AOI21_X1 _18546_ ( .A(_02725_ ), .B1(_02698_ ), .B2(\EXU.r2_i [8] ), .ZN(_02726_ ) );
INV_X1 _18547_ ( .A(\LSU.ls_axi_wdata [8] ), .ZN(_02727_ ) );
OAI22_X1 _18548_ ( .A1(_02726_ ), .A2(_02706_ ), .B1(_02727_ ), .B2(_02715_ ), .ZN(_00921_ ) );
BUF_X4 _18549_ ( .A(_02663_ ), .Z(_02728_ ) );
NAND4_X1 _18550_ ( .A1(_02698_ ), .A2(\EXU.r2_i [7] ), .A3(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ), .A4(_02728_ ), .ZN(_02729_ ) );
INV_X1 _18551_ ( .A(\LSU.ls_axi_wdata [7] ), .ZN(_02730_ ) );
OAI21_X1 _18552_ ( .A(_02729_ ), .B1(_02730_ ), .B2(_02667_ ), .ZN(_00922_ ) );
NAND4_X1 _18553_ ( .A1(_02698_ ), .A2(\EXU.r2_i [6] ), .A3(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ), .A4(_02728_ ), .ZN(_02731_ ) );
INV_X1 _18554_ ( .A(\LSU.ls_axi_wdata [6] ), .ZN(_02732_ ) );
OAI21_X1 _18555_ ( .A(_02731_ ), .B1(_02732_ ), .B2(_02667_ ), .ZN(_00923_ ) );
NAND4_X1 _18556_ ( .A1(_02660_ ), .A2(\EXU.r2_i [5] ), .A3(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ), .A4(_02728_ ), .ZN(_02733_ ) );
INV_X1 _18557_ ( .A(\LSU.ls_axi_wdata [5] ), .ZN(_02734_ ) );
OAI21_X1 _18558_ ( .A(_02733_ ), .B1(_02734_ ), .B2(_02667_ ), .ZN(_00924_ ) );
NAND4_X1 _18559_ ( .A1(_02660_ ), .A2(\EXU.r2_i [4] ), .A3(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ), .A4(_02728_ ), .ZN(_02735_ ) );
INV_X1 _18560_ ( .A(\LSU.ls_axi_wdata [4] ), .ZN(_02736_ ) );
OAI21_X1 _18561_ ( .A(_02735_ ), .B1(_02736_ ), .B2(_02667_ ), .ZN(_00925_ ) );
NAND4_X1 _18562_ ( .A1(_02660_ ), .A2(\EXU.r2_i [3] ), .A3(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ), .A4(_02728_ ), .ZN(_02737_ ) );
INV_X1 _18563_ ( .A(\LSU.ls_axi_wdata [3] ), .ZN(_02738_ ) );
OAI21_X1 _18564_ ( .A(_02737_ ), .B1(_02738_ ), .B2(_02667_ ), .ZN(_00926_ ) );
NAND4_X1 _18565_ ( .A1(_02660_ ), .A2(\EXU.r2_i [2] ), .A3(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ), .A4(_02728_ ), .ZN(_02739_ ) );
INV_X1 _18566_ ( .A(\LSU.ls_axi_wdata [2] ), .ZN(_02740_ ) );
OAI21_X1 _18567_ ( .A(_02739_ ), .B1(_02740_ ), .B2(_02667_ ), .ZN(_00927_ ) );
NAND3_X1 _18568_ ( .A1(_02649_ ), .A2(\EXU.r2_i [4] ), .A3(_02650_ ), .ZN(_02741_ ) );
NAND3_X1 _18569_ ( .A1(_02619_ ), .A2(\EXU.r2_i [20] ), .A3(_02650_ ), .ZN(_02742_ ) );
OAI211_X1 _18570_ ( .A(_02741_ ), .B(_02742_ ), .C1(_02672_ ), .C2(_02677_ ), .ZN(_02743_ ) );
AOI21_X1 _18571_ ( .A(_02743_ ), .B1(\EXU.r2_i [28] ), .B2(_02683_ ), .ZN(_02744_ ) );
INV_X1 _18572_ ( .A(\LSU.ls_axi_wdata [28] ), .ZN(_02745_ ) );
OAI22_X1 _18573_ ( .A1(_02744_ ), .A2(_02706_ ), .B1(_02745_ ), .B2(_02715_ ), .ZN(_00928_ ) );
NAND4_X1 _18574_ ( .A1(_02660_ ), .A2(\EXU.r2_i [1] ), .A3(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ), .A4(_02728_ ), .ZN(_02746_ ) );
INV_X1 _18575_ ( .A(\LSU.ls_axi_wdata [1] ), .ZN(_02747_ ) );
OAI21_X1 _18576_ ( .A(_02746_ ), .B1(_02747_ ), .B2(_02667_ ), .ZN(_00929_ ) );
NAND4_X1 _18577_ ( .A1(_02660_ ), .A2(\EXU.r2_i [0] ), .A3(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ), .A4(_02728_ ), .ZN(_02748_ ) );
INV_X1 _18578_ ( .A(\LSU.ls_axi_wdata [0] ), .ZN(_02749_ ) );
OAI21_X1 _18579_ ( .A(_02748_ ), .B1(_02749_ ), .B2(_02667_ ), .ZN(_00930_ ) );
NAND3_X1 _18580_ ( .A1(_02649_ ), .A2(\EXU.r2_i [3] ), .A3(_02622_ ), .ZN(_02750_ ) );
OAI221_X1 _18581_ ( .A(_02750_ ), .B1(_02653_ ), .B2(_05700_ ), .C1(_02656_ ), .C2(_02681_ ), .ZN(_02751_ ) );
AOI21_X1 _18582_ ( .A(_02751_ ), .B1(\EXU.r2_i [27] ), .B2(_02683_ ), .ZN(_02752_ ) );
INV_X1 _18583_ ( .A(\LSU.ls_axi_wdata [27] ), .ZN(_02753_ ) );
OAI22_X1 _18584_ ( .A1(_02752_ ), .A2(_02706_ ), .B1(_02753_ ), .B2(_02715_ ), .ZN(_00931_ ) );
NAND3_X1 _18585_ ( .A1(_02649_ ), .A2(\EXU.r2_i [2] ), .A3(_02650_ ), .ZN(_02754_ ) );
NAND3_X1 _18586_ ( .A1(_02619_ ), .A2(\EXU.r2_i [18] ), .A3(_02650_ ), .ZN(_02755_ ) );
OAI211_X1 _18587_ ( .A(_02754_ ), .B(_02755_ ), .C1(_02672_ ), .C2(_02686_ ), .ZN(_02756_ ) );
AOI21_X1 _18588_ ( .A(_02756_ ), .B1(\EXU.r2_i [26] ), .B2(_02683_ ), .ZN(_02757_ ) );
INV_X1 _18589_ ( .A(\LSU.ls_axi_wdata [26] ), .ZN(_02758_ ) );
OAI22_X1 _18590_ ( .A1(_02757_ ), .A2(_02706_ ), .B1(_02758_ ), .B2(_02715_ ), .ZN(_00932_ ) );
NAND3_X1 _18591_ ( .A1(_02649_ ), .A2(\EXU.r2_i [1] ), .A3(_02622_ ), .ZN(_02759_ ) );
OAI221_X1 _18592_ ( .A(_02759_ ), .B1(_02653_ ), .B2(_05694_ ), .C1(_02656_ ), .C2(_05672_ ), .ZN(_02760_ ) );
AOI21_X1 _18593_ ( .A(_02760_ ), .B1(\EXU.r2_i [25] ), .B2(_02683_ ), .ZN(_02761_ ) );
INV_X1 _18594_ ( .A(\LSU.ls_axi_wdata [25] ), .ZN(_02762_ ) );
OAI22_X1 _18595_ ( .A1(_02761_ ), .A2(_02664_ ), .B1(_02762_ ), .B2(_02715_ ), .ZN(_00933_ ) );
NAND3_X1 _18596_ ( .A1(_02649_ ), .A2(\EXU.r2_i [0] ), .A3(_02650_ ), .ZN(_02763_ ) );
NAND3_X1 _18597_ ( .A1(_02619_ ), .A2(\EXU.r2_i [16] ), .A3(_02650_ ), .ZN(_02764_ ) );
OAI211_X1 _18598_ ( .A(_02763_ ), .B(_02764_ ), .C1(_02656_ ), .C2(_02693_ ), .ZN(_02765_ ) );
AOI21_X1 _18599_ ( .A(_02765_ ), .B1(\EXU.r2_i [24] ), .B2(_02683_ ), .ZN(_02766_ ) );
INV_X1 _18600_ ( .A(\LSU.ls_axi_wdata [24] ), .ZN(_02767_ ) );
OAI22_X1 _18601_ ( .A1(_02766_ ), .A2(_02664_ ), .B1(_02767_ ), .B2(_02715_ ), .ZN(_00934_ ) );
OAI22_X1 _18602_ ( .A1(_02672_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_16_A_$_ANDNOT__Y_B ), .B1(_02654_ ), .B2(_02657_ ), .ZN(_02768_ ) );
AOI21_X1 _18603_ ( .A(_02768_ ), .B1(\EXU.r2_i [23] ), .B2(_02659_ ), .ZN(_02769_ ) );
INV_X1 _18604_ ( .A(\LSU.ls_axi_wdata [23] ), .ZN(_02770_ ) );
OAI22_X1 _18605_ ( .A1(_02769_ ), .A2(_02664_ ), .B1(_02770_ ), .B2(_02728_ ), .ZN(_00935_ ) );
OAI22_X1 _18606_ ( .A1(_02672_ ), .A2(\LSU.ls_wdata_i_$_MUX__Y_17_A_$_ANDNOT__Y_B ), .B1(_02654_ ), .B2(_05663_ ), .ZN(_02771_ ) );
AOI21_X1 _18607_ ( .A(_02771_ ), .B1(\EXU.r2_i [22] ), .B2(_02659_ ), .ZN(_02772_ ) );
INV_X1 _18608_ ( .A(\LSU.ls_axi_wdata [22] ), .ZN(_02773_ ) );
OAI22_X1 _18609_ ( .A1(_02772_ ), .A2(_02664_ ), .B1(_02773_ ), .B2(_02728_ ), .ZN(_00936_ ) );
MUX2_X1 _18610_ ( .A(\LSU.ls_axi_wlast ), .B(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ), .S(_02559_ ), .Z(_00937_ ) );
MUX2_X1 _18611_ ( .A(\LSU.ls_axi_wvalid ), .B(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ), .S(_02663_ ), .Z(_00938_ ) );
BUF_X2 _18612_ ( .A(_02646_ ), .Z(\LSU.ls_axi_rready_$_ANDNOT__A_Y ) );
AND2_X2 _18613_ ( .A1(_02655_ ), .A2(_06006_ ), .ZN(_02774_ ) );
NOR2_X1 _18614_ ( .A1(_07688_ ), .A2(_04058_ ), .ZN(_02775_ ) );
AND3_X1 _18615_ ( .A1(_02774_ ), .A2(_04716_ ), .A3(_02775_ ), .ZN(_02776_ ) );
AND3_X1 _18616_ ( .A1(_02618_ ), .A2(_06006_ ), .A3(_02622_ ), .ZN(_02777_ ) );
AND2_X1 _18617_ ( .A1(_02777_ ), .A2(_04711_ ), .ZN(_02778_ ) );
AND2_X1 _18618_ ( .A1(_02778_ ), .A2(_02775_ ), .ZN(_02779_ ) );
AND2_X1 _18619_ ( .A1(_02659_ ), .A2(_06006_ ), .ZN(_02780_ ) );
BUF_X4 _18620_ ( .A(_02780_ ), .Z(_02781_ ) );
NOR2_X1 _18621_ ( .A1(_07726_ ), .A2(_04058_ ), .ZN(_02782_ ) );
AND3_X1 _18622_ ( .A1(_02781_ ), .A2(_04716_ ), .A3(_02782_ ), .ZN(_02783_ ) );
NOR3_X1 _18623_ ( .A1(_02776_ ), .A2(_02779_ ), .A3(_02783_ ), .ZN(_02784_ ) );
BUF_X4 _18624_ ( .A(_02784_ ), .Z(_02785_ ) );
AND2_X2 _18625_ ( .A1(_02781_ ), .A2(_04711_ ), .ZN(_02786_ ) );
NOR2_X1 _18626_ ( .A1(_07756_ ), .A2(_04105_ ), .ZN(_02787_ ) );
NAND2_X2 _18627_ ( .A1(_02786_ ), .A2(_02787_ ), .ZN(_02788_ ) );
BUF_X4 _18628_ ( .A(_02788_ ), .Z(_02789_ ) );
AND2_X1 _18629_ ( .A1(_02774_ ), .A2(_04711_ ), .ZN(_02790_ ) );
BUF_X4 _18630_ ( .A(_02790_ ), .Z(_02791_ ) );
NOR2_X1 _18631_ ( .A1(_07790_ ), .A2(_04105_ ), .ZN(_02792_ ) );
NOR3_X1 _18632_ ( .A1(_02618_ ), .A2(_04414_ ), .A3(_02623_ ), .ZN(_02793_ ) );
CLKBUF_X2 _18633_ ( .A(_02793_ ), .Z(_02794_ ) );
AND2_X1 _18634_ ( .A1(_02794_ ), .A2(_04711_ ), .ZN(_02795_ ) );
AOI22_X2 _18635_ ( .A1(_02791_ ), .A2(_02792_ ), .B1(_02782_ ), .B2(_02795_ ), .ZN(_02796_ ) );
BUF_X4 _18636_ ( .A(_02796_ ), .Z(_02797_ ) );
BUF_X4 _18637_ ( .A(_02781_ ), .Z(_02798_ ) );
BUF_X4 _18638_ ( .A(_05525_ ), .Z(_02799_ ) );
BUF_X4 _18639_ ( .A(_02799_ ), .Z(_02800_ ) );
NAND3_X1 _18640_ ( .A1(_02798_ ), .A2(_02800_ ), .A3(_02775_ ), .ZN(_02801_ ) );
NAND4_X1 _18641_ ( .A1(_02785_ ), .A2(_02789_ ), .A3(_02797_ ), .A4(_02801_ ), .ZN(_02802_ ) );
MUX2_X1 _18642_ ( .A(\EXU.ls_rdata_i [31] ), .B(_02802_ ), .S(_02647_ ), .Z(_00939_ ) );
NOR2_X1 _18643_ ( .A1(_07701_ ), .A2(_04105_ ), .ZN(_02803_ ) );
NAND3_X1 _18644_ ( .A1(_02798_ ), .A2(_02800_ ), .A3(_02803_ ), .ZN(_02804_ ) );
NAND4_X1 _18645_ ( .A1(_02785_ ), .A2(_02789_ ), .A3(_02797_ ), .A4(_02804_ ), .ZN(_02805_ ) );
MUX2_X1 _18646_ ( .A(\EXU.ls_rdata_i [30] ), .B(_02805_ ), .S(_02647_ ), .Z(_00940_ ) );
BUF_X2 _18647_ ( .A(_04058_ ), .Z(_02806_ ) );
BUF_X4 _18648_ ( .A(_02806_ ), .Z(_02807_ ) );
NOR2_X1 _18649_ ( .A1(_07707_ ), .A2(_02807_ ), .ZN(_02808_ ) );
NAND3_X1 _18650_ ( .A1(_02798_ ), .A2(_02800_ ), .A3(_02808_ ), .ZN(_02809_ ) );
NAND4_X1 _18651_ ( .A1(_02785_ ), .A2(_02789_ ), .A3(_02797_ ), .A4(_02809_ ), .ZN(_02810_ ) );
MUX2_X1 _18652_ ( .A(\EXU.ls_rdata_i [21] ), .B(_02810_ ), .S(_02647_ ), .Z(_00941_ ) );
NOR2_X1 _18653_ ( .A1(_07710_ ), .A2(_07831_ ), .ZN(_02811_ ) );
NAND3_X1 _18654_ ( .A1(_02798_ ), .A2(_02800_ ), .A3(_02811_ ), .ZN(_02812_ ) );
NAND4_X1 _18655_ ( .A1(_02785_ ), .A2(_02789_ ), .A3(_02797_ ), .A4(_02812_ ), .ZN(_02813_ ) );
MUX2_X1 _18656_ ( .A(\EXU.ls_rdata_i [20] ), .B(_02813_ ), .S(_02647_ ), .Z(_00942_ ) );
NOR2_X1 _18657_ ( .A1(_07713_ ), .A2(_07831_ ), .ZN(_02814_ ) );
NAND3_X1 _18658_ ( .A1(_02798_ ), .A2(_02800_ ), .A3(_02814_ ), .ZN(_02815_ ) );
NAND4_X1 _18659_ ( .A1(_02785_ ), .A2(_02789_ ), .A3(_02797_ ), .A4(_02815_ ), .ZN(_02816_ ) );
MUX2_X1 _18660_ ( .A(\EXU.ls_rdata_i [19] ), .B(_02816_ ), .S(_02647_ ), .Z(_00943_ ) );
NOR2_X1 _18661_ ( .A1(_07716_ ), .A2(_02807_ ), .ZN(_02817_ ) );
NAND3_X1 _18662_ ( .A1(_02798_ ), .A2(_02800_ ), .A3(_02817_ ), .ZN(_02818_ ) );
NAND4_X1 _18663_ ( .A1(_02785_ ), .A2(_02789_ ), .A3(_02797_ ), .A4(_02818_ ), .ZN(_02819_ ) );
MUX2_X1 _18664_ ( .A(\EXU.ls_rdata_i [18] ), .B(_02819_ ), .S(_02647_ ), .Z(_00944_ ) );
NOR2_X1 _18665_ ( .A1(_07719_ ), .A2(_02807_ ), .ZN(_02820_ ) );
NAND3_X1 _18666_ ( .A1(_02798_ ), .A2(_02799_ ), .A3(_02820_ ), .ZN(_02821_ ) );
NAND4_X1 _18667_ ( .A1(_02785_ ), .A2(_02789_ ), .A3(_02797_ ), .A4(_02821_ ), .ZN(_02822_ ) );
BUF_X4 _18668_ ( .A(_02646_ ), .Z(_02823_ ) );
MUX2_X1 _18669_ ( .A(\EXU.ls_rdata_i [17] ), .B(_02822_ ), .S(_02823_ ), .Z(_00945_ ) );
NOR2_X1 _18670_ ( .A1(_07723_ ), .A2(_02807_ ), .ZN(_02824_ ) );
NAND3_X1 _18671_ ( .A1(_02798_ ), .A2(_02799_ ), .A3(_02824_ ), .ZN(_02825_ ) );
NAND4_X1 _18672_ ( .A1(_02785_ ), .A2(_02789_ ), .A3(_02797_ ), .A4(_02825_ ), .ZN(_02826_ ) );
MUX2_X1 _18673_ ( .A(\EXU.ls_rdata_i [16] ), .B(_02826_ ), .S(_02823_ ), .Z(_00946_ ) );
NAND3_X1 _18674_ ( .A1(_02781_ ), .A2(_02799_ ), .A3(_02782_ ), .ZN(_02827_ ) );
AND3_X1 _18675_ ( .A1(_02796_ ), .A2(_02788_ ), .A3(_02827_ ), .ZN(_02828_ ) );
NOR2_X1 _18676_ ( .A1(_02779_ ), .A2(_02783_ ), .ZN(_02829_ ) );
AND2_X1 _18677_ ( .A1(_02781_ ), .A2(_04716_ ), .ZN(_02830_ ) );
BUF_X2 _18678_ ( .A(_02830_ ), .Z(_02831_ ) );
INV_X1 _18679_ ( .A(_02831_ ), .ZN(_02832_ ) );
AND4_X1 _18680_ ( .A1(_06007_ ), .A2(_02655_ ), .A3(_05543_ ), .A4(_02775_ ), .ZN(_02833_ ) );
AND4_X1 _18681_ ( .A1(_06007_ ), .A2(_02659_ ), .A3(_05543_ ), .A4(_02782_ ), .ZN(_02834_ ) );
NOR2_X1 _18682_ ( .A1(_02833_ ), .A2(_02834_ ), .ZN(_02835_ ) );
AND2_X1 _18683_ ( .A1(_02774_ ), .A2(_04716_ ), .ZN(_02836_ ) );
NOR2_X1 _18684_ ( .A1(_02835_ ), .A2(_02836_ ), .ZN(_02837_ ) );
OAI21_X1 _18685_ ( .A(_02832_ ), .B1(_02837_ ), .B2(_02776_ ), .ZN(_02838_ ) );
NAND3_X1 _18686_ ( .A1(_02828_ ), .A2(_02829_ ), .A3(_02838_ ), .ZN(_02839_ ) );
MUX2_X1 _18687_ ( .A(\EXU.ls_rdata_i [15] ), .B(_02839_ ), .S(_02823_ ), .Z(_00947_ ) );
AND2_X1 _18688_ ( .A1(_02774_ ), .A2(_05543_ ), .ZN(_02840_ ) );
NOR2_X1 _18689_ ( .A1(_02836_ ), .A2(_02840_ ), .ZN(_02841_ ) );
INV_X1 _18690_ ( .A(_02841_ ), .ZN(_02842_ ) );
NAND3_X1 _18691_ ( .A1(_02842_ ), .A2(_02832_ ), .A3(_02803_ ), .ZN(_02843_ ) );
AND2_X2 _18692_ ( .A1(_02796_ ), .A2(_02788_ ), .ZN(_02844_ ) );
INV_X1 _18693_ ( .A(_02779_ ), .ZN(_02845_ ) );
NAND2_X1 _18694_ ( .A1(_02780_ ), .A2(_05543_ ), .ZN(_02846_ ) );
BUF_X2 _18695_ ( .A(_06007_ ), .Z(_02847_ ) );
OAI211_X1 _18696_ ( .A(_02659_ ), .B(_02847_ ), .C1(_05528_ ), .C2(_02799_ ), .ZN(_02848_ ) );
NAND2_X1 _18697_ ( .A1(_02846_ ), .A2(_02848_ ), .ZN(_02849_ ) );
NOR2_X1 _18698_ ( .A1(_07730_ ), .A2(_04058_ ), .ZN(_02850_ ) );
NAND2_X1 _18699_ ( .A1(_02849_ ), .A2(_02850_ ), .ZN(_02851_ ) );
NAND4_X1 _18700_ ( .A1(_02843_ ), .A2(_02844_ ), .A3(_02845_ ), .A4(_02851_ ), .ZN(_02852_ ) );
NAND2_X1 _18701_ ( .A1(_02852_ ), .A2(\LSU.ls_axi_rready_$_ANDNOT__A_Y ), .ZN(_02853_ ) );
OAI21_X1 _18702_ ( .A(_02853_ ), .B1(_06556_ ), .B2(\LSU.ls_axi_rready_$_ANDNOT__A_Y ), .ZN(_00948_ ) );
OR2_X1 _18703_ ( .A1(_07740_ ), .A2(_02806_ ), .ZN(_02854_ ) );
OR3_X1 _18704_ ( .A1(_02841_ ), .A2(_02831_ ), .A3(_02854_ ), .ZN(_02855_ ) );
NOR2_X1 _18705_ ( .A1(_07733_ ), .A2(_02806_ ), .ZN(_02856_ ) );
NAND2_X1 _18706_ ( .A1(_02849_ ), .A2(_02856_ ), .ZN(_02857_ ) );
NAND4_X1 _18707_ ( .A1(_02855_ ), .A2(_02844_ ), .A3(_02845_ ), .A4(_02857_ ), .ZN(_02858_ ) );
MUX2_X1 _18708_ ( .A(\EXU.ls_rdata_i [13] ), .B(_02858_ ), .S(_02823_ ), .Z(_00949_ ) );
NOR2_X1 _18709_ ( .A1(_07775_ ), .A2(_02807_ ), .ZN(_02859_ ) );
NAND3_X1 _18710_ ( .A1(_02842_ ), .A2(_02832_ ), .A3(_02859_ ), .ZN(_02860_ ) );
NOR2_X1 _18711_ ( .A1(_07737_ ), .A2(_02806_ ), .ZN(_02861_ ) );
NAND2_X1 _18712_ ( .A1(_02849_ ), .A2(_02861_ ), .ZN(_02862_ ) );
NAND4_X1 _18713_ ( .A1(_02860_ ), .A2(_02844_ ), .A3(_02845_ ), .A4(_02862_ ), .ZN(_02863_ ) );
MUX2_X1 _18714_ ( .A(\EXU.ls_rdata_i [12] ), .B(_02863_ ), .S(_02823_ ), .Z(_00950_ ) );
AND2_X2 _18715_ ( .A1(_02781_ ), .A2(_02799_ ), .ZN(_02864_ ) );
INV_X1 _18716_ ( .A(_02864_ ), .ZN(_02865_ ) );
OR2_X1 _18717_ ( .A1(_02865_ ), .A2(_02854_ ), .ZN(_02866_ ) );
NAND4_X1 _18718_ ( .A1(_02785_ ), .A2(_02866_ ), .A3(_02788_ ), .A4(_02796_ ), .ZN(_02867_ ) );
MUX2_X1 _18719_ ( .A(\EXU.ls_rdata_i [29] ), .B(_02867_ ), .S(_02823_ ), .Z(_00951_ ) );
NOR2_X1 _18720_ ( .A1(_07778_ ), .A2(_04105_ ), .ZN(_02868_ ) );
NAND3_X1 _18721_ ( .A1(_02842_ ), .A2(_02832_ ), .A3(_02868_ ), .ZN(_02869_ ) );
NAND3_X1 _18722_ ( .A1(_02869_ ), .A2(_02844_ ), .A3(_02845_ ), .ZN(_02870_ ) );
NOR2_X1 _18723_ ( .A1(_07743_ ), .A2(_04105_ ), .ZN(_02871_ ) );
AND2_X1 _18724_ ( .A1(_02849_ ), .A2(_02871_ ), .ZN(_02872_ ) );
OAI21_X1 _18725_ ( .A(_02647_ ), .B1(_02870_ ), .B2(_02872_ ), .ZN(_02873_ ) );
OAI21_X1 _18726_ ( .A(_02873_ ), .B1(_06764_ ), .B2(\LSU.ls_axi_rready_$_ANDNOT__A_Y ), .ZN(_00952_ ) );
OR2_X1 _18727_ ( .A1(_07781_ ), .A2(_02806_ ), .ZN(_02874_ ) );
OR3_X1 _18728_ ( .A1(_02841_ ), .A2(_02831_ ), .A3(_02874_ ), .ZN(_02875_ ) );
NOR2_X1 _18729_ ( .A1(_07746_ ), .A2(_02806_ ), .ZN(_02876_ ) );
NAND2_X1 _18730_ ( .A1(_02849_ ), .A2(_02876_ ), .ZN(_02877_ ) );
NAND4_X1 _18731_ ( .A1(_02875_ ), .A2(_02844_ ), .A3(_02845_ ), .A4(_02877_ ), .ZN(_02878_ ) );
NAND2_X1 _18732_ ( .A1(_02878_ ), .A2(\LSU.ls_axi_rready_$_ANDNOT__A_Y ), .ZN(_02879_ ) );
OAI21_X1 _18733_ ( .A(_02879_ ), .B1(_06810_ ), .B2(\LSU.ls_axi_rready_$_ANDNOT__A_Y ), .ZN(_00953_ ) );
OR2_X1 _18734_ ( .A1(_07784_ ), .A2(_02806_ ), .ZN(_02880_ ) );
OR3_X1 _18735_ ( .A1(_02841_ ), .A2(_02831_ ), .A3(_02880_ ), .ZN(_02881_ ) );
NOR2_X1 _18736_ ( .A1(_07749_ ), .A2(_04105_ ), .ZN(_02882_ ) );
NAND2_X1 _18737_ ( .A1(_02849_ ), .A2(_02882_ ), .ZN(_02883_ ) );
NAND4_X1 _18738_ ( .A1(_02881_ ), .A2(_02844_ ), .A3(_02845_ ), .A4(_02883_ ), .ZN(_02884_ ) );
MUX2_X1 _18739_ ( .A(\EXU.ls_rdata_i [9] ), .B(_02884_ ), .S(_02823_ ), .Z(_00954_ ) );
OR2_X1 _18740_ ( .A1(_07787_ ), .A2(_02806_ ), .ZN(_02885_ ) );
OR3_X1 _18741_ ( .A1(_02841_ ), .A2(_02831_ ), .A3(_02885_ ), .ZN(_02886_ ) );
NOR2_X1 _18742_ ( .A1(_07752_ ), .A2(_02806_ ), .ZN(_02887_ ) );
NAND2_X1 _18743_ ( .A1(_02849_ ), .A2(_02887_ ), .ZN(_02888_ ) );
NAND4_X1 _18744_ ( .A1(_02886_ ), .A2(_02844_ ), .A3(_02845_ ), .A4(_02888_ ), .ZN(_02889_ ) );
NAND2_X1 _18745_ ( .A1(_02889_ ), .A2(\LSU.ls_axi_rready_$_ANDNOT__A_Y ), .ZN(_02890_ ) );
OAI21_X1 _18746_ ( .A(_02890_ ), .B1(_06917_ ), .B2(\LSU.ls_axi_rready_$_ANDNOT__A_Y ), .ZN(_00955_ ) );
BUF_X4 _18747_ ( .A(_02786_ ), .Z(_02891_ ) );
OAI21_X1 _18748_ ( .A(_02787_ ), .B1(_02891_ ), .B2(_02864_ ), .ZN(_02892_ ) );
AND2_X1 _18749_ ( .A1(_02795_ ), .A2(_02782_ ), .ZN(_02893_ ) );
AND2_X1 _18750_ ( .A1(_02791_ ), .A2(_02792_ ), .ZN(_02894_ ) );
INV_X1 _18751_ ( .A(_02894_ ), .ZN(_02895_ ) );
NAND2_X1 _18752_ ( .A1(_02774_ ), .A2(_05570_ ), .ZN(_02896_ ) );
NAND2_X1 _18753_ ( .A1(_02841_ ), .A2(_02896_ ), .ZN(_02897_ ) );
NAND2_X1 _18754_ ( .A1(_02897_ ), .A2(_02792_ ), .ZN(_02898_ ) );
NAND2_X1 _18755_ ( .A1(_02780_ ), .A2(_05570_ ), .ZN(_02899_ ) );
NAND2_X1 _18756_ ( .A1(_02846_ ), .A2(_02899_ ), .ZN(_02900_ ) );
OAI21_X1 _18757_ ( .A(_02787_ ), .B1(_02900_ ), .B2(_02831_ ), .ZN(_02901_ ) );
BUF_X2 _18758_ ( .A(_05570_ ), .Z(_02902_ ) );
NAND3_X1 _18759_ ( .A1(_02777_ ), .A2(_02902_ ), .A3(_02775_ ), .ZN(_02903_ ) );
NAND3_X1 _18760_ ( .A1(_02794_ ), .A2(_02902_ ), .A3(_02782_ ), .ZN(_02904_ ) );
AND2_X1 _18761_ ( .A1(_02903_ ), .A2(_02904_ ), .ZN(_02905_ ) );
NAND3_X1 _18762_ ( .A1(_02898_ ), .A2(_02901_ ), .A3(_02905_ ), .ZN(_02906_ ) );
INV_X1 _18763_ ( .A(_02778_ ), .ZN(_02907_ ) );
BUF_X4 _18764_ ( .A(_02907_ ), .Z(_02908_ ) );
AOI21_X1 _18765_ ( .A(_02779_ ), .B1(_02906_ ), .B2(_02908_ ), .ZN(_02909_ ) );
OAI21_X1 _18766_ ( .A(_02895_ ), .B1(_02909_ ), .B2(_02791_ ), .ZN(_02910_ ) );
INV_X1 _18767_ ( .A(_02795_ ), .ZN(_02911_ ) );
AOI21_X1 _18768_ ( .A(_02893_ ), .B1(_02910_ ), .B2(_02911_ ), .ZN(_02912_ ) );
OAI21_X1 _18769_ ( .A(_02892_ ), .B1(_02912_ ), .B2(_02891_ ), .ZN(_02913_ ) );
MUX2_X1 _18770_ ( .A(\EXU.ls_rdata_i [7] ), .B(_02913_ ), .S(_02823_ ), .Z(_00956_ ) );
NOR2_X1 _18771_ ( .A1(_07759_ ), .A2(_02807_ ), .ZN(_02914_ ) );
OAI21_X1 _18772_ ( .A(_02914_ ), .B1(_02891_ ), .B2(_02864_ ), .ZN(_02915_ ) );
CLKBUF_X2 _18773_ ( .A(_04711_ ), .Z(_02916_ ) );
AND3_X1 _18774_ ( .A1(_02794_ ), .A2(_02916_ ), .A3(_02850_ ), .ZN(_02917_ ) );
BUF_X2 _18775_ ( .A(_04711_ ), .Z(_02918_ ) );
NOR2_X1 _18776_ ( .A1(_07793_ ), .A2(_02807_ ), .ZN(_02919_ ) );
NAND3_X1 _18777_ ( .A1(_02774_ ), .A2(_02918_ ), .A3(_02919_ ), .ZN(_02920_ ) );
AND3_X1 _18778_ ( .A1(_02777_ ), .A2(_04711_ ), .A3(_02803_ ), .ZN(_02921_ ) );
NAND2_X1 _18779_ ( .A1(_02897_ ), .A2(_02919_ ), .ZN(_02922_ ) );
OAI21_X1 _18780_ ( .A(_02914_ ), .B1(_02900_ ), .B2(_02831_ ), .ZN(_02923_ ) );
AND3_X1 _18781_ ( .A1(_02793_ ), .A2(_02902_ ), .A3(_02850_ ), .ZN(_02924_ ) );
AND2_X1 _18782_ ( .A1(_02777_ ), .A2(_05570_ ), .ZN(_02925_ ) );
AOI21_X1 _18783_ ( .A(_02924_ ), .B1(_02803_ ), .B2(_02925_ ), .ZN(_02926_ ) );
NAND3_X1 _18784_ ( .A1(_02922_ ), .A2(_02923_ ), .A3(_02926_ ), .ZN(_02927_ ) );
AOI21_X1 _18785_ ( .A(_02921_ ), .B1(_02927_ ), .B2(_02908_ ), .ZN(_02928_ ) );
OAI21_X1 _18786_ ( .A(_02920_ ), .B1(_02928_ ), .B2(_02791_ ), .ZN(_02929_ ) );
AOI21_X1 _18787_ ( .A(_02917_ ), .B1(_02929_ ), .B2(_02911_ ), .ZN(_02930_ ) );
OAI21_X1 _18788_ ( .A(_02915_ ), .B1(_02930_ ), .B2(_02891_ ), .ZN(_02931_ ) );
MUX2_X1 _18789_ ( .A(\EXU.ls_rdata_i [6] ), .B(_02931_ ), .S(_02823_ ), .Z(_00957_ ) );
NOR2_X1 _18790_ ( .A1(_07762_ ), .A2(_02807_ ), .ZN(_02932_ ) );
OAI21_X1 _18791_ ( .A(_02932_ ), .B1(_02786_ ), .B2(_02864_ ), .ZN(_02933_ ) );
AND3_X1 _18792_ ( .A1(_02794_ ), .A2(_02916_ ), .A3(_02856_ ), .ZN(_02934_ ) );
NAND3_X1 _18793_ ( .A1(_02774_ ), .A2(_02918_ ), .A3(_02808_ ), .ZN(_02935_ ) );
NOR2_X1 _18794_ ( .A1(_02908_ ), .A2(_02854_ ), .ZN(_02936_ ) );
NAND2_X1 _18795_ ( .A1(_02897_ ), .A2(_02808_ ), .ZN(_02937_ ) );
OAI21_X1 _18796_ ( .A(_02932_ ), .B1(_02900_ ), .B2(_02831_ ), .ZN(_02938_ ) );
INV_X1 _18797_ ( .A(_02925_ ), .ZN(_02939_ ) );
NOR2_X1 _18798_ ( .A1(_02939_ ), .A2(_02854_ ), .ZN(_02940_ ) );
AND3_X1 _18799_ ( .A1(_02794_ ), .A2(_02902_ ), .A3(_02856_ ), .ZN(_02941_ ) );
NOR2_X1 _18800_ ( .A1(_02940_ ), .A2(_02941_ ), .ZN(_02942_ ) );
NAND3_X1 _18801_ ( .A1(_02937_ ), .A2(_02938_ ), .A3(_02942_ ), .ZN(_02943_ ) );
AOI21_X1 _18802_ ( .A(_02936_ ), .B1(_02943_ ), .B2(_02908_ ), .ZN(_02944_ ) );
OAI21_X1 _18803_ ( .A(_02935_ ), .B1(_02944_ ), .B2(_02791_ ), .ZN(_02945_ ) );
AOI21_X1 _18804_ ( .A(_02934_ ), .B1(_02945_ ), .B2(_02911_ ), .ZN(_02946_ ) );
OAI21_X1 _18805_ ( .A(_02933_ ), .B1(_02946_ ), .B2(_02891_ ), .ZN(_02947_ ) );
MUX2_X1 _18806_ ( .A(\EXU.ls_rdata_i [5] ), .B(_02947_ ), .S(_02823_ ), .Z(_00958_ ) );
NAND2_X1 _18807_ ( .A1(_02897_ ), .A2(_02811_ ), .ZN(_02948_ ) );
NOR2_X1 _18808_ ( .A1(_07765_ ), .A2(_07831_ ), .ZN(_02949_ ) );
OAI21_X1 _18809_ ( .A(_02949_ ), .B1(_02900_ ), .B2(_02831_ ), .ZN(_02950_ ) );
AND3_X1 _18810_ ( .A1(_02793_ ), .A2(_02902_ ), .A3(_02861_ ), .ZN(_02951_ ) );
AOI21_X1 _18811_ ( .A(_02951_ ), .B1(_02859_ ), .B2(_02925_ ), .ZN(_02952_ ) );
NAND3_X1 _18812_ ( .A1(_02948_ ), .A2(_02950_ ), .A3(_02952_ ), .ZN(_02953_ ) );
NAND2_X1 _18813_ ( .A1(_02953_ ), .A2(_02908_ ), .ZN(_02954_ ) );
AND2_X1 _18814_ ( .A1(_02618_ ), .A2(_02622_ ), .ZN(_02955_ ) );
NAND4_X1 _18815_ ( .A1(_02955_ ), .A2(_02847_ ), .A3(_02916_ ), .A4(_02859_ ), .ZN(_02956_ ) );
AOI21_X1 _18816_ ( .A(_02791_ ), .B1(_02954_ ), .B2(_02956_ ), .ZN(_02957_ ) );
AND4_X1 _18817_ ( .A1(_02847_ ), .A2(_02655_ ), .A3(_02916_ ), .A4(_02811_ ), .ZN(_02958_ ) );
OAI21_X1 _18818_ ( .A(_02911_ ), .B1(_02957_ ), .B2(_02958_ ), .ZN(_02959_ ) );
NAND4_X1 _18819_ ( .A1(_02652_ ), .A2(_02847_ ), .A3(_02918_ ), .A4(_02861_ ), .ZN(_02960_ ) );
AOI21_X1 _18820_ ( .A(_02891_ ), .B1(_02959_ ), .B2(_02960_ ), .ZN(_02961_ ) );
OAI211_X1 _18821_ ( .A(_02798_ ), .B(_02949_ ), .C1(_02918_ ), .C2(_02800_ ), .ZN(_02962_ ) );
INV_X1 _18822_ ( .A(_02962_ ), .ZN(_02963_ ) );
OAI21_X1 _18823_ ( .A(_02647_ ), .B1(_02961_ ), .B2(_02963_ ), .ZN(_02964_ ) );
OAI21_X1 _18824_ ( .A(_02964_ ), .B1(_07095_ ), .B2(\LSU.ls_axi_rready_$_ANDNOT__A_Y ), .ZN(_00959_ ) );
NAND2_X1 _18825_ ( .A1(_02897_ ), .A2(_02814_ ), .ZN(_02965_ ) );
NOR2_X1 _18826_ ( .A1(_07769_ ), .A2(_02807_ ), .ZN(_02966_ ) );
OAI21_X1 _18827_ ( .A(_02966_ ), .B1(_02900_ ), .B2(_02831_ ), .ZN(_02967_ ) );
NAND3_X1 _18828_ ( .A1(_02777_ ), .A2(_02902_ ), .A3(_02868_ ), .ZN(_02968_ ) );
NAND3_X1 _18829_ ( .A1(_02794_ ), .A2(_02902_ ), .A3(_02871_ ), .ZN(_02969_ ) );
AND2_X1 _18830_ ( .A1(_02968_ ), .A2(_02969_ ), .ZN(_02970_ ) );
NAND3_X1 _18831_ ( .A1(_02965_ ), .A2(_02967_ ), .A3(_02970_ ), .ZN(_02971_ ) );
NAND2_X1 _18832_ ( .A1(_02971_ ), .A2(_02908_ ), .ZN(_02972_ ) );
NAND4_X1 _18833_ ( .A1(_02955_ ), .A2(_02847_ ), .A3(_02916_ ), .A4(_02868_ ), .ZN(_02973_ ) );
AOI21_X1 _18834_ ( .A(_02791_ ), .B1(_02972_ ), .B2(_02973_ ), .ZN(_02974_ ) );
AND4_X1 _18835_ ( .A1(_02847_ ), .A2(_02655_ ), .A3(_02916_ ), .A4(_02814_ ), .ZN(_02975_ ) );
OAI21_X1 _18836_ ( .A(_02911_ ), .B1(_02974_ ), .B2(_02975_ ), .ZN(_02976_ ) );
NAND4_X1 _18837_ ( .A1(_02652_ ), .A2(_02847_ ), .A3(_02918_ ), .A4(_02871_ ), .ZN(_02977_ ) );
AOI21_X1 _18838_ ( .A(_02891_ ), .B1(_02976_ ), .B2(_02977_ ), .ZN(_02978_ ) );
OAI211_X1 _18839_ ( .A(_02798_ ), .B(_02966_ ), .C1(_02918_ ), .C2(_02800_ ), .ZN(_02979_ ) );
INV_X1 _18840_ ( .A(_02979_ ), .ZN(_02980_ ) );
OAI21_X1 _18841_ ( .A(_02647_ ), .B1(_02978_ ), .B2(_02980_ ), .ZN(_02981_ ) );
OAI21_X1 _18842_ ( .A(_02981_ ), .B1(_07140_ ), .B2(\LSU.ls_axi_rready_$_ANDNOT__A_Y ), .ZN(_00960_ ) );
NOR2_X1 _18843_ ( .A1(_07772_ ), .A2(_02807_ ), .ZN(_02982_ ) );
OAI21_X1 _18844_ ( .A(_02982_ ), .B1(_02786_ ), .B2(_02864_ ), .ZN(_02983_ ) );
AND3_X1 _18845_ ( .A1(_02794_ ), .A2(_02916_ ), .A3(_02876_ ), .ZN(_02984_ ) );
NAND3_X1 _18846_ ( .A1(_02774_ ), .A2(_02918_ ), .A3(_02817_ ), .ZN(_02985_ ) );
NOR2_X1 _18847_ ( .A1(_02908_ ), .A2(_02874_ ), .ZN(_02986_ ) );
NAND2_X1 _18848_ ( .A1(_02897_ ), .A2(_02817_ ), .ZN(_02987_ ) );
OAI21_X1 _18849_ ( .A(_02982_ ), .B1(_02900_ ), .B2(_02830_ ), .ZN(_02988_ ) );
NOR2_X1 _18850_ ( .A1(_02939_ ), .A2(_02874_ ), .ZN(_02989_ ) );
AND3_X1 _18851_ ( .A1(_02793_ ), .A2(_02902_ ), .A3(_02876_ ), .ZN(_02990_ ) );
NOR2_X1 _18852_ ( .A1(_02989_ ), .A2(_02990_ ), .ZN(_02991_ ) );
NAND3_X1 _18853_ ( .A1(_02987_ ), .A2(_02988_ ), .A3(_02991_ ), .ZN(_02992_ ) );
AOI21_X1 _18854_ ( .A(_02986_ ), .B1(_02992_ ), .B2(_02908_ ), .ZN(_02993_ ) );
OAI21_X1 _18855_ ( .A(_02985_ ), .B1(_02993_ ), .B2(_02791_ ), .ZN(_02994_ ) );
AOI21_X1 _18856_ ( .A(_02984_ ), .B1(_02994_ ), .B2(_02911_ ), .ZN(_02995_ ) );
OAI21_X1 _18857_ ( .A(_02983_ ), .B1(_02995_ ), .B2(_02891_ ), .ZN(_02996_ ) );
BUF_X4 _18858_ ( .A(_02646_ ), .Z(_02997_ ) );
MUX2_X1 _18859_ ( .A(\EXU.ls_rdata_i [2] ), .B(_02996_ ), .S(_02997_ ), .Z(_00961_ ) );
NAND3_X1 _18860_ ( .A1(_02781_ ), .A2(_02799_ ), .A3(_02859_ ), .ZN(_02998_ ) );
NAND4_X1 _18861_ ( .A1(_02785_ ), .A2(_02789_ ), .A3(_02797_ ), .A4(_02998_ ), .ZN(_02999_ ) );
MUX2_X1 _18862_ ( .A(\EXU.ls_rdata_i [28] ), .B(_02999_ ), .S(_02997_ ), .Z(_00962_ ) );
NOR2_X1 _18863_ ( .A1(_02786_ ), .A2(_02864_ ), .ZN(_03000_ ) );
INV_X1 _18864_ ( .A(_04089_ ), .ZN(_03001_ ) );
INV_X1 _18865_ ( .A(_04074_ ), .ZN(_03002_ ) );
INV_X1 _18866_ ( .A(_04098_ ), .ZN(_03003_ ) );
AOI211_X1 _18867_ ( .A(_04201_ ), .B(_03001_ ), .C1(_03002_ ), .C2(_03003_ ), .ZN(_03004_ ) );
AOI21_X1 _18868_ ( .A(_03004_ ), .B1(\io_master_rdata [1] ), .B2(_07540_ ), .ZN(_03005_ ) );
OR2_X1 _18869_ ( .A1(_03005_ ), .A2(_02806_ ), .ZN(_03006_ ) );
OR2_X1 _18870_ ( .A1(_03000_ ), .A2(_03006_ ), .ZN(_03007_ ) );
AND3_X1 _18871_ ( .A1(_02794_ ), .A2(_02916_ ), .A3(_02882_ ), .ZN(_03008_ ) );
NAND3_X1 _18872_ ( .A1(_02774_ ), .A2(_02918_ ), .A3(_02820_ ), .ZN(_03009_ ) );
NOR2_X1 _18873_ ( .A1(_02907_ ), .A2(_02880_ ), .ZN(_03010_ ) );
NAND2_X1 _18874_ ( .A1(_02897_ ), .A2(_02820_ ), .ZN(_03011_ ) );
NOR2_X1 _18875_ ( .A1(_02900_ ), .A2(_02830_ ), .ZN(_03012_ ) );
OR2_X1 _18876_ ( .A1(_03012_ ), .A2(_03006_ ), .ZN(_03013_ ) );
NAND3_X1 _18877_ ( .A1(_02794_ ), .A2(_02902_ ), .A3(_02882_ ), .ZN(_03014_ ) );
OR2_X1 _18878_ ( .A1(_02939_ ), .A2(_02880_ ), .ZN(_03015_ ) );
NAND4_X1 _18879_ ( .A1(_03011_ ), .A2(_03013_ ), .A3(_03014_ ), .A4(_03015_ ), .ZN(_03016_ ) );
AOI21_X1 _18880_ ( .A(_03010_ ), .B1(_03016_ ), .B2(_02908_ ), .ZN(_03017_ ) );
OAI21_X1 _18881_ ( .A(_03009_ ), .B1(_03017_ ), .B2(_02791_ ), .ZN(_03018_ ) );
AOI21_X1 _18882_ ( .A(_03008_ ), .B1(_03018_ ), .B2(_02911_ ), .ZN(_03019_ ) );
OAI21_X1 _18883_ ( .A(_03007_ ), .B1(_03019_ ), .B2(_02891_ ), .ZN(_03020_ ) );
MUX2_X1 _18884_ ( .A(\EXU.ls_rdata_i [1] ), .B(_03020_ ), .S(_02997_ ), .Z(_00963_ ) );
AND3_X1 _18885_ ( .A1(_02794_ ), .A2(_02916_ ), .A3(_02887_ ), .ZN(_03021_ ) );
NAND3_X1 _18886_ ( .A1(_02774_ ), .A2(_02916_ ), .A3(_02824_ ), .ZN(_03022_ ) );
NOR2_X1 _18887_ ( .A1(_02907_ ), .A2(_02885_ ), .ZN(_03023_ ) );
NAND2_X1 _18888_ ( .A1(_02897_ ), .A2(_02824_ ), .ZN(_03024_ ) );
AOI211_X1 _18889_ ( .A(_04206_ ), .B(_03001_ ), .C1(_03002_ ), .C2(_03003_ ), .ZN(_03025_ ) );
AOI21_X1 _18890_ ( .A(_03025_ ), .B1(\io_master_rdata [0] ), .B2(_07540_ ), .ZN(_03026_ ) );
OR2_X1 _18891_ ( .A1(_03026_ ), .A2(_04105_ ), .ZN(_03027_ ) );
OR2_X1 _18892_ ( .A1(_03012_ ), .A2(_03027_ ), .ZN(_03028_ ) );
NOR2_X1 _18893_ ( .A1(_02939_ ), .A2(_02885_ ), .ZN(_03029_ ) );
AND3_X1 _18894_ ( .A1(_02793_ ), .A2(_02902_ ), .A3(_02887_ ), .ZN(_03030_ ) );
NOR2_X1 _18895_ ( .A1(_03029_ ), .A2(_03030_ ), .ZN(_03031_ ) );
NAND3_X1 _18896_ ( .A1(_03024_ ), .A2(_03028_ ), .A3(_03031_ ), .ZN(_03032_ ) );
AOI21_X1 _18897_ ( .A(_03023_ ), .B1(_03032_ ), .B2(_02908_ ), .ZN(_03033_ ) );
OAI21_X1 _18898_ ( .A(_03022_ ), .B1(_03033_ ), .B2(_02791_ ), .ZN(_03034_ ) );
AOI21_X1 _18899_ ( .A(_03021_ ), .B1(_03034_ ), .B2(_02911_ ), .ZN(_03035_ ) );
OAI22_X1 _18900_ ( .A1(_03035_ ), .A2(_02891_ ), .B1(_03000_ ), .B2(_03027_ ), .ZN(_03036_ ) );
MUX2_X1 _18901_ ( .A(\EXU.ls_rdata_i [0] ), .B(_03036_ ), .S(_02997_ ), .Z(_00964_ ) );
NAND3_X1 _18902_ ( .A1(_02781_ ), .A2(_02799_ ), .A3(_02868_ ), .ZN(_03037_ ) );
NAND4_X1 _18903_ ( .A1(_02784_ ), .A2(_02789_ ), .A3(_02797_ ), .A4(_03037_ ), .ZN(_03038_ ) );
MUX2_X1 _18904_ ( .A(\EXU.ls_rdata_i [27] ), .B(_03038_ ), .S(_02997_ ), .Z(_00965_ ) );
OR2_X1 _18905_ ( .A1(_02865_ ), .A2(_02874_ ), .ZN(_03039_ ) );
NAND4_X1 _18906_ ( .A1(_02784_ ), .A2(_03039_ ), .A3(_02788_ ), .A4(_02796_ ), .ZN(_03040_ ) );
MUX2_X1 _18907_ ( .A(\EXU.ls_rdata_i [26] ), .B(_03040_ ), .S(_02997_ ), .Z(_00966_ ) );
OR2_X1 _18908_ ( .A1(_02865_ ), .A2(_02880_ ), .ZN(_03041_ ) );
NAND4_X1 _18909_ ( .A1(_02784_ ), .A2(_03041_ ), .A3(_02788_ ), .A4(_02796_ ), .ZN(_03042_ ) );
MUX2_X1 _18910_ ( .A(\EXU.ls_rdata_i [25] ), .B(_03042_ ), .S(_02997_ ), .Z(_00967_ ) );
OR2_X1 _18911_ ( .A1(_02865_ ), .A2(_02885_ ), .ZN(_03043_ ) );
NAND4_X1 _18912_ ( .A1(_02784_ ), .A2(_03043_ ), .A3(_02788_ ), .A4(_02796_ ), .ZN(_03044_ ) );
MUX2_X1 _18913_ ( .A(\EXU.ls_rdata_i [24] ), .B(_03044_ ), .S(_02997_ ), .Z(_00968_ ) );
NAND3_X1 _18914_ ( .A1(_02781_ ), .A2(_02799_ ), .A3(_02792_ ), .ZN(_03045_ ) );
NAND4_X1 _18915_ ( .A1(_02784_ ), .A2(_02788_ ), .A3(_02796_ ), .A4(_03045_ ), .ZN(_03046_ ) );
MUX2_X1 _18916_ ( .A(\EXU.ls_rdata_i [23] ), .B(_03046_ ), .S(_02997_ ), .Z(_00969_ ) );
NAND3_X1 _18917_ ( .A1(_02781_ ), .A2(_02799_ ), .A3(_02919_ ), .ZN(_03047_ ) );
NAND4_X1 _18918_ ( .A1(_02784_ ), .A2(_02788_ ), .A3(_02796_ ), .A4(_03047_ ), .ZN(_03048_ ) );
MUX2_X1 _18919_ ( .A(\EXU.ls_rdata_i [22] ), .B(_03048_ ), .S(_02997_ ), .Z(_00970_ ) );
INV_X1 _18920_ ( .A(_05436_ ), .ZN(_03049_ ) );
AND2_X2 _18921_ ( .A1(_03049_ ), .A2(\EXU.gpr_wen_o ), .ZN(_03050_ ) );
BUF_X4 _18922_ ( .A(_03050_ ), .Z(_03051_ ) );
AND4_X1 _18923_ ( .A1(\EXU.rd_o [3] ), .A2(_05430_ ), .A3(_05434_ ), .A4(\EXU.rd_o [1] ), .ZN(_03052_ ) );
AND2_X2 _18924_ ( .A1(_03051_ ), .A2(_03052_ ), .ZN(_03053_ ) );
BUF_X4 _18925_ ( .A(_03053_ ), .Z(_03054_ ) );
MUX2_X1 _18926_ ( .A(\RFU.rf[10][31] ), .B(\EXU.xrd_o [31] ), .S(_03054_ ), .Z(_00971_ ) );
MUX2_X1 _18927_ ( .A(\RFU.rf[10][30] ), .B(\EXU.xrd_o [30] ), .S(_03054_ ), .Z(_00972_ ) );
MUX2_X1 _18928_ ( .A(\RFU.rf[10][21] ), .B(\EXU.xrd_o [21] ), .S(_03054_ ), .Z(_00973_ ) );
MUX2_X1 _18929_ ( .A(\RFU.rf[10][20] ), .B(\EXU.xrd_o [20] ), .S(_03054_ ), .Z(_00974_ ) );
MUX2_X1 _18930_ ( .A(\RFU.rf[10][19] ), .B(\EXU.xrd_o [19] ), .S(_03054_ ), .Z(_00975_ ) );
MUX2_X1 _18931_ ( .A(\RFU.rf[10][18] ), .B(\EXU.xrd_o [18] ), .S(_03054_ ), .Z(_00976_ ) );
MUX2_X1 _18932_ ( .A(\RFU.rf[10][17] ), .B(\EXU.xrd_o [17] ), .S(_03054_ ), .Z(_00977_ ) );
MUX2_X1 _18933_ ( .A(\RFU.rf[10][16] ), .B(\EXU.xrd_o [16] ), .S(_03054_ ), .Z(_00978_ ) );
MUX2_X1 _18934_ ( .A(\RFU.rf[10][15] ), .B(\EXU.xrd_o [15] ), .S(_03054_ ), .Z(_00979_ ) );
MUX2_X1 _18935_ ( .A(\RFU.rf[10][14] ), .B(\EXU.xrd_o [14] ), .S(_03054_ ), .Z(_00980_ ) );
BUF_X4 _18936_ ( .A(_03053_ ), .Z(_03055_ ) );
MUX2_X1 _18937_ ( .A(\RFU.rf[10][13] ), .B(\EXU.xrd_o [13] ), .S(_03055_ ), .Z(_00981_ ) );
MUX2_X1 _18938_ ( .A(\RFU.rf[10][12] ), .B(\EXU.xrd_o [12] ), .S(_03055_ ), .Z(_00982_ ) );
MUX2_X1 _18939_ ( .A(\RFU.rf[10][29] ), .B(\EXU.xrd_o [29] ), .S(_03055_ ), .Z(_00983_ ) );
MUX2_X1 _18940_ ( .A(\RFU.rf[10][11] ), .B(\EXU.xrd_o [11] ), .S(_03055_ ), .Z(_00984_ ) );
MUX2_X1 _18941_ ( .A(\RFU.rf[10][10] ), .B(\EXU.xrd_o [10] ), .S(_03055_ ), .Z(_00985_ ) );
MUX2_X1 _18942_ ( .A(\RFU.rf[10][9] ), .B(\EXU.xrd_o [9] ), .S(_03055_ ), .Z(_00986_ ) );
MUX2_X1 _18943_ ( .A(\RFU.rf[10][8] ), .B(\EXU.xrd_o [8] ), .S(_03055_ ), .Z(_00987_ ) );
MUX2_X1 _18944_ ( .A(\RFU.rf[10][7] ), .B(\EXU.xrd_o [7] ), .S(_03055_ ), .Z(_00988_ ) );
MUX2_X1 _18945_ ( .A(\RFU.rf[10][6] ), .B(\EXU.xrd_o [6] ), .S(_03055_ ), .Z(_00989_ ) );
MUX2_X1 _18946_ ( .A(\RFU.rf[10][5] ), .B(\EXU.xrd_o [5] ), .S(_03055_ ), .Z(_00990_ ) );
BUF_X4 _18947_ ( .A(_03053_ ), .Z(_03056_ ) );
MUX2_X1 _18948_ ( .A(\RFU.rf[10][4] ), .B(\EXU.xrd_o [4] ), .S(_03056_ ), .Z(_00991_ ) );
MUX2_X1 _18949_ ( .A(\RFU.rf[10][3] ), .B(\EXU.xrd_o [3] ), .S(_03056_ ), .Z(_00992_ ) );
MUX2_X1 _18950_ ( .A(\RFU.rf[10][2] ), .B(\EXU.xrd_o [2] ), .S(_03056_ ), .Z(_00993_ ) );
MUX2_X1 _18951_ ( .A(\RFU.rf[10][28] ), .B(\EXU.xrd_o [28] ), .S(_03056_ ), .Z(_00994_ ) );
MUX2_X1 _18952_ ( .A(\RFU.rf[10][1] ), .B(\EXU.xrd_o [1] ), .S(_03056_ ), .Z(_00995_ ) );
MUX2_X1 _18953_ ( .A(\RFU.rf[10][0] ), .B(\EXU.xrd_o [0] ), .S(_03056_ ), .Z(_00996_ ) );
MUX2_X1 _18954_ ( .A(\RFU.rf[10][27] ), .B(\EXU.xrd_o [27] ), .S(_03056_ ), .Z(_00997_ ) );
MUX2_X1 _18955_ ( .A(\RFU.rf[10][26] ), .B(\EXU.xrd_o [26] ), .S(_03056_ ), .Z(_00998_ ) );
MUX2_X1 _18956_ ( .A(\RFU.rf[10][25] ), .B(\EXU.xrd_o [25] ), .S(_03056_ ), .Z(_00999_ ) );
MUX2_X1 _18957_ ( .A(\RFU.rf[10][24] ), .B(\EXU.xrd_o [24] ), .S(_03056_ ), .Z(_01000_ ) );
MUX2_X1 _18958_ ( .A(\RFU.rf[10][23] ), .B(\EXU.xrd_o [23] ), .S(_03053_ ), .Z(_01001_ ) );
MUX2_X1 _18959_ ( .A(\RFU.rf[10][22] ), .B(\EXU.xrd_o [22] ), .S(_03053_ ), .Z(_01002_ ) );
AND4_X1 _18960_ ( .A1(\EXU.rd_o [3] ), .A2(_05430_ ), .A3(\EXU.rd_o [1] ), .A4(\EXU.rd_o [0] ), .ZN(_03057_ ) );
AND2_X2 _18961_ ( .A1(_03051_ ), .A2(_03057_ ), .ZN(_03058_ ) );
BUF_X4 _18962_ ( .A(_03058_ ), .Z(_03059_ ) );
MUX2_X1 _18963_ ( .A(\RFU.rf[11][31] ), .B(\EXU.xrd_o [31] ), .S(_03059_ ), .Z(_01003_ ) );
MUX2_X1 _18964_ ( .A(\RFU.rf[11][30] ), .B(\EXU.xrd_o [30] ), .S(_03059_ ), .Z(_01004_ ) );
MUX2_X1 _18965_ ( .A(\RFU.rf[11][21] ), .B(\EXU.xrd_o [21] ), .S(_03059_ ), .Z(_01005_ ) );
MUX2_X1 _18966_ ( .A(\RFU.rf[11][20] ), .B(\EXU.xrd_o [20] ), .S(_03059_ ), .Z(_01006_ ) );
MUX2_X1 _18967_ ( .A(\RFU.rf[11][19] ), .B(\EXU.xrd_o [19] ), .S(_03059_ ), .Z(_01007_ ) );
MUX2_X1 _18968_ ( .A(\RFU.rf[11][18] ), .B(\EXU.xrd_o [18] ), .S(_03059_ ), .Z(_01008_ ) );
MUX2_X1 _18969_ ( .A(\RFU.rf[11][17] ), .B(\EXU.xrd_o [17] ), .S(_03059_ ), .Z(_01009_ ) );
MUX2_X1 _18970_ ( .A(\RFU.rf[11][16] ), .B(\EXU.xrd_o [16] ), .S(_03059_ ), .Z(_01010_ ) );
MUX2_X1 _18971_ ( .A(\RFU.rf[11][15] ), .B(\EXU.xrd_o [15] ), .S(_03059_ ), .Z(_01011_ ) );
MUX2_X1 _18972_ ( .A(\RFU.rf[11][14] ), .B(\EXU.xrd_o [14] ), .S(_03059_ ), .Z(_01012_ ) );
BUF_X4 _18973_ ( .A(_03058_ ), .Z(_03060_ ) );
MUX2_X1 _18974_ ( .A(\RFU.rf[11][13] ), .B(\EXU.xrd_o [13] ), .S(_03060_ ), .Z(_01013_ ) );
MUX2_X1 _18975_ ( .A(\RFU.rf[11][12] ), .B(\EXU.xrd_o [12] ), .S(_03060_ ), .Z(_01014_ ) );
MUX2_X1 _18976_ ( .A(\RFU.rf[11][29] ), .B(\EXU.xrd_o [29] ), .S(_03060_ ), .Z(_01015_ ) );
MUX2_X1 _18977_ ( .A(\RFU.rf[11][11] ), .B(\EXU.xrd_o [11] ), .S(_03060_ ), .Z(_01016_ ) );
MUX2_X1 _18978_ ( .A(\RFU.rf[11][10] ), .B(\EXU.xrd_o [10] ), .S(_03060_ ), .Z(_01017_ ) );
MUX2_X1 _18979_ ( .A(\RFU.rf[11][9] ), .B(\EXU.xrd_o [9] ), .S(_03060_ ), .Z(_01018_ ) );
MUX2_X1 _18980_ ( .A(\RFU.rf[11][8] ), .B(\EXU.xrd_o [8] ), .S(_03060_ ), .Z(_01019_ ) );
MUX2_X1 _18981_ ( .A(\RFU.rf[11][7] ), .B(\EXU.xrd_o [7] ), .S(_03060_ ), .Z(_01020_ ) );
MUX2_X1 _18982_ ( .A(\RFU.rf[11][6] ), .B(\EXU.xrd_o [6] ), .S(_03060_ ), .Z(_01021_ ) );
MUX2_X1 _18983_ ( .A(\RFU.rf[11][5] ), .B(\EXU.xrd_o [5] ), .S(_03060_ ), .Z(_01022_ ) );
BUF_X4 _18984_ ( .A(_03058_ ), .Z(_03061_ ) );
MUX2_X1 _18985_ ( .A(\RFU.rf[11][4] ), .B(\EXU.xrd_o [4] ), .S(_03061_ ), .Z(_01023_ ) );
MUX2_X1 _18986_ ( .A(\RFU.rf[11][3] ), .B(\EXU.xrd_o [3] ), .S(_03061_ ), .Z(_01024_ ) );
MUX2_X1 _18987_ ( .A(\RFU.rf[11][2] ), .B(\EXU.xrd_o [2] ), .S(_03061_ ), .Z(_01025_ ) );
MUX2_X1 _18988_ ( .A(\RFU.rf[11][28] ), .B(\EXU.xrd_o [28] ), .S(_03061_ ), .Z(_01026_ ) );
MUX2_X1 _18989_ ( .A(\RFU.rf[11][1] ), .B(\EXU.xrd_o [1] ), .S(_03061_ ), .Z(_01027_ ) );
MUX2_X1 _18990_ ( .A(\RFU.rf[11][0] ), .B(\EXU.xrd_o [0] ), .S(_03061_ ), .Z(_01028_ ) );
MUX2_X1 _18991_ ( .A(\RFU.rf[11][27] ), .B(\EXU.xrd_o [27] ), .S(_03061_ ), .Z(_01029_ ) );
MUX2_X1 _18992_ ( .A(\RFU.rf[11][26] ), .B(\EXU.xrd_o [26] ), .S(_03061_ ), .Z(_01030_ ) );
MUX2_X1 _18993_ ( .A(\RFU.rf[11][25] ), .B(\EXU.xrd_o [25] ), .S(_03061_ ), .Z(_01031_ ) );
MUX2_X1 _18994_ ( .A(\RFU.rf[11][24] ), .B(\EXU.xrd_o [24] ), .S(_03061_ ), .Z(_01032_ ) );
MUX2_X1 _18995_ ( .A(\RFU.rf[11][23] ), .B(\EXU.xrd_o [23] ), .S(_03058_ ), .Z(_01033_ ) );
MUX2_X1 _18996_ ( .A(\RFU.rf[11][22] ), .B(\EXU.xrd_o [22] ), .S(_03058_ ), .Z(_01034_ ) );
AND4_X1 _18997_ ( .A1(\EXU.rd_o [3] ), .A2(_05432_ ), .A3(_05434_ ), .A4(\EXU.rd_o [2] ), .ZN(_03062_ ) );
NAND2_X1 _18998_ ( .A1(_03051_ ), .A2(_03062_ ), .ZN(_03063_ ) );
BUF_X4 _18999_ ( .A(_03063_ ), .Z(_03064_ ) );
MUX2_X1 _19000_ ( .A(\EXU.xrd_o [31] ), .B(\RFU.rf[12][31] ), .S(_03064_ ), .Z(_01035_ ) );
MUX2_X1 _19001_ ( .A(\EXU.xrd_o [30] ), .B(\RFU.rf[12][30] ), .S(_03064_ ), .Z(_01036_ ) );
MUX2_X1 _19002_ ( .A(\EXU.xrd_o [21] ), .B(\RFU.rf[12][21] ), .S(_03064_ ), .Z(_01037_ ) );
MUX2_X1 _19003_ ( .A(\EXU.xrd_o [20] ), .B(\RFU.rf[12][20] ), .S(_03064_ ), .Z(_01038_ ) );
MUX2_X1 _19004_ ( .A(\EXU.xrd_o [19] ), .B(\RFU.rf[12][19] ), .S(_03064_ ), .Z(_01039_ ) );
MUX2_X1 _19005_ ( .A(\EXU.xrd_o [18] ), .B(\RFU.rf[12][18] ), .S(_03064_ ), .Z(_01040_ ) );
MUX2_X1 _19006_ ( .A(\EXU.xrd_o [17] ), .B(\RFU.rf[12][17] ), .S(_03064_ ), .Z(_01041_ ) );
MUX2_X1 _19007_ ( .A(\EXU.xrd_o [16] ), .B(\RFU.rf[12][16] ), .S(_03064_ ), .Z(_01042_ ) );
MUX2_X1 _19008_ ( .A(\EXU.xrd_o [15] ), .B(\RFU.rf[12][15] ), .S(_03064_ ), .Z(_01043_ ) );
MUX2_X1 _19009_ ( .A(\EXU.xrd_o [14] ), .B(\RFU.rf[12][14] ), .S(_03064_ ), .Z(_01044_ ) );
BUF_X4 _19010_ ( .A(_03063_ ), .Z(_03065_ ) );
MUX2_X1 _19011_ ( .A(\EXU.xrd_o [13] ), .B(\RFU.rf[12][13] ), .S(_03065_ ), .Z(_01045_ ) );
MUX2_X1 _19012_ ( .A(\EXU.xrd_o [12] ), .B(\RFU.rf[12][12] ), .S(_03065_ ), .Z(_01046_ ) );
MUX2_X1 _19013_ ( .A(\EXU.xrd_o [29] ), .B(\RFU.rf[12][29] ), .S(_03065_ ), .Z(_01047_ ) );
MUX2_X1 _19014_ ( .A(\EXU.xrd_o [11] ), .B(\RFU.rf[12][11] ), .S(_03065_ ), .Z(_01048_ ) );
MUX2_X1 _19015_ ( .A(\EXU.xrd_o [10] ), .B(\RFU.rf[12][10] ), .S(_03065_ ), .Z(_01049_ ) );
MUX2_X1 _19016_ ( .A(\EXU.xrd_o [9] ), .B(\RFU.rf[12][9] ), .S(_03065_ ), .Z(_01050_ ) );
MUX2_X1 _19017_ ( .A(\EXU.xrd_o [8] ), .B(\RFU.rf[12][8] ), .S(_03065_ ), .Z(_01051_ ) );
MUX2_X1 _19018_ ( .A(\EXU.xrd_o [7] ), .B(\RFU.rf[12][7] ), .S(_03065_ ), .Z(_01052_ ) );
MUX2_X1 _19019_ ( .A(\EXU.xrd_o [6] ), .B(\RFU.rf[12][6] ), .S(_03065_ ), .Z(_01053_ ) );
MUX2_X1 _19020_ ( .A(\EXU.xrd_o [5] ), .B(\RFU.rf[12][5] ), .S(_03065_ ), .Z(_01054_ ) );
BUF_X4 _19021_ ( .A(_03063_ ), .Z(_03066_ ) );
MUX2_X1 _19022_ ( .A(\EXU.xrd_o [4] ), .B(\RFU.rf[12][4] ), .S(_03066_ ), .Z(_01055_ ) );
MUX2_X1 _19023_ ( .A(\EXU.xrd_o [3] ), .B(\RFU.rf[12][3] ), .S(_03066_ ), .Z(_01056_ ) );
MUX2_X1 _19024_ ( .A(\EXU.xrd_o [2] ), .B(\RFU.rf[12][2] ), .S(_03066_ ), .Z(_01057_ ) );
MUX2_X1 _19025_ ( .A(\EXU.xrd_o [28] ), .B(\RFU.rf[12][28] ), .S(_03066_ ), .Z(_01058_ ) );
MUX2_X1 _19026_ ( .A(\EXU.xrd_o [1] ), .B(\RFU.rf[12][1] ), .S(_03066_ ), .Z(_01059_ ) );
MUX2_X1 _19027_ ( .A(\EXU.xrd_o [0] ), .B(\RFU.rf[12][0] ), .S(_03066_ ), .Z(_01060_ ) );
MUX2_X1 _19028_ ( .A(\EXU.xrd_o [27] ), .B(\RFU.rf[12][27] ), .S(_03066_ ), .Z(_01061_ ) );
MUX2_X1 _19029_ ( .A(\EXU.xrd_o [26] ), .B(\RFU.rf[12][26] ), .S(_03066_ ), .Z(_01062_ ) );
MUX2_X1 _19030_ ( .A(\EXU.xrd_o [25] ), .B(\RFU.rf[12][25] ), .S(_03066_ ), .Z(_01063_ ) );
MUX2_X1 _19031_ ( .A(\EXU.xrd_o [24] ), .B(\RFU.rf[12][24] ), .S(_03066_ ), .Z(_01064_ ) );
MUX2_X1 _19032_ ( .A(\EXU.xrd_o [23] ), .B(\RFU.rf[12][23] ), .S(_03063_ ), .Z(_01065_ ) );
MUX2_X1 _19033_ ( .A(\EXU.xrd_o [22] ), .B(\RFU.rf[12][22] ), .S(_03063_ ), .Z(_01066_ ) );
AND4_X1 _19034_ ( .A1(\EXU.rd_o [3] ), .A2(_05432_ ), .A3(\EXU.rd_o [2] ), .A4(\EXU.rd_o [0] ), .ZN(_03067_ ) );
AND2_X2 _19035_ ( .A1(_03051_ ), .A2(_03067_ ), .ZN(_03068_ ) );
BUF_X4 _19036_ ( .A(_03068_ ), .Z(_03069_ ) );
MUX2_X1 _19037_ ( .A(\RFU.rf[13][31] ), .B(\EXU.xrd_o [31] ), .S(_03069_ ), .Z(_01067_ ) );
MUX2_X1 _19038_ ( .A(\RFU.rf[13][30] ), .B(\EXU.xrd_o [30] ), .S(_03069_ ), .Z(_01068_ ) );
MUX2_X1 _19039_ ( .A(\RFU.rf[13][21] ), .B(\EXU.xrd_o [21] ), .S(_03069_ ), .Z(_01069_ ) );
MUX2_X1 _19040_ ( .A(\RFU.rf[13][20] ), .B(\EXU.xrd_o [20] ), .S(_03069_ ), .Z(_01070_ ) );
MUX2_X1 _19041_ ( .A(\RFU.rf[13][19] ), .B(\EXU.xrd_o [19] ), .S(_03069_ ), .Z(_01071_ ) );
MUX2_X1 _19042_ ( .A(\RFU.rf[13][18] ), .B(\EXU.xrd_o [18] ), .S(_03069_ ), .Z(_01072_ ) );
MUX2_X1 _19043_ ( .A(\RFU.rf[13][17] ), .B(\EXU.xrd_o [17] ), .S(_03069_ ), .Z(_01073_ ) );
MUX2_X1 _19044_ ( .A(\RFU.rf[13][16] ), .B(\EXU.xrd_o [16] ), .S(_03069_ ), .Z(_01074_ ) );
MUX2_X1 _19045_ ( .A(\RFU.rf[13][15] ), .B(\EXU.xrd_o [15] ), .S(_03069_ ), .Z(_01075_ ) );
MUX2_X1 _19046_ ( .A(\RFU.rf[13][14] ), .B(\EXU.xrd_o [14] ), .S(_03069_ ), .Z(_01076_ ) );
BUF_X4 _19047_ ( .A(_03068_ ), .Z(_03070_ ) );
MUX2_X1 _19048_ ( .A(\RFU.rf[13][13] ), .B(\EXU.xrd_o [13] ), .S(_03070_ ), .Z(_01077_ ) );
MUX2_X1 _19049_ ( .A(\RFU.rf[13][12] ), .B(\EXU.xrd_o [12] ), .S(_03070_ ), .Z(_01078_ ) );
MUX2_X1 _19050_ ( .A(\RFU.rf[13][29] ), .B(\EXU.xrd_o [29] ), .S(_03070_ ), .Z(_01079_ ) );
MUX2_X1 _19051_ ( .A(\RFU.rf[13][11] ), .B(\EXU.xrd_o [11] ), .S(_03070_ ), .Z(_01080_ ) );
MUX2_X1 _19052_ ( .A(\RFU.rf[13][10] ), .B(\EXU.xrd_o [10] ), .S(_03070_ ), .Z(_01081_ ) );
MUX2_X1 _19053_ ( .A(\RFU.rf[13][9] ), .B(\EXU.xrd_o [9] ), .S(_03070_ ), .Z(_01082_ ) );
MUX2_X1 _19054_ ( .A(\RFU.rf[13][8] ), .B(\EXU.xrd_o [8] ), .S(_03070_ ), .Z(_01083_ ) );
MUX2_X1 _19055_ ( .A(\RFU.rf[13][7] ), .B(\EXU.xrd_o [7] ), .S(_03070_ ), .Z(_01084_ ) );
MUX2_X1 _19056_ ( .A(\RFU.rf[13][6] ), .B(\EXU.xrd_o [6] ), .S(_03070_ ), .Z(_01085_ ) );
MUX2_X1 _19057_ ( .A(\RFU.rf[13][5] ), .B(\EXU.xrd_o [5] ), .S(_03070_ ), .Z(_01086_ ) );
BUF_X4 _19058_ ( .A(_03068_ ), .Z(_03071_ ) );
MUX2_X1 _19059_ ( .A(\RFU.rf[13][4] ), .B(\EXU.xrd_o [4] ), .S(_03071_ ), .Z(_01087_ ) );
MUX2_X1 _19060_ ( .A(\RFU.rf[13][3] ), .B(\EXU.xrd_o [3] ), .S(_03071_ ), .Z(_01088_ ) );
MUX2_X1 _19061_ ( .A(\RFU.rf[13][2] ), .B(\EXU.xrd_o [2] ), .S(_03071_ ), .Z(_01089_ ) );
MUX2_X1 _19062_ ( .A(\RFU.rf[13][28] ), .B(\EXU.xrd_o [28] ), .S(_03071_ ), .Z(_01090_ ) );
MUX2_X1 _19063_ ( .A(\RFU.rf[13][1] ), .B(\EXU.xrd_o [1] ), .S(_03071_ ), .Z(_01091_ ) );
MUX2_X1 _19064_ ( .A(\RFU.rf[13][0] ), .B(\EXU.xrd_o [0] ), .S(_03071_ ), .Z(_01092_ ) );
MUX2_X1 _19065_ ( .A(\RFU.rf[13][27] ), .B(\EXU.xrd_o [27] ), .S(_03071_ ), .Z(_01093_ ) );
MUX2_X1 _19066_ ( .A(\RFU.rf[13][26] ), .B(\EXU.xrd_o [26] ), .S(_03071_ ), .Z(_01094_ ) );
MUX2_X1 _19067_ ( .A(\RFU.rf[13][25] ), .B(\EXU.xrd_o [25] ), .S(_03071_ ), .Z(_01095_ ) );
MUX2_X1 _19068_ ( .A(\RFU.rf[13][24] ), .B(\EXU.xrd_o [24] ), .S(_03071_ ), .Z(_01096_ ) );
MUX2_X1 _19069_ ( .A(\RFU.rf[13][23] ), .B(\EXU.xrd_o [23] ), .S(_03068_ ), .Z(_01097_ ) );
MUX2_X1 _19070_ ( .A(\RFU.rf[13][22] ), .B(\EXU.xrd_o [22] ), .S(_03068_ ), .Z(_01098_ ) );
AND4_X1 _19071_ ( .A1(\EXU.rd_o [3] ), .A2(_05434_ ), .A3(\EXU.rd_o [2] ), .A4(\EXU.rd_o [1] ), .ZN(_03072_ ) );
AND2_X2 _19072_ ( .A1(_03051_ ), .A2(_03072_ ), .ZN(_03073_ ) );
BUF_X4 _19073_ ( .A(_03073_ ), .Z(_03074_ ) );
MUX2_X1 _19074_ ( .A(\RFU.rf[14][31] ), .B(\EXU.xrd_o [31] ), .S(_03074_ ), .Z(_01099_ ) );
MUX2_X1 _19075_ ( .A(\RFU.rf[14][30] ), .B(\EXU.xrd_o [30] ), .S(_03074_ ), .Z(_01100_ ) );
MUX2_X1 _19076_ ( .A(\RFU.rf[14][21] ), .B(\EXU.xrd_o [21] ), .S(_03074_ ), .Z(_01101_ ) );
MUX2_X1 _19077_ ( .A(\RFU.rf[14][20] ), .B(\EXU.xrd_o [20] ), .S(_03074_ ), .Z(_01102_ ) );
MUX2_X1 _19078_ ( .A(\RFU.rf[14][19] ), .B(\EXU.xrd_o [19] ), .S(_03074_ ), .Z(_01103_ ) );
MUX2_X1 _19079_ ( .A(\RFU.rf[14][18] ), .B(\EXU.xrd_o [18] ), .S(_03074_ ), .Z(_01104_ ) );
MUX2_X1 _19080_ ( .A(\RFU.rf[14][17] ), .B(\EXU.xrd_o [17] ), .S(_03074_ ), .Z(_01105_ ) );
MUX2_X1 _19081_ ( .A(\RFU.rf[14][16] ), .B(\EXU.xrd_o [16] ), .S(_03074_ ), .Z(_01106_ ) );
MUX2_X1 _19082_ ( .A(\RFU.rf[14][15] ), .B(\EXU.xrd_o [15] ), .S(_03074_ ), .Z(_01107_ ) );
MUX2_X1 _19083_ ( .A(\RFU.rf[14][14] ), .B(\EXU.xrd_o [14] ), .S(_03074_ ), .Z(_01108_ ) );
BUF_X4 _19084_ ( .A(_03073_ ), .Z(_03075_ ) );
MUX2_X1 _19085_ ( .A(\RFU.rf[14][13] ), .B(\EXU.xrd_o [13] ), .S(_03075_ ), .Z(_01109_ ) );
MUX2_X1 _19086_ ( .A(\RFU.rf[14][12] ), .B(\EXU.xrd_o [12] ), .S(_03075_ ), .Z(_01110_ ) );
MUX2_X1 _19087_ ( .A(\RFU.rf[14][29] ), .B(\EXU.xrd_o [29] ), .S(_03075_ ), .Z(_01111_ ) );
MUX2_X1 _19088_ ( .A(\RFU.rf[14][11] ), .B(\EXU.xrd_o [11] ), .S(_03075_ ), .Z(_01112_ ) );
MUX2_X1 _19089_ ( .A(\RFU.rf[14][10] ), .B(\EXU.xrd_o [10] ), .S(_03075_ ), .Z(_01113_ ) );
MUX2_X1 _19090_ ( .A(\RFU.rf[14][9] ), .B(\EXU.xrd_o [9] ), .S(_03075_ ), .Z(_01114_ ) );
MUX2_X1 _19091_ ( .A(\RFU.rf[14][8] ), .B(\EXU.xrd_o [8] ), .S(_03075_ ), .Z(_01115_ ) );
MUX2_X1 _19092_ ( .A(\RFU.rf[14][7] ), .B(\EXU.xrd_o [7] ), .S(_03075_ ), .Z(_01116_ ) );
MUX2_X1 _19093_ ( .A(\RFU.rf[14][6] ), .B(\EXU.xrd_o [6] ), .S(_03075_ ), .Z(_01117_ ) );
MUX2_X1 _19094_ ( .A(\RFU.rf[14][5] ), .B(\EXU.xrd_o [5] ), .S(_03075_ ), .Z(_01118_ ) );
BUF_X4 _19095_ ( .A(_03073_ ), .Z(_03076_ ) );
MUX2_X1 _19096_ ( .A(\RFU.rf[14][4] ), .B(\EXU.xrd_o [4] ), .S(_03076_ ), .Z(_01119_ ) );
MUX2_X1 _19097_ ( .A(\RFU.rf[14][3] ), .B(\EXU.xrd_o [3] ), .S(_03076_ ), .Z(_01120_ ) );
MUX2_X1 _19098_ ( .A(\RFU.rf[14][2] ), .B(\EXU.xrd_o [2] ), .S(_03076_ ), .Z(_01121_ ) );
MUX2_X1 _19099_ ( .A(\RFU.rf[14][28] ), .B(\EXU.xrd_o [28] ), .S(_03076_ ), .Z(_01122_ ) );
MUX2_X1 _19100_ ( .A(\RFU.rf[14][1] ), .B(\EXU.xrd_o [1] ), .S(_03076_ ), .Z(_01123_ ) );
MUX2_X1 _19101_ ( .A(\RFU.rf[14][0] ), .B(\EXU.xrd_o [0] ), .S(_03076_ ), .Z(_01124_ ) );
MUX2_X1 _19102_ ( .A(\RFU.rf[14][27] ), .B(\EXU.xrd_o [27] ), .S(_03076_ ), .Z(_01125_ ) );
MUX2_X1 _19103_ ( .A(\RFU.rf[14][26] ), .B(\EXU.xrd_o [26] ), .S(_03076_ ), .Z(_01126_ ) );
MUX2_X1 _19104_ ( .A(\RFU.rf[14][25] ), .B(\EXU.xrd_o [25] ), .S(_03076_ ), .Z(_01127_ ) );
MUX2_X1 _19105_ ( .A(\RFU.rf[14][24] ), .B(\EXU.xrd_o [24] ), .S(_03076_ ), .Z(_01128_ ) );
MUX2_X1 _19106_ ( .A(\RFU.rf[14][23] ), .B(\EXU.xrd_o [23] ), .S(_03073_ ), .Z(_01129_ ) );
MUX2_X1 _19107_ ( .A(\RFU.rf[14][22] ), .B(\EXU.xrd_o [22] ), .S(_03073_ ), .Z(_01130_ ) );
AND4_X1 _19108_ ( .A1(\EXU.rd_o [3] ), .A2(\EXU.rd_o [2] ), .A3(\EXU.rd_o [1] ), .A4(\EXU.rd_o [0] ), .ZN(_03077_ ) );
AND2_X2 _19109_ ( .A1(_03051_ ), .A2(_03077_ ), .ZN(_03078_ ) );
BUF_X4 _19110_ ( .A(_03078_ ), .Z(_03079_ ) );
MUX2_X1 _19111_ ( .A(\RFU.rf[15][31] ), .B(\EXU.xrd_o [31] ), .S(_03079_ ), .Z(_01131_ ) );
MUX2_X1 _19112_ ( .A(\RFU.rf[15][30] ), .B(\EXU.xrd_o [30] ), .S(_03079_ ), .Z(_01132_ ) );
MUX2_X1 _19113_ ( .A(\RFU.rf[15][21] ), .B(\EXU.xrd_o [21] ), .S(_03079_ ), .Z(_01133_ ) );
MUX2_X1 _19114_ ( .A(\RFU.rf[15][20] ), .B(\EXU.xrd_o [20] ), .S(_03079_ ), .Z(_01134_ ) );
MUX2_X1 _19115_ ( .A(\RFU.rf[15][19] ), .B(\EXU.xrd_o [19] ), .S(_03079_ ), .Z(_01135_ ) );
MUX2_X1 _19116_ ( .A(\RFU.rf[15][18] ), .B(\EXU.xrd_o [18] ), .S(_03079_ ), .Z(_01136_ ) );
MUX2_X1 _19117_ ( .A(\RFU.rf[15][17] ), .B(\EXU.xrd_o [17] ), .S(_03079_ ), .Z(_01137_ ) );
MUX2_X1 _19118_ ( .A(\RFU.rf[15][16] ), .B(\EXU.xrd_o [16] ), .S(_03079_ ), .Z(_01138_ ) );
MUX2_X1 _19119_ ( .A(\RFU.rf[15][15] ), .B(\EXU.xrd_o [15] ), .S(_03079_ ), .Z(_01139_ ) );
MUX2_X1 _19120_ ( .A(\RFU.rf[15][14] ), .B(\EXU.xrd_o [14] ), .S(_03079_ ), .Z(_01140_ ) );
BUF_X4 _19121_ ( .A(_03078_ ), .Z(_03080_ ) );
MUX2_X1 _19122_ ( .A(\RFU.rf[15][13] ), .B(\EXU.xrd_o [13] ), .S(_03080_ ), .Z(_01141_ ) );
MUX2_X1 _19123_ ( .A(\RFU.rf[15][12] ), .B(\EXU.xrd_o [12] ), .S(_03080_ ), .Z(_01142_ ) );
MUX2_X1 _19124_ ( .A(\RFU.rf[15][29] ), .B(\EXU.xrd_o [29] ), .S(_03080_ ), .Z(_01143_ ) );
MUX2_X1 _19125_ ( .A(\RFU.rf[15][11] ), .B(\EXU.xrd_o [11] ), .S(_03080_ ), .Z(_01144_ ) );
MUX2_X1 _19126_ ( .A(\RFU.rf[15][10] ), .B(\EXU.xrd_o [10] ), .S(_03080_ ), .Z(_01145_ ) );
MUX2_X1 _19127_ ( .A(\RFU.rf[15][9] ), .B(\EXU.xrd_o [9] ), .S(_03080_ ), .Z(_01146_ ) );
MUX2_X1 _19128_ ( .A(\RFU.rf[15][8] ), .B(\EXU.xrd_o [8] ), .S(_03080_ ), .Z(_01147_ ) );
MUX2_X1 _19129_ ( .A(\RFU.rf[15][7] ), .B(\EXU.xrd_o [7] ), .S(_03080_ ), .Z(_01148_ ) );
MUX2_X1 _19130_ ( .A(\RFU.rf[15][6] ), .B(\EXU.xrd_o [6] ), .S(_03080_ ), .Z(_01149_ ) );
MUX2_X1 _19131_ ( .A(\RFU.rf[15][5] ), .B(\EXU.xrd_o [5] ), .S(_03080_ ), .Z(_01150_ ) );
BUF_X4 _19132_ ( .A(_03078_ ), .Z(_03081_ ) );
MUX2_X1 _19133_ ( .A(\RFU.rf[15][4] ), .B(\EXU.xrd_o [4] ), .S(_03081_ ), .Z(_01151_ ) );
MUX2_X1 _19134_ ( .A(\RFU.rf[15][3] ), .B(\EXU.xrd_o [3] ), .S(_03081_ ), .Z(_01152_ ) );
MUX2_X1 _19135_ ( .A(\RFU.rf[15][2] ), .B(\EXU.xrd_o [2] ), .S(_03081_ ), .Z(_01153_ ) );
MUX2_X1 _19136_ ( .A(\RFU.rf[15][28] ), .B(\EXU.xrd_o [28] ), .S(_03081_ ), .Z(_01154_ ) );
MUX2_X1 _19137_ ( .A(\RFU.rf[15][1] ), .B(\EXU.xrd_o [1] ), .S(_03081_ ), .Z(_01155_ ) );
MUX2_X1 _19138_ ( .A(\RFU.rf[15][0] ), .B(\EXU.xrd_o [0] ), .S(_03081_ ), .Z(_01156_ ) );
MUX2_X1 _19139_ ( .A(\RFU.rf[15][27] ), .B(\EXU.xrd_o [27] ), .S(_03081_ ), .Z(_01157_ ) );
MUX2_X1 _19140_ ( .A(\RFU.rf[15][26] ), .B(\EXU.xrd_o [26] ), .S(_03081_ ), .Z(_01158_ ) );
MUX2_X1 _19141_ ( .A(\RFU.rf[15][25] ), .B(\EXU.xrd_o [25] ), .S(_03081_ ), .Z(_01159_ ) );
MUX2_X1 _19142_ ( .A(\RFU.rf[15][24] ), .B(\EXU.xrd_o [24] ), .S(_03081_ ), .Z(_01160_ ) );
MUX2_X1 _19143_ ( .A(\RFU.rf[15][23] ), .B(\EXU.xrd_o [23] ), .S(_03078_ ), .Z(_01161_ ) );
MUX2_X1 _19144_ ( .A(\RFU.rf[15][22] ), .B(\EXU.xrd_o [22] ), .S(_03078_ ), .Z(_01162_ ) );
AND4_X1 _19145_ ( .A1(_05428_ ), .A2(_05430_ ), .A3(_05432_ ), .A4(\EXU.rd_o [0] ), .ZN(_03082_ ) );
NAND2_X1 _19146_ ( .A1(_03050_ ), .A2(_03082_ ), .ZN(_03083_ ) );
BUF_X4 _19147_ ( .A(_03083_ ), .Z(_03084_ ) );
MUX2_X1 _19148_ ( .A(\EXU.xrd_o [31] ), .B(\RFU.rf[1][31] ), .S(_03084_ ), .Z(_01163_ ) );
MUX2_X1 _19149_ ( .A(\EXU.xrd_o [30] ), .B(\RFU.rf[1][30] ), .S(_03084_ ), .Z(_01164_ ) );
MUX2_X1 _19150_ ( .A(\EXU.xrd_o [21] ), .B(\RFU.rf[1][21] ), .S(_03084_ ), .Z(_01165_ ) );
MUX2_X1 _19151_ ( .A(\EXU.xrd_o [20] ), .B(\RFU.rf[1][20] ), .S(_03084_ ), .Z(_01166_ ) );
MUX2_X1 _19152_ ( .A(\EXU.xrd_o [19] ), .B(\RFU.rf[1][19] ), .S(_03084_ ), .Z(_01167_ ) );
MUX2_X1 _19153_ ( .A(\EXU.xrd_o [18] ), .B(\RFU.rf[1][18] ), .S(_03084_ ), .Z(_01168_ ) );
MUX2_X1 _19154_ ( .A(\EXU.xrd_o [17] ), .B(\RFU.rf[1][17] ), .S(_03084_ ), .Z(_01169_ ) );
MUX2_X1 _19155_ ( .A(\EXU.xrd_o [16] ), .B(\RFU.rf[1][16] ), .S(_03084_ ), .Z(_01170_ ) );
MUX2_X1 _19156_ ( .A(\EXU.xrd_o [15] ), .B(\RFU.rf[1][15] ), .S(_03084_ ), .Z(_01171_ ) );
MUX2_X1 _19157_ ( .A(\EXU.xrd_o [14] ), .B(\RFU.rf[1][14] ), .S(_03084_ ), .Z(_01172_ ) );
BUF_X4 _19158_ ( .A(_03083_ ), .Z(_03085_ ) );
MUX2_X1 _19159_ ( .A(\EXU.xrd_o [13] ), .B(\RFU.rf[1][13] ), .S(_03085_ ), .Z(_01173_ ) );
MUX2_X1 _19160_ ( .A(\EXU.xrd_o [12] ), .B(\RFU.rf[1][12] ), .S(_03085_ ), .Z(_01174_ ) );
MUX2_X1 _19161_ ( .A(\EXU.xrd_o [29] ), .B(\RFU.rf[1][29] ), .S(_03085_ ), .Z(_01175_ ) );
MUX2_X1 _19162_ ( .A(\EXU.xrd_o [11] ), .B(\RFU.rf[1][11] ), .S(_03085_ ), .Z(_01176_ ) );
MUX2_X1 _19163_ ( .A(\EXU.xrd_o [10] ), .B(\RFU.rf[1][10] ), .S(_03085_ ), .Z(_01177_ ) );
MUX2_X1 _19164_ ( .A(\EXU.xrd_o [9] ), .B(\RFU.rf[1][9] ), .S(_03085_ ), .Z(_01178_ ) );
MUX2_X1 _19165_ ( .A(\EXU.xrd_o [8] ), .B(\RFU.rf[1][8] ), .S(_03085_ ), .Z(_01179_ ) );
MUX2_X1 _19166_ ( .A(\EXU.xrd_o [7] ), .B(\RFU.rf[1][7] ), .S(_03085_ ), .Z(_01180_ ) );
MUX2_X1 _19167_ ( .A(\EXU.xrd_o [6] ), .B(\RFU.rf[1][6] ), .S(_03085_ ), .Z(_01181_ ) );
MUX2_X1 _19168_ ( .A(\EXU.xrd_o [5] ), .B(\RFU.rf[1][5] ), .S(_03085_ ), .Z(_01182_ ) );
BUF_X4 _19169_ ( .A(_03083_ ), .Z(_03086_ ) );
MUX2_X1 _19170_ ( .A(\EXU.xrd_o [4] ), .B(\RFU.rf[1][4] ), .S(_03086_ ), .Z(_01183_ ) );
MUX2_X1 _19171_ ( .A(\EXU.xrd_o [3] ), .B(\RFU.rf[1][3] ), .S(_03086_ ), .Z(_01184_ ) );
MUX2_X1 _19172_ ( .A(\EXU.xrd_o [2] ), .B(\RFU.rf[1][2] ), .S(_03086_ ), .Z(_01185_ ) );
MUX2_X1 _19173_ ( .A(\EXU.xrd_o [28] ), .B(\RFU.rf[1][28] ), .S(_03086_ ), .Z(_01186_ ) );
MUX2_X1 _19174_ ( .A(\EXU.xrd_o [1] ), .B(\RFU.rf[1][1] ), .S(_03086_ ), .Z(_01187_ ) );
MUX2_X1 _19175_ ( .A(\EXU.xrd_o [0] ), .B(\RFU.rf[1][0] ), .S(_03086_ ), .Z(_01188_ ) );
MUX2_X1 _19176_ ( .A(\EXU.xrd_o [27] ), .B(\RFU.rf[1][27] ), .S(_03086_ ), .Z(_01189_ ) );
MUX2_X1 _19177_ ( .A(\EXU.xrd_o [26] ), .B(\RFU.rf[1][26] ), .S(_03086_ ), .Z(_01190_ ) );
MUX2_X1 _19178_ ( .A(\EXU.xrd_o [25] ), .B(\RFU.rf[1][25] ), .S(_03086_ ), .Z(_01191_ ) );
MUX2_X1 _19179_ ( .A(\EXU.xrd_o [24] ), .B(\RFU.rf[1][24] ), .S(_03086_ ), .Z(_01192_ ) );
MUX2_X1 _19180_ ( .A(\EXU.xrd_o [23] ), .B(\RFU.rf[1][23] ), .S(_03083_ ), .Z(_01193_ ) );
MUX2_X1 _19181_ ( .A(\EXU.xrd_o [22] ), .B(\RFU.rf[1][22] ), .S(_03083_ ), .Z(_01194_ ) );
AND4_X1 _19182_ ( .A1(_05428_ ), .A2(_05430_ ), .A3(_05434_ ), .A4(\EXU.rd_o [1] ), .ZN(_03087_ ) );
NAND2_X1 _19183_ ( .A1(_03050_ ), .A2(_03087_ ), .ZN(_03088_ ) );
BUF_X4 _19184_ ( .A(_03088_ ), .Z(_03089_ ) );
MUX2_X1 _19185_ ( .A(\EXU.xrd_o [31] ), .B(\RFU.rf[2][31] ), .S(_03089_ ), .Z(_01195_ ) );
MUX2_X1 _19186_ ( .A(\EXU.xrd_o [30] ), .B(\RFU.rf[2][30] ), .S(_03089_ ), .Z(_01196_ ) );
MUX2_X1 _19187_ ( .A(\EXU.xrd_o [21] ), .B(\RFU.rf[2][21] ), .S(_03089_ ), .Z(_01197_ ) );
MUX2_X1 _19188_ ( .A(\EXU.xrd_o [20] ), .B(\RFU.rf[2][20] ), .S(_03089_ ), .Z(_01198_ ) );
MUX2_X1 _19189_ ( .A(\EXU.xrd_o [19] ), .B(\RFU.rf[2][19] ), .S(_03089_ ), .Z(_01199_ ) );
MUX2_X1 _19190_ ( .A(\EXU.xrd_o [18] ), .B(\RFU.rf[2][18] ), .S(_03089_ ), .Z(_01200_ ) );
MUX2_X1 _19191_ ( .A(\EXU.xrd_o [17] ), .B(\RFU.rf[2][17] ), .S(_03089_ ), .Z(_01201_ ) );
MUX2_X1 _19192_ ( .A(\EXU.xrd_o [16] ), .B(\RFU.rf[2][16] ), .S(_03089_ ), .Z(_01202_ ) );
MUX2_X1 _19193_ ( .A(\EXU.xrd_o [15] ), .B(\RFU.rf[2][15] ), .S(_03089_ ), .Z(_01203_ ) );
MUX2_X1 _19194_ ( .A(\EXU.xrd_o [14] ), .B(\RFU.rf[2][14] ), .S(_03089_ ), .Z(_01204_ ) );
BUF_X4 _19195_ ( .A(_03088_ ), .Z(_03090_ ) );
MUX2_X1 _19196_ ( .A(\EXU.xrd_o [13] ), .B(\RFU.rf[2][13] ), .S(_03090_ ), .Z(_01205_ ) );
MUX2_X1 _19197_ ( .A(\EXU.xrd_o [12] ), .B(\RFU.rf[2][12] ), .S(_03090_ ), .Z(_01206_ ) );
MUX2_X1 _19198_ ( .A(\EXU.xrd_o [29] ), .B(\RFU.rf[2][29] ), .S(_03090_ ), .Z(_01207_ ) );
MUX2_X1 _19199_ ( .A(\EXU.xrd_o [11] ), .B(\RFU.rf[2][11] ), .S(_03090_ ), .Z(_01208_ ) );
MUX2_X1 _19200_ ( .A(\EXU.xrd_o [10] ), .B(\RFU.rf[2][10] ), .S(_03090_ ), .Z(_01209_ ) );
MUX2_X1 _19201_ ( .A(\EXU.xrd_o [9] ), .B(\RFU.rf[2][9] ), .S(_03090_ ), .Z(_01210_ ) );
MUX2_X1 _19202_ ( .A(\EXU.xrd_o [8] ), .B(\RFU.rf[2][8] ), .S(_03090_ ), .Z(_01211_ ) );
MUX2_X1 _19203_ ( .A(\EXU.xrd_o [7] ), .B(\RFU.rf[2][7] ), .S(_03090_ ), .Z(_01212_ ) );
MUX2_X1 _19204_ ( .A(\EXU.xrd_o [6] ), .B(\RFU.rf[2][6] ), .S(_03090_ ), .Z(_01213_ ) );
MUX2_X1 _19205_ ( .A(\EXU.xrd_o [5] ), .B(\RFU.rf[2][5] ), .S(_03090_ ), .Z(_01214_ ) );
BUF_X4 _19206_ ( .A(_03088_ ), .Z(_03091_ ) );
MUX2_X1 _19207_ ( .A(\EXU.xrd_o [4] ), .B(\RFU.rf[2][4] ), .S(_03091_ ), .Z(_01215_ ) );
MUX2_X1 _19208_ ( .A(\EXU.xrd_o [3] ), .B(\RFU.rf[2][3] ), .S(_03091_ ), .Z(_01216_ ) );
MUX2_X1 _19209_ ( .A(\EXU.xrd_o [2] ), .B(\RFU.rf[2][2] ), .S(_03091_ ), .Z(_01217_ ) );
MUX2_X1 _19210_ ( .A(\EXU.xrd_o [28] ), .B(\RFU.rf[2][28] ), .S(_03091_ ), .Z(_01218_ ) );
MUX2_X1 _19211_ ( .A(\EXU.xrd_o [1] ), .B(\RFU.rf[2][1] ), .S(_03091_ ), .Z(_01219_ ) );
MUX2_X1 _19212_ ( .A(\EXU.xrd_o [0] ), .B(\RFU.rf[2][0] ), .S(_03091_ ), .Z(_01220_ ) );
MUX2_X1 _19213_ ( .A(\EXU.xrd_o [27] ), .B(\RFU.rf[2][27] ), .S(_03091_ ), .Z(_01221_ ) );
MUX2_X1 _19214_ ( .A(\EXU.xrd_o [26] ), .B(\RFU.rf[2][26] ), .S(_03091_ ), .Z(_01222_ ) );
MUX2_X1 _19215_ ( .A(\EXU.xrd_o [25] ), .B(\RFU.rf[2][25] ), .S(_03091_ ), .Z(_01223_ ) );
MUX2_X1 _19216_ ( .A(\EXU.xrd_o [24] ), .B(\RFU.rf[2][24] ), .S(_03091_ ), .Z(_01224_ ) );
MUX2_X1 _19217_ ( .A(\EXU.xrd_o [23] ), .B(\RFU.rf[2][23] ), .S(_03088_ ), .Z(_01225_ ) );
MUX2_X1 _19218_ ( .A(\EXU.xrd_o [22] ), .B(\RFU.rf[2][22] ), .S(_03088_ ), .Z(_01226_ ) );
AND4_X1 _19219_ ( .A1(_05428_ ), .A2(_05430_ ), .A3(\EXU.rd_o [1] ), .A4(\EXU.rd_o [0] ), .ZN(_03092_ ) );
NAND2_X1 _19220_ ( .A1(_03050_ ), .A2(_03092_ ), .ZN(_03093_ ) );
BUF_X4 _19221_ ( .A(_03093_ ), .Z(_03094_ ) );
MUX2_X1 _19222_ ( .A(\EXU.xrd_o [31] ), .B(\RFU.rf[3][31] ), .S(_03094_ ), .Z(_01227_ ) );
MUX2_X1 _19223_ ( .A(\EXU.xrd_o [30] ), .B(\RFU.rf[3][30] ), .S(_03094_ ), .Z(_01228_ ) );
MUX2_X1 _19224_ ( .A(\EXU.xrd_o [21] ), .B(\RFU.rf[3][21] ), .S(_03094_ ), .Z(_01229_ ) );
MUX2_X1 _19225_ ( .A(\EXU.xrd_o [20] ), .B(\RFU.rf[3][20] ), .S(_03094_ ), .Z(_01230_ ) );
MUX2_X1 _19226_ ( .A(\EXU.xrd_o [19] ), .B(\RFU.rf[3][19] ), .S(_03094_ ), .Z(_01231_ ) );
MUX2_X1 _19227_ ( .A(\EXU.xrd_o [18] ), .B(\RFU.rf[3][18] ), .S(_03094_ ), .Z(_01232_ ) );
MUX2_X1 _19228_ ( .A(\EXU.xrd_o [17] ), .B(\RFU.rf[3][17] ), .S(_03094_ ), .Z(_01233_ ) );
MUX2_X1 _19229_ ( .A(\EXU.xrd_o [16] ), .B(\RFU.rf[3][16] ), .S(_03094_ ), .Z(_01234_ ) );
MUX2_X1 _19230_ ( .A(\EXU.xrd_o [15] ), .B(\RFU.rf[3][15] ), .S(_03094_ ), .Z(_01235_ ) );
MUX2_X1 _19231_ ( .A(\EXU.xrd_o [14] ), .B(\RFU.rf[3][14] ), .S(_03094_ ), .Z(_01236_ ) );
BUF_X4 _19232_ ( .A(_03093_ ), .Z(_03095_ ) );
MUX2_X1 _19233_ ( .A(\EXU.xrd_o [13] ), .B(\RFU.rf[3][13] ), .S(_03095_ ), .Z(_01237_ ) );
MUX2_X1 _19234_ ( .A(\EXU.xrd_o [12] ), .B(\RFU.rf[3][12] ), .S(_03095_ ), .Z(_01238_ ) );
MUX2_X1 _19235_ ( .A(\EXU.xrd_o [29] ), .B(\RFU.rf[3][29] ), .S(_03095_ ), .Z(_01239_ ) );
MUX2_X1 _19236_ ( .A(\EXU.xrd_o [11] ), .B(\RFU.rf[3][11] ), .S(_03095_ ), .Z(_01240_ ) );
MUX2_X1 _19237_ ( .A(\EXU.xrd_o [10] ), .B(\RFU.rf[3][10] ), .S(_03095_ ), .Z(_01241_ ) );
MUX2_X1 _19238_ ( .A(\EXU.xrd_o [9] ), .B(\RFU.rf[3][9] ), .S(_03095_ ), .Z(_01242_ ) );
MUX2_X1 _19239_ ( .A(\EXU.xrd_o [8] ), .B(\RFU.rf[3][8] ), .S(_03095_ ), .Z(_01243_ ) );
MUX2_X1 _19240_ ( .A(\EXU.xrd_o [7] ), .B(\RFU.rf[3][7] ), .S(_03095_ ), .Z(_01244_ ) );
MUX2_X1 _19241_ ( .A(\EXU.xrd_o [6] ), .B(\RFU.rf[3][6] ), .S(_03095_ ), .Z(_01245_ ) );
MUX2_X1 _19242_ ( .A(\EXU.xrd_o [5] ), .B(\RFU.rf[3][5] ), .S(_03095_ ), .Z(_01246_ ) );
BUF_X4 _19243_ ( .A(_03093_ ), .Z(_03096_ ) );
MUX2_X1 _19244_ ( .A(\EXU.xrd_o [4] ), .B(\RFU.rf[3][4] ), .S(_03096_ ), .Z(_01247_ ) );
MUX2_X1 _19245_ ( .A(\EXU.xrd_o [3] ), .B(\RFU.rf[3][3] ), .S(_03096_ ), .Z(_01248_ ) );
MUX2_X1 _19246_ ( .A(\EXU.xrd_o [2] ), .B(\RFU.rf[3][2] ), .S(_03096_ ), .Z(_01249_ ) );
MUX2_X1 _19247_ ( .A(\EXU.xrd_o [28] ), .B(\RFU.rf[3][28] ), .S(_03096_ ), .Z(_01250_ ) );
MUX2_X1 _19248_ ( .A(\EXU.xrd_o [1] ), .B(\RFU.rf[3][1] ), .S(_03096_ ), .Z(_01251_ ) );
MUX2_X1 _19249_ ( .A(\EXU.xrd_o [0] ), .B(\RFU.rf[3][0] ), .S(_03096_ ), .Z(_01252_ ) );
MUX2_X1 _19250_ ( .A(\EXU.xrd_o [27] ), .B(\RFU.rf[3][27] ), .S(_03096_ ), .Z(_01253_ ) );
MUX2_X1 _19251_ ( .A(\EXU.xrd_o [26] ), .B(\RFU.rf[3][26] ), .S(_03096_ ), .Z(_01254_ ) );
MUX2_X1 _19252_ ( .A(\EXU.xrd_o [25] ), .B(\RFU.rf[3][25] ), .S(_03096_ ), .Z(_01255_ ) );
MUX2_X1 _19253_ ( .A(\EXU.xrd_o [24] ), .B(\RFU.rf[3][24] ), .S(_03096_ ), .Z(_01256_ ) );
MUX2_X1 _19254_ ( .A(\EXU.xrd_o [23] ), .B(\RFU.rf[3][23] ), .S(_03093_ ), .Z(_01257_ ) );
MUX2_X1 _19255_ ( .A(\EXU.xrd_o [22] ), .B(\RFU.rf[3][22] ), .S(_03093_ ), .Z(_01258_ ) );
AND4_X1 _19256_ ( .A1(_05428_ ), .A2(_05432_ ), .A3(_05434_ ), .A4(\EXU.rd_o [2] ), .ZN(_03097_ ) );
NAND2_X1 _19257_ ( .A1(_03050_ ), .A2(_03097_ ), .ZN(_03098_ ) );
BUF_X4 _19258_ ( .A(_03098_ ), .Z(_03099_ ) );
MUX2_X1 _19259_ ( .A(\EXU.xrd_o [31] ), .B(\RFU.rf[4][31] ), .S(_03099_ ), .Z(_01259_ ) );
MUX2_X1 _19260_ ( .A(\EXU.xrd_o [30] ), .B(\RFU.rf[4][30] ), .S(_03099_ ), .Z(_01260_ ) );
MUX2_X1 _19261_ ( .A(\EXU.xrd_o [21] ), .B(\RFU.rf[4][21] ), .S(_03099_ ), .Z(_01261_ ) );
MUX2_X1 _19262_ ( .A(\EXU.xrd_o [20] ), .B(\RFU.rf[4][20] ), .S(_03099_ ), .Z(_01262_ ) );
MUX2_X1 _19263_ ( .A(\EXU.xrd_o [19] ), .B(\RFU.rf[4][19] ), .S(_03099_ ), .Z(_01263_ ) );
MUX2_X1 _19264_ ( .A(\EXU.xrd_o [18] ), .B(\RFU.rf[4][18] ), .S(_03099_ ), .Z(_01264_ ) );
MUX2_X1 _19265_ ( .A(\EXU.xrd_o [17] ), .B(\RFU.rf[4][17] ), .S(_03099_ ), .Z(_01265_ ) );
MUX2_X1 _19266_ ( .A(\EXU.xrd_o [16] ), .B(\RFU.rf[4][16] ), .S(_03099_ ), .Z(_01266_ ) );
MUX2_X1 _19267_ ( .A(\EXU.xrd_o [15] ), .B(\RFU.rf[4][15] ), .S(_03099_ ), .Z(_01267_ ) );
MUX2_X1 _19268_ ( .A(\EXU.xrd_o [14] ), .B(\RFU.rf[4][14] ), .S(_03099_ ), .Z(_01268_ ) );
BUF_X4 _19269_ ( .A(_03098_ ), .Z(_03100_ ) );
MUX2_X1 _19270_ ( .A(\EXU.xrd_o [13] ), .B(\RFU.rf[4][13] ), .S(_03100_ ), .Z(_01269_ ) );
MUX2_X1 _19271_ ( .A(\EXU.xrd_o [12] ), .B(\RFU.rf[4][12] ), .S(_03100_ ), .Z(_01270_ ) );
MUX2_X1 _19272_ ( .A(\EXU.xrd_o [29] ), .B(\RFU.rf[4][29] ), .S(_03100_ ), .Z(_01271_ ) );
MUX2_X1 _19273_ ( .A(\EXU.xrd_o [11] ), .B(\RFU.rf[4][11] ), .S(_03100_ ), .Z(_01272_ ) );
MUX2_X1 _19274_ ( .A(\EXU.xrd_o [10] ), .B(\RFU.rf[4][10] ), .S(_03100_ ), .Z(_01273_ ) );
MUX2_X1 _19275_ ( .A(\EXU.xrd_o [9] ), .B(\RFU.rf[4][9] ), .S(_03100_ ), .Z(_01274_ ) );
MUX2_X1 _19276_ ( .A(\EXU.xrd_o [8] ), .B(\RFU.rf[4][8] ), .S(_03100_ ), .Z(_01275_ ) );
MUX2_X1 _19277_ ( .A(\EXU.xrd_o [7] ), .B(\RFU.rf[4][7] ), .S(_03100_ ), .Z(_01276_ ) );
MUX2_X1 _19278_ ( .A(\EXU.xrd_o [6] ), .B(\RFU.rf[4][6] ), .S(_03100_ ), .Z(_01277_ ) );
MUX2_X1 _19279_ ( .A(\EXU.xrd_o [5] ), .B(\RFU.rf[4][5] ), .S(_03100_ ), .Z(_01278_ ) );
BUF_X4 _19280_ ( .A(_03098_ ), .Z(_03101_ ) );
MUX2_X1 _19281_ ( .A(\EXU.xrd_o [4] ), .B(\RFU.rf[4][4] ), .S(_03101_ ), .Z(_01279_ ) );
MUX2_X1 _19282_ ( .A(\EXU.xrd_o [3] ), .B(\RFU.rf[4][3] ), .S(_03101_ ), .Z(_01280_ ) );
MUX2_X1 _19283_ ( .A(\EXU.xrd_o [2] ), .B(\RFU.rf[4][2] ), .S(_03101_ ), .Z(_01281_ ) );
MUX2_X1 _19284_ ( .A(\EXU.xrd_o [28] ), .B(\RFU.rf[4][28] ), .S(_03101_ ), .Z(_01282_ ) );
MUX2_X1 _19285_ ( .A(\EXU.xrd_o [1] ), .B(\RFU.rf[4][1] ), .S(_03101_ ), .Z(_01283_ ) );
MUX2_X1 _19286_ ( .A(\EXU.xrd_o [0] ), .B(\RFU.rf[4][0] ), .S(_03101_ ), .Z(_01284_ ) );
MUX2_X1 _19287_ ( .A(\EXU.xrd_o [27] ), .B(\RFU.rf[4][27] ), .S(_03101_ ), .Z(_01285_ ) );
MUX2_X1 _19288_ ( .A(\EXU.xrd_o [26] ), .B(\RFU.rf[4][26] ), .S(_03101_ ), .Z(_01286_ ) );
MUX2_X1 _19289_ ( .A(\EXU.xrd_o [25] ), .B(\RFU.rf[4][25] ), .S(_03101_ ), .Z(_01287_ ) );
MUX2_X1 _19290_ ( .A(\EXU.xrd_o [24] ), .B(\RFU.rf[4][24] ), .S(_03101_ ), .Z(_01288_ ) );
MUX2_X1 _19291_ ( .A(\EXU.xrd_o [23] ), .B(\RFU.rf[4][23] ), .S(_03098_ ), .Z(_01289_ ) );
MUX2_X1 _19292_ ( .A(\EXU.xrd_o [22] ), .B(\RFU.rf[4][22] ), .S(_03098_ ), .Z(_01290_ ) );
AND4_X1 _19293_ ( .A1(_05428_ ), .A2(_05432_ ), .A3(\EXU.rd_o [2] ), .A4(\EXU.rd_o [0] ), .ZN(_03102_ ) );
AND2_X2 _19294_ ( .A1(_03051_ ), .A2(_03102_ ), .ZN(_03103_ ) );
BUF_X4 _19295_ ( .A(_03103_ ), .Z(_03104_ ) );
MUX2_X1 _19296_ ( .A(\RFU.rf[5][31] ), .B(\EXU.xrd_o [31] ), .S(_03104_ ), .Z(_01291_ ) );
MUX2_X1 _19297_ ( .A(\RFU.rf[5][30] ), .B(\EXU.xrd_o [30] ), .S(_03104_ ), .Z(_01292_ ) );
MUX2_X1 _19298_ ( .A(\RFU.rf[5][21] ), .B(\EXU.xrd_o [21] ), .S(_03104_ ), .Z(_01293_ ) );
MUX2_X1 _19299_ ( .A(\RFU.rf[5][20] ), .B(\EXU.xrd_o [20] ), .S(_03104_ ), .Z(_01294_ ) );
MUX2_X1 _19300_ ( .A(\RFU.rf[5][19] ), .B(\EXU.xrd_o [19] ), .S(_03104_ ), .Z(_01295_ ) );
MUX2_X1 _19301_ ( .A(\RFU.rf[5][18] ), .B(\EXU.xrd_o [18] ), .S(_03104_ ), .Z(_01296_ ) );
MUX2_X1 _19302_ ( .A(\RFU.rf[5][17] ), .B(\EXU.xrd_o [17] ), .S(_03104_ ), .Z(_01297_ ) );
MUX2_X1 _19303_ ( .A(\RFU.rf[5][16] ), .B(\EXU.xrd_o [16] ), .S(_03104_ ), .Z(_01298_ ) );
MUX2_X1 _19304_ ( .A(\RFU.rf[5][15] ), .B(\EXU.xrd_o [15] ), .S(_03104_ ), .Z(_01299_ ) );
MUX2_X1 _19305_ ( .A(\RFU.rf[5][14] ), .B(\EXU.xrd_o [14] ), .S(_03104_ ), .Z(_01300_ ) );
BUF_X4 _19306_ ( .A(_03103_ ), .Z(_03105_ ) );
MUX2_X1 _19307_ ( .A(\RFU.rf[5][13] ), .B(\EXU.xrd_o [13] ), .S(_03105_ ), .Z(_01301_ ) );
MUX2_X1 _19308_ ( .A(\RFU.rf[5][12] ), .B(\EXU.xrd_o [12] ), .S(_03105_ ), .Z(_01302_ ) );
MUX2_X1 _19309_ ( .A(\RFU.rf[5][29] ), .B(\EXU.xrd_o [29] ), .S(_03105_ ), .Z(_01303_ ) );
MUX2_X1 _19310_ ( .A(\RFU.rf[5][11] ), .B(\EXU.xrd_o [11] ), .S(_03105_ ), .Z(_01304_ ) );
MUX2_X1 _19311_ ( .A(\RFU.rf[5][10] ), .B(\EXU.xrd_o [10] ), .S(_03105_ ), .Z(_01305_ ) );
MUX2_X1 _19312_ ( .A(\RFU.rf[5][9] ), .B(\EXU.xrd_o [9] ), .S(_03105_ ), .Z(_01306_ ) );
MUX2_X1 _19313_ ( .A(\RFU.rf[5][8] ), .B(\EXU.xrd_o [8] ), .S(_03105_ ), .Z(_01307_ ) );
MUX2_X1 _19314_ ( .A(\RFU.rf[5][7] ), .B(\EXU.xrd_o [7] ), .S(_03105_ ), .Z(_01308_ ) );
MUX2_X1 _19315_ ( .A(\RFU.rf[5][6] ), .B(\EXU.xrd_o [6] ), .S(_03105_ ), .Z(_01309_ ) );
MUX2_X1 _19316_ ( .A(\RFU.rf[5][5] ), .B(\EXU.xrd_o [5] ), .S(_03105_ ), .Z(_01310_ ) );
BUF_X4 _19317_ ( .A(_03103_ ), .Z(_03106_ ) );
MUX2_X1 _19318_ ( .A(\RFU.rf[5][4] ), .B(\EXU.xrd_o [4] ), .S(_03106_ ), .Z(_01311_ ) );
MUX2_X1 _19319_ ( .A(\RFU.rf[5][3] ), .B(\EXU.xrd_o [3] ), .S(_03106_ ), .Z(_01312_ ) );
MUX2_X1 _19320_ ( .A(\RFU.rf[5][2] ), .B(\EXU.xrd_o [2] ), .S(_03106_ ), .Z(_01313_ ) );
MUX2_X1 _19321_ ( .A(\RFU.rf[5][28] ), .B(\EXU.xrd_o [28] ), .S(_03106_ ), .Z(_01314_ ) );
MUX2_X1 _19322_ ( .A(\RFU.rf[5][1] ), .B(\EXU.xrd_o [1] ), .S(_03106_ ), .Z(_01315_ ) );
MUX2_X1 _19323_ ( .A(\RFU.rf[5][0] ), .B(\EXU.xrd_o [0] ), .S(_03106_ ), .Z(_01316_ ) );
MUX2_X1 _19324_ ( .A(\RFU.rf[5][27] ), .B(\EXU.xrd_o [27] ), .S(_03106_ ), .Z(_01317_ ) );
MUX2_X1 _19325_ ( .A(\RFU.rf[5][26] ), .B(\EXU.xrd_o [26] ), .S(_03106_ ), .Z(_01318_ ) );
MUX2_X1 _19326_ ( .A(\RFU.rf[5][25] ), .B(\EXU.xrd_o [25] ), .S(_03106_ ), .Z(_01319_ ) );
MUX2_X1 _19327_ ( .A(\RFU.rf[5][24] ), .B(\EXU.xrd_o [24] ), .S(_03106_ ), .Z(_01320_ ) );
MUX2_X1 _19328_ ( .A(\RFU.rf[5][23] ), .B(\EXU.xrd_o [23] ), .S(_03103_ ), .Z(_01321_ ) );
MUX2_X1 _19329_ ( .A(\RFU.rf[5][22] ), .B(\EXU.xrd_o [22] ), .S(_03103_ ), .Z(_01322_ ) );
AND4_X1 _19330_ ( .A1(_05428_ ), .A2(_05434_ ), .A3(\EXU.rd_o [2] ), .A4(\EXU.rd_o [1] ), .ZN(_03107_ ) );
AND2_X2 _19331_ ( .A1(_03051_ ), .A2(_03107_ ), .ZN(_03108_ ) );
BUF_X4 _19332_ ( .A(_03108_ ), .Z(_03109_ ) );
MUX2_X1 _19333_ ( .A(\RFU.rf[6][31] ), .B(\EXU.xrd_o [31] ), .S(_03109_ ), .Z(_01323_ ) );
MUX2_X1 _19334_ ( .A(\RFU.rf[6][30] ), .B(\EXU.xrd_o [30] ), .S(_03109_ ), .Z(_01324_ ) );
MUX2_X1 _19335_ ( .A(\RFU.rf[6][21] ), .B(\EXU.xrd_o [21] ), .S(_03109_ ), .Z(_01325_ ) );
MUX2_X1 _19336_ ( .A(\RFU.rf[6][20] ), .B(\EXU.xrd_o [20] ), .S(_03109_ ), .Z(_01326_ ) );
MUX2_X1 _19337_ ( .A(\RFU.rf[6][19] ), .B(\EXU.xrd_o [19] ), .S(_03109_ ), .Z(_01327_ ) );
MUX2_X1 _19338_ ( .A(\RFU.rf[6][18] ), .B(\EXU.xrd_o [18] ), .S(_03109_ ), .Z(_01328_ ) );
MUX2_X1 _19339_ ( .A(\RFU.rf[6][17] ), .B(\EXU.xrd_o [17] ), .S(_03109_ ), .Z(_01329_ ) );
MUX2_X1 _19340_ ( .A(\RFU.rf[6][16] ), .B(\EXU.xrd_o [16] ), .S(_03109_ ), .Z(_01330_ ) );
MUX2_X1 _19341_ ( .A(\RFU.rf[6][15] ), .B(\EXU.xrd_o [15] ), .S(_03109_ ), .Z(_01331_ ) );
MUX2_X1 _19342_ ( .A(\RFU.rf[6][14] ), .B(\EXU.xrd_o [14] ), .S(_03109_ ), .Z(_01332_ ) );
BUF_X4 _19343_ ( .A(_03108_ ), .Z(_03110_ ) );
MUX2_X1 _19344_ ( .A(\RFU.rf[6][13] ), .B(\EXU.xrd_o [13] ), .S(_03110_ ), .Z(_01333_ ) );
MUX2_X1 _19345_ ( .A(\RFU.rf[6][12] ), .B(\EXU.xrd_o [12] ), .S(_03110_ ), .Z(_01334_ ) );
MUX2_X1 _19346_ ( .A(\RFU.rf[6][29] ), .B(\EXU.xrd_o [29] ), .S(_03110_ ), .Z(_01335_ ) );
MUX2_X1 _19347_ ( .A(\RFU.rf[6][11] ), .B(\EXU.xrd_o [11] ), .S(_03110_ ), .Z(_01336_ ) );
MUX2_X1 _19348_ ( .A(\RFU.rf[6][10] ), .B(\EXU.xrd_o [10] ), .S(_03110_ ), .Z(_01337_ ) );
MUX2_X1 _19349_ ( .A(\RFU.rf[6][9] ), .B(\EXU.xrd_o [9] ), .S(_03110_ ), .Z(_01338_ ) );
MUX2_X1 _19350_ ( .A(\RFU.rf[6][8] ), .B(\EXU.xrd_o [8] ), .S(_03110_ ), .Z(_01339_ ) );
MUX2_X1 _19351_ ( .A(\RFU.rf[6][7] ), .B(\EXU.xrd_o [7] ), .S(_03110_ ), .Z(_01340_ ) );
MUX2_X1 _19352_ ( .A(\RFU.rf[6][6] ), .B(\EXU.xrd_o [6] ), .S(_03110_ ), .Z(_01341_ ) );
MUX2_X1 _19353_ ( .A(\RFU.rf[6][5] ), .B(\EXU.xrd_o [5] ), .S(_03110_ ), .Z(_01342_ ) );
BUF_X4 _19354_ ( .A(_03108_ ), .Z(_03111_ ) );
MUX2_X1 _19355_ ( .A(\RFU.rf[6][4] ), .B(\EXU.xrd_o [4] ), .S(_03111_ ), .Z(_01343_ ) );
MUX2_X1 _19356_ ( .A(\RFU.rf[6][3] ), .B(\EXU.xrd_o [3] ), .S(_03111_ ), .Z(_01344_ ) );
MUX2_X1 _19357_ ( .A(\RFU.rf[6][2] ), .B(\EXU.xrd_o [2] ), .S(_03111_ ), .Z(_01345_ ) );
MUX2_X1 _19358_ ( .A(\RFU.rf[6][28] ), .B(\EXU.xrd_o [28] ), .S(_03111_ ), .Z(_01346_ ) );
MUX2_X1 _19359_ ( .A(\RFU.rf[6][1] ), .B(\EXU.xrd_o [1] ), .S(_03111_ ), .Z(_01347_ ) );
MUX2_X1 _19360_ ( .A(\RFU.rf[6][0] ), .B(\EXU.xrd_o [0] ), .S(_03111_ ), .Z(_01348_ ) );
MUX2_X1 _19361_ ( .A(\RFU.rf[6][27] ), .B(\EXU.xrd_o [27] ), .S(_03111_ ), .Z(_01349_ ) );
MUX2_X1 _19362_ ( .A(\RFU.rf[6][26] ), .B(\EXU.xrd_o [26] ), .S(_03111_ ), .Z(_01350_ ) );
MUX2_X1 _19363_ ( .A(\RFU.rf[6][25] ), .B(\EXU.xrd_o [25] ), .S(_03111_ ), .Z(_01351_ ) );
MUX2_X1 _19364_ ( .A(\RFU.rf[6][24] ), .B(\EXU.xrd_o [24] ), .S(_03111_ ), .Z(_01352_ ) );
MUX2_X1 _19365_ ( .A(\RFU.rf[6][23] ), .B(\EXU.xrd_o [23] ), .S(_03108_ ), .Z(_01353_ ) );
MUX2_X1 _19366_ ( .A(\RFU.rf[6][22] ), .B(\EXU.xrd_o [22] ), .S(_03108_ ), .Z(_01354_ ) );
AND4_X1 _19367_ ( .A1(_05428_ ), .A2(\EXU.rd_o [2] ), .A3(\EXU.rd_o [1] ), .A4(\EXU.rd_o [0] ), .ZN(_03112_ ) );
AND2_X2 _19368_ ( .A1(_03051_ ), .A2(_03112_ ), .ZN(_03113_ ) );
BUF_X4 _19369_ ( .A(_03113_ ), .Z(_03114_ ) );
MUX2_X1 _19370_ ( .A(\RFU.rf[7][31] ), .B(\EXU.xrd_o [31] ), .S(_03114_ ), .Z(_01355_ ) );
MUX2_X1 _19371_ ( .A(\RFU.rf[7][30] ), .B(\EXU.xrd_o [30] ), .S(_03114_ ), .Z(_01356_ ) );
MUX2_X1 _19372_ ( .A(\RFU.rf[7][21] ), .B(\EXU.xrd_o [21] ), .S(_03114_ ), .Z(_01357_ ) );
MUX2_X1 _19373_ ( .A(\RFU.rf[7][20] ), .B(\EXU.xrd_o [20] ), .S(_03114_ ), .Z(_01358_ ) );
MUX2_X1 _19374_ ( .A(\RFU.rf[7][19] ), .B(\EXU.xrd_o [19] ), .S(_03114_ ), .Z(_01359_ ) );
MUX2_X1 _19375_ ( .A(\RFU.rf[7][18] ), .B(\EXU.xrd_o [18] ), .S(_03114_ ), .Z(_01360_ ) );
MUX2_X1 _19376_ ( .A(\RFU.rf[7][17] ), .B(\EXU.xrd_o [17] ), .S(_03114_ ), .Z(_01361_ ) );
MUX2_X1 _19377_ ( .A(\RFU.rf[7][16] ), .B(\EXU.xrd_o [16] ), .S(_03114_ ), .Z(_01362_ ) );
MUX2_X1 _19378_ ( .A(\RFU.rf[7][15] ), .B(\EXU.xrd_o [15] ), .S(_03114_ ), .Z(_01363_ ) );
MUX2_X1 _19379_ ( .A(\RFU.rf[7][14] ), .B(\EXU.xrd_o [14] ), .S(_03114_ ), .Z(_01364_ ) );
BUF_X4 _19380_ ( .A(_03113_ ), .Z(_03115_ ) );
MUX2_X1 _19381_ ( .A(\RFU.rf[7][13] ), .B(\EXU.xrd_o [13] ), .S(_03115_ ), .Z(_01365_ ) );
MUX2_X1 _19382_ ( .A(\RFU.rf[7][12] ), .B(\EXU.xrd_o [12] ), .S(_03115_ ), .Z(_01366_ ) );
MUX2_X1 _19383_ ( .A(\RFU.rf[7][29] ), .B(\EXU.xrd_o [29] ), .S(_03115_ ), .Z(_01367_ ) );
MUX2_X1 _19384_ ( .A(\RFU.rf[7][11] ), .B(\EXU.xrd_o [11] ), .S(_03115_ ), .Z(_01368_ ) );
MUX2_X1 _19385_ ( .A(\RFU.rf[7][10] ), .B(\EXU.xrd_o [10] ), .S(_03115_ ), .Z(_01369_ ) );
MUX2_X1 _19386_ ( .A(\RFU.rf[7][9] ), .B(\EXU.xrd_o [9] ), .S(_03115_ ), .Z(_01370_ ) );
MUX2_X1 _19387_ ( .A(\RFU.rf[7][8] ), .B(\EXU.xrd_o [8] ), .S(_03115_ ), .Z(_01371_ ) );
MUX2_X1 _19388_ ( .A(\RFU.rf[7][7] ), .B(\EXU.xrd_o [7] ), .S(_03115_ ), .Z(_01372_ ) );
MUX2_X1 _19389_ ( .A(\RFU.rf[7][6] ), .B(\EXU.xrd_o [6] ), .S(_03115_ ), .Z(_01373_ ) );
MUX2_X1 _19390_ ( .A(\RFU.rf[7][5] ), .B(\EXU.xrd_o [5] ), .S(_03115_ ), .Z(_01374_ ) );
BUF_X4 _19391_ ( .A(_03113_ ), .Z(_03116_ ) );
MUX2_X1 _19392_ ( .A(\RFU.rf[7][4] ), .B(\EXU.xrd_o [4] ), .S(_03116_ ), .Z(_01375_ ) );
MUX2_X1 _19393_ ( .A(\RFU.rf[7][3] ), .B(\EXU.xrd_o [3] ), .S(_03116_ ), .Z(_01376_ ) );
MUX2_X1 _19394_ ( .A(\RFU.rf[7][2] ), .B(\EXU.xrd_o [2] ), .S(_03116_ ), .Z(_01377_ ) );
MUX2_X1 _19395_ ( .A(\RFU.rf[7][28] ), .B(\EXU.xrd_o [28] ), .S(_03116_ ), .Z(_01378_ ) );
MUX2_X1 _19396_ ( .A(\RFU.rf[7][1] ), .B(\EXU.xrd_o [1] ), .S(_03116_ ), .Z(_01379_ ) );
MUX2_X1 _19397_ ( .A(\RFU.rf[7][0] ), .B(\EXU.xrd_o [0] ), .S(_03116_ ), .Z(_01380_ ) );
MUX2_X1 _19398_ ( .A(\RFU.rf[7][27] ), .B(\EXU.xrd_o [27] ), .S(_03116_ ), .Z(_01381_ ) );
MUX2_X1 _19399_ ( .A(\RFU.rf[7][26] ), .B(\EXU.xrd_o [26] ), .S(_03116_ ), .Z(_01382_ ) );
MUX2_X1 _19400_ ( .A(\RFU.rf[7][25] ), .B(\EXU.xrd_o [25] ), .S(_03116_ ), .Z(_01383_ ) );
MUX2_X1 _19401_ ( .A(\RFU.rf[7][24] ), .B(\EXU.xrd_o [24] ), .S(_03116_ ), .Z(_01384_ ) );
MUX2_X1 _19402_ ( .A(\RFU.rf[7][23] ), .B(\EXU.xrd_o [23] ), .S(_03113_ ), .Z(_01385_ ) );
MUX2_X1 _19403_ ( .A(\RFU.rf[7][22] ), .B(\EXU.xrd_o [22] ), .S(_03113_ ), .Z(_01386_ ) );
NOR4_X1 _19404_ ( .A1(_05428_ ), .A2(\EXU.rd_o [2] ), .A3(\EXU.rd_o [1] ), .A4(\EXU.rd_o [0] ), .ZN(_03117_ ) );
NAND2_X1 _19405_ ( .A1(_03050_ ), .A2(_03117_ ), .ZN(_03118_ ) );
BUF_X4 _19406_ ( .A(_03118_ ), .Z(_03119_ ) );
MUX2_X1 _19407_ ( .A(\EXU.xrd_o [31] ), .B(\RFU.rf[8][31] ), .S(_03119_ ), .Z(_01387_ ) );
MUX2_X1 _19408_ ( .A(\EXU.xrd_o [30] ), .B(\RFU.rf[8][30] ), .S(_03119_ ), .Z(_01388_ ) );
MUX2_X1 _19409_ ( .A(\EXU.xrd_o [21] ), .B(\RFU.rf[8][21] ), .S(_03119_ ), .Z(_01389_ ) );
MUX2_X1 _19410_ ( .A(\EXU.xrd_o [20] ), .B(\RFU.rf[8][20] ), .S(_03119_ ), .Z(_01390_ ) );
MUX2_X1 _19411_ ( .A(\EXU.xrd_o [19] ), .B(\RFU.rf[8][19] ), .S(_03119_ ), .Z(_01391_ ) );
MUX2_X1 _19412_ ( .A(\EXU.xrd_o [18] ), .B(\RFU.rf[8][18] ), .S(_03119_ ), .Z(_01392_ ) );
MUX2_X1 _19413_ ( .A(\EXU.xrd_o [17] ), .B(\RFU.rf[8][17] ), .S(_03119_ ), .Z(_01393_ ) );
MUX2_X1 _19414_ ( .A(\EXU.xrd_o [16] ), .B(\RFU.rf[8][16] ), .S(_03119_ ), .Z(_01394_ ) );
MUX2_X1 _19415_ ( .A(\EXU.xrd_o [15] ), .B(\RFU.rf[8][15] ), .S(_03119_ ), .Z(_01395_ ) );
MUX2_X1 _19416_ ( .A(\EXU.xrd_o [14] ), .B(\RFU.rf[8][14] ), .S(_03119_ ), .Z(_01396_ ) );
BUF_X4 _19417_ ( .A(_03118_ ), .Z(_03120_ ) );
MUX2_X1 _19418_ ( .A(\EXU.xrd_o [13] ), .B(\RFU.rf[8][13] ), .S(_03120_ ), .Z(_01397_ ) );
MUX2_X1 _19419_ ( .A(\EXU.xrd_o [12] ), .B(\RFU.rf[8][12] ), .S(_03120_ ), .Z(_01398_ ) );
MUX2_X1 _19420_ ( .A(\EXU.xrd_o [29] ), .B(\RFU.rf[8][29] ), .S(_03120_ ), .Z(_01399_ ) );
MUX2_X1 _19421_ ( .A(\EXU.xrd_o [11] ), .B(\RFU.rf[8][11] ), .S(_03120_ ), .Z(_01400_ ) );
MUX2_X1 _19422_ ( .A(\EXU.xrd_o [10] ), .B(\RFU.rf[8][10] ), .S(_03120_ ), .Z(_01401_ ) );
MUX2_X1 _19423_ ( .A(\EXU.xrd_o [9] ), .B(\RFU.rf[8][9] ), .S(_03120_ ), .Z(_01402_ ) );
MUX2_X1 _19424_ ( .A(\EXU.xrd_o [8] ), .B(\RFU.rf[8][8] ), .S(_03120_ ), .Z(_01403_ ) );
MUX2_X1 _19425_ ( .A(\EXU.xrd_o [7] ), .B(\RFU.rf[8][7] ), .S(_03120_ ), .Z(_01404_ ) );
MUX2_X1 _19426_ ( .A(\EXU.xrd_o [6] ), .B(\RFU.rf[8][6] ), .S(_03120_ ), .Z(_01405_ ) );
MUX2_X1 _19427_ ( .A(\EXU.xrd_o [5] ), .B(\RFU.rf[8][5] ), .S(_03120_ ), .Z(_01406_ ) );
BUF_X4 _19428_ ( .A(_03118_ ), .Z(_03121_ ) );
MUX2_X1 _19429_ ( .A(\EXU.xrd_o [4] ), .B(\RFU.rf[8][4] ), .S(_03121_ ), .Z(_01407_ ) );
MUX2_X1 _19430_ ( .A(\EXU.xrd_o [3] ), .B(\RFU.rf[8][3] ), .S(_03121_ ), .Z(_01408_ ) );
MUX2_X1 _19431_ ( .A(\EXU.xrd_o [2] ), .B(\RFU.rf[8][2] ), .S(_03121_ ), .Z(_01409_ ) );
MUX2_X1 _19432_ ( .A(\EXU.xrd_o [28] ), .B(\RFU.rf[8][28] ), .S(_03121_ ), .Z(_01410_ ) );
MUX2_X1 _19433_ ( .A(\EXU.xrd_o [1] ), .B(\RFU.rf[8][1] ), .S(_03121_ ), .Z(_01411_ ) );
MUX2_X1 _19434_ ( .A(\EXU.xrd_o [0] ), .B(\RFU.rf[8][0] ), .S(_03121_ ), .Z(_01412_ ) );
MUX2_X1 _19435_ ( .A(\EXU.xrd_o [27] ), .B(\RFU.rf[8][27] ), .S(_03121_ ), .Z(_01413_ ) );
MUX2_X1 _19436_ ( .A(\EXU.xrd_o [26] ), .B(\RFU.rf[8][26] ), .S(_03121_ ), .Z(_01414_ ) );
MUX2_X1 _19437_ ( .A(\EXU.xrd_o [25] ), .B(\RFU.rf[8][25] ), .S(_03121_ ), .Z(_01415_ ) );
MUX2_X1 _19438_ ( .A(\EXU.xrd_o [24] ), .B(\RFU.rf[8][24] ), .S(_03121_ ), .Z(_01416_ ) );
MUX2_X1 _19439_ ( .A(\EXU.xrd_o [23] ), .B(\RFU.rf[8][23] ), .S(_03118_ ), .Z(_01417_ ) );
MUX2_X1 _19440_ ( .A(\EXU.xrd_o [22] ), .B(\RFU.rf[8][22] ), .S(_03118_ ), .Z(_01418_ ) );
AND4_X1 _19441_ ( .A1(\EXU.rd_o [3] ), .A2(_05430_ ), .A3(_05432_ ), .A4(\EXU.rd_o [0] ), .ZN(_03122_ ) );
AND2_X2 _19442_ ( .A1(_03051_ ), .A2(_03122_ ), .ZN(_03123_ ) );
BUF_X4 _19443_ ( .A(_03123_ ), .Z(_03124_ ) );
MUX2_X1 _19444_ ( .A(\RFU.rf[9][31] ), .B(\EXU.xrd_o [31] ), .S(_03124_ ), .Z(_01419_ ) );
MUX2_X1 _19445_ ( .A(\RFU.rf[9][30] ), .B(\EXU.xrd_o [30] ), .S(_03124_ ), .Z(_01420_ ) );
MUX2_X1 _19446_ ( .A(\RFU.rf[9][21] ), .B(\EXU.xrd_o [21] ), .S(_03124_ ), .Z(_01421_ ) );
MUX2_X1 _19447_ ( .A(\RFU.rf[9][20] ), .B(\EXU.xrd_o [20] ), .S(_03124_ ), .Z(_01422_ ) );
MUX2_X1 _19448_ ( .A(\RFU.rf[9][19] ), .B(\EXU.xrd_o [19] ), .S(_03124_ ), .Z(_01423_ ) );
MUX2_X1 _19449_ ( .A(\RFU.rf[9][18] ), .B(\EXU.xrd_o [18] ), .S(_03124_ ), .Z(_01424_ ) );
MUX2_X1 _19450_ ( .A(\RFU.rf[9][17] ), .B(\EXU.xrd_o [17] ), .S(_03124_ ), .Z(_01425_ ) );
MUX2_X1 _19451_ ( .A(\RFU.rf[9][16] ), .B(\EXU.xrd_o [16] ), .S(_03124_ ), .Z(_01426_ ) );
MUX2_X1 _19452_ ( .A(\RFU.rf[9][15] ), .B(\EXU.xrd_o [15] ), .S(_03124_ ), .Z(_01427_ ) );
MUX2_X1 _19453_ ( .A(\RFU.rf[9][14] ), .B(\EXU.xrd_o [14] ), .S(_03124_ ), .Z(_01428_ ) );
BUF_X4 _19454_ ( .A(_03123_ ), .Z(_03125_ ) );
MUX2_X1 _19455_ ( .A(\RFU.rf[9][13] ), .B(\EXU.xrd_o [13] ), .S(_03125_ ), .Z(_01429_ ) );
MUX2_X1 _19456_ ( .A(\RFU.rf[9][12] ), .B(\EXU.xrd_o [12] ), .S(_03125_ ), .Z(_01430_ ) );
MUX2_X1 _19457_ ( .A(\RFU.rf[9][29] ), .B(\EXU.xrd_o [29] ), .S(_03125_ ), .Z(_01431_ ) );
MUX2_X1 _19458_ ( .A(\RFU.rf[9][11] ), .B(\EXU.xrd_o [11] ), .S(_03125_ ), .Z(_01432_ ) );
MUX2_X1 _19459_ ( .A(\RFU.rf[9][10] ), .B(\EXU.xrd_o [10] ), .S(_03125_ ), .Z(_01433_ ) );
MUX2_X1 _19460_ ( .A(\RFU.rf[9][9] ), .B(\EXU.xrd_o [9] ), .S(_03125_ ), .Z(_01434_ ) );
MUX2_X1 _19461_ ( .A(\RFU.rf[9][8] ), .B(\EXU.xrd_o [8] ), .S(_03125_ ), .Z(_01435_ ) );
MUX2_X1 _19462_ ( .A(\RFU.rf[9][7] ), .B(\EXU.xrd_o [7] ), .S(_03125_ ), .Z(_01436_ ) );
MUX2_X1 _19463_ ( .A(\RFU.rf[9][6] ), .B(\EXU.xrd_o [6] ), .S(_03125_ ), .Z(_01437_ ) );
MUX2_X1 _19464_ ( .A(\RFU.rf[9][5] ), .B(\EXU.xrd_o [5] ), .S(_03125_ ), .Z(_01438_ ) );
BUF_X4 _19465_ ( .A(_03123_ ), .Z(_03126_ ) );
MUX2_X1 _19466_ ( .A(\RFU.rf[9][4] ), .B(\EXU.xrd_o [4] ), .S(_03126_ ), .Z(_01439_ ) );
MUX2_X1 _19467_ ( .A(\RFU.rf[9][3] ), .B(\EXU.xrd_o [3] ), .S(_03126_ ), .Z(_01440_ ) );
MUX2_X1 _19468_ ( .A(\RFU.rf[9][2] ), .B(\EXU.xrd_o [2] ), .S(_03126_ ), .Z(_01441_ ) );
MUX2_X1 _19469_ ( .A(\RFU.rf[9][28] ), .B(\EXU.xrd_o [28] ), .S(_03126_ ), .Z(_01442_ ) );
MUX2_X1 _19470_ ( .A(\RFU.rf[9][1] ), .B(\EXU.xrd_o [1] ), .S(_03126_ ), .Z(_01443_ ) );
MUX2_X1 _19471_ ( .A(\RFU.rf[9][0] ), .B(\EXU.xrd_o [0] ), .S(_03126_ ), .Z(_01444_ ) );
MUX2_X1 _19472_ ( .A(\RFU.rf[9][27] ), .B(\EXU.xrd_o [27] ), .S(_03126_ ), .Z(_01445_ ) );
MUX2_X1 _19473_ ( .A(\RFU.rf[9][26] ), .B(\EXU.xrd_o [26] ), .S(_03126_ ), .Z(_01446_ ) );
MUX2_X1 _19474_ ( .A(\RFU.rf[9][25] ), .B(\EXU.xrd_o [25] ), .S(_03126_ ), .Z(_01447_ ) );
MUX2_X1 _19475_ ( .A(\RFU.rf[9][24] ), .B(\EXU.xrd_o [24] ), .S(_03126_ ), .Z(_01448_ ) );
MUX2_X1 _19476_ ( .A(\RFU.rf[9][23] ), .B(\EXU.xrd_o [23] ), .S(_03123_ ), .Z(_01449_ ) );
MUX2_X1 _19477_ ( .A(\RFU.rf[9][22] ), .B(\EXU.xrd_o [22] ), .S(_03123_ ), .Z(_01450_ ) );
MUX2_X1 _19478_ ( .A(\ICACHE.s_axi_araddr [15] ), .B(_07636_ ), .S(_03833_ ), .Z(_00515_ ) );
MUX2_X1 _19479_ ( .A(\ICACHE.s_axi_araddr [14] ), .B(_07586_ ), .S(_03833_ ), .Z(_00516_ ) );
NOR2_X1 _19480_ ( .A1(_03833_ ), .A2(\ICACHE.s_axi_araddr [5] ), .ZN(_03127_ ) );
CLKBUF_X2 _19481_ ( .A(_03808_ ), .Z(\CLINT.c_axi_arready_$_DFF_P__Q_D ) );
AOI21_X1 _19482_ ( .A(_03127_ ), .B1(_07607_ ), .B2(\CLINT.c_axi_arready_$_DFF_P__Q_D ), .ZN(_00517_ ) );
OAI21_X1 _19483_ ( .A(_07796_ ), .B1(\CLINT.c_axi_arready_$_DFF_P__Q_D ), .B2(_07549_ ), .ZN(_00518_ ) );
MUX2_X1 _19484_ ( .A(\ICACHE.s_axi_araddr [3] ), .B(_01600_ ), .S(_03833_ ), .Z(_00519_ ) );
MUX2_X1 _19485_ ( .A(\ICACHE.s_axi_araddr [2] ), .B(_01601_ ), .S(_03833_ ), .Z(_00520_ ) );
MUX2_X1 _19486_ ( .A(\ICACHE.s_axi_araddr [13] ), .B(_07595_ ), .S(_03844_ ), .Z(_00521_ ) );
NAND2_X1 _19487_ ( .A1(fanout_net_11 ), .A2(\ICACHE.s_axi_araddr [12] ), .ZN(_03128_ ) );
OAI21_X1 _19488_ ( .A(_03128_ ), .B1(_07613_ ), .B2(fanout_net_11 ), .ZN(_00522_ ) );
NAND2_X1 _19489_ ( .A1(fanout_net_11 ), .A2(\ICACHE.s_axi_araddr [11] ), .ZN(_03129_ ) );
OAI21_X1 _19490_ ( .A(_03129_ ), .B1(_07620_ ), .B2(fanout_net_11 ), .ZN(_00523_ ) );
MUX2_X1 _19491_ ( .A(\ICACHE.s_axi_araddr [10] ), .B(_07579_ ), .S(_03844_ ), .Z(_00524_ ) );
MUX2_X1 _19492_ ( .A(\ICACHE.s_axi_araddr [9] ), .B(_07628_ ), .S(_03844_ ), .Z(_00525_ ) );
MUX2_X1 _19493_ ( .A(\ICACHE.s_axi_araddr [8] ), .B(_07564_ ), .S(_03844_ ), .Z(_00526_ ) );
MUX2_X1 _19494_ ( .A(\ICACHE.s_axi_araddr [7] ), .B(_07571_ ), .S(_03844_ ), .Z(_00527_ ) );
MUX2_X1 _19495_ ( .A(\ICACHE.s_axi_araddr [6] ), .B(_07557_ ), .S(_03844_ ), .Z(_00528_ ) );
INV_X1 _19496_ ( .A(\CLINT.c_axi_rvalid ), .ZN(_03130_ ) );
OR2_X1 _19497_ ( .A1(_07831_ ), .A2(\LSU.ls_axi_rready_$_NOT__A_Y ), .ZN(_03131_ ) );
OR3_X1 _19498_ ( .A1(_04055_ ), .A2(\ICACHE.m_axi_arready ), .A3(\Xbar.state [2] ), .ZN(_03132_ ) );
AND2_X1 _19499_ ( .A1(_03131_ ), .A2(_03132_ ), .ZN(_03133_ ) );
NOR3_X1 _19500_ ( .A1(_07540_ ), .A2(_03130_ ), .A3(_03133_ ), .ZN(_03134_ ) );
NOR2_X1 _19501_ ( .A1(_04106_ ), .A2(_04107_ ), .ZN(_03135_ ) );
AOI211_X1 _19502_ ( .A(_03135_ ), .B(_03001_ ), .C1(_03002_ ), .C2(_03003_ ), .ZN(_03136_ ) );
NAND2_X1 _19503_ ( .A1(_03136_ ), .A2(\CLINT.c_axi_arready ), .ZN(_03137_ ) );
AOI211_X1 _19504_ ( .A(fanout_net_11 ), .B(_03134_ ), .C1(_03137_ ), .C2(_03130_ ), .ZN(_00132_ ) );
AND2_X4 _19505_ ( .A1(\CLINT.mtime [1] ), .A2(\CLINT.mtime [0] ), .ZN(_03138_ ) );
AND2_X4 _19506_ ( .A1(_03138_ ), .A2(\CLINT.mtime [2] ), .ZN(_03139_ ) );
AND2_X4 _19507_ ( .A1(_03139_ ), .A2(\CLINT.mtime [3] ), .ZN(_03140_ ) );
AND2_X1 _19508_ ( .A1(\CLINT.mtime [5] ), .A2(\CLINT.mtime [4] ), .ZN(_03141_ ) );
AND2_X4 _19509_ ( .A1(_03140_ ), .A2(_03141_ ), .ZN(_03142_ ) );
AND2_X4 _19510_ ( .A1(_03142_ ), .A2(\CLINT.mtime [6] ), .ZN(_03143_ ) );
AND2_X4 _19511_ ( .A1(_03143_ ), .A2(\CLINT.mtime [7] ), .ZN(_03144_ ) );
AND4_X1 _19512_ ( .A1(\CLINT.mtime [15] ), .A2(\CLINT.mtime [14] ), .A3(\CLINT.mtime [13] ), .A4(\CLINT.mtime [12] ), .ZN(_03145_ ) );
AND2_X1 _19513_ ( .A1(\CLINT.mtime [9] ), .A2(\CLINT.mtime [8] ), .ZN(_03146_ ) );
AND4_X1 _19514_ ( .A1(\CLINT.mtime [11] ), .A2(_03145_ ), .A3(\CLINT.mtime [10] ), .A4(_03146_ ), .ZN(_03147_ ) );
AND2_X1 _19515_ ( .A1(_03144_ ), .A2(_03147_ ), .ZN(_03148_ ) );
AND2_X1 _19516_ ( .A1(\CLINT.mtime [29] ), .A2(\CLINT.mtime [28] ), .ZN(_03149_ ) );
AND3_X1 _19517_ ( .A1(_03149_ ), .A2(\CLINT.mtime [30] ), .A3(\CLINT.mtime [31] ), .ZN(_03150_ ) );
AND2_X1 _19518_ ( .A1(\CLINT.mtime [25] ), .A2(\CLINT.mtime [24] ), .ZN(_03151_ ) );
AND3_X1 _19519_ ( .A1(_03151_ ), .A2(\CLINT.mtime [27] ), .A3(\CLINT.mtime [26] ), .ZN(_03152_ ) );
AND4_X1 _19520_ ( .A1(\CLINT.mtime [21] ), .A2(\CLINT.mtime [20] ), .A3(\CLINT.mtime [23] ), .A4(\CLINT.mtime [22] ), .ZN(_03153_ ) );
NAND2_X1 _19521_ ( .A1(\CLINT.mtime [19] ), .A2(\CLINT.mtime [18] ), .ZN(_03154_ ) );
INV_X1 _19522_ ( .A(\CLINT.mtime [17] ), .ZN(_03155_ ) );
INV_X1 _19523_ ( .A(\CLINT.mtime [16] ), .ZN(_03156_ ) );
NOR3_X1 _19524_ ( .A1(_03154_ ), .A2(_03155_ ), .A3(_03156_ ), .ZN(_03157_ ) );
AND4_X2 _19525_ ( .A1(_03150_ ), .A2(_03152_ ), .A3(_03153_ ), .A4(_03157_ ), .ZN(_03158_ ) );
AND2_X2 _19526_ ( .A1(_03148_ ), .A2(_03158_ ), .ZN(_03159_ ) );
AND2_X1 _19527_ ( .A1(\CLINT.mtime [45] ), .A2(\CLINT.mtime [44] ), .ZN(_03160_ ) );
AND3_X1 _19528_ ( .A1(_03160_ ), .A2(\CLINT.mtime [47] ), .A3(\CLINT.mtime [46] ), .ZN(_03161_ ) );
AND2_X1 _19529_ ( .A1(\CLINT.mtime [41] ), .A2(\CLINT.mtime [40] ), .ZN(_03162_ ) );
AND3_X1 _19530_ ( .A1(_03162_ ), .A2(\CLINT.mtime [43] ), .A3(\CLINT.mtime [42] ), .ZN(_03163_ ) );
AND4_X1 _19531_ ( .A1(\CLINT.mtime [39] ), .A2(\CLINT.mtime [38] ), .A3(\CLINT.mtime [37] ), .A4(\CLINT.mtime [36] ), .ZN(_03164_ ) );
NAND2_X1 _19532_ ( .A1(\CLINT.mtime [33] ), .A2(\CLINT.mtime [32] ), .ZN(_03165_ ) );
INV_X1 _19533_ ( .A(\CLINT.mtime [35] ), .ZN(_03166_ ) );
INV_X1 _19534_ ( .A(\CLINT.mtime [34] ), .ZN(_03167_ ) );
NOR3_X1 _19535_ ( .A1(_03165_ ), .A2(_03166_ ), .A3(_03167_ ), .ZN(_03168_ ) );
AND4_X1 _19536_ ( .A1(_03161_ ), .A2(_03163_ ), .A3(_03164_ ), .A4(_03168_ ), .ZN(_03169_ ) );
AND2_X1 _19537_ ( .A1(_03159_ ), .A2(_03169_ ), .ZN(_03170_ ) );
AND2_X1 _19538_ ( .A1(\CLINT.mtime [51] ), .A2(\CLINT.mtime [50] ), .ZN(_03171_ ) );
NAND3_X1 _19539_ ( .A1(_03171_ ), .A2(\CLINT.mtime [49] ), .A3(\CLINT.mtime [48] ), .ZN(_03172_ ) );
NAND4_X1 _19540_ ( .A1(\CLINT.mtime [53] ), .A2(\CLINT.mtime [52] ), .A3(\CLINT.mtime [55] ), .A4(\CLINT.mtime [54] ), .ZN(_03173_ ) );
NOR2_X1 _19541_ ( .A1(_03172_ ), .A2(_03173_ ), .ZN(_03174_ ) );
AND2_X1 _19542_ ( .A1(_03170_ ), .A2(_03174_ ), .ZN(_03175_ ) );
INV_X1 _19543_ ( .A(_03175_ ), .ZN(_03176_ ) );
NAND4_X1 _19544_ ( .A1(\CLINT.mtime [59] ), .A2(\CLINT.mtime [58] ), .A3(\CLINT.mtime [57] ), .A4(\CLINT.mtime [56] ), .ZN(_03177_ ) );
NOR2_X1 _19545_ ( .A1(_03176_ ), .A2(_03177_ ), .ZN(_03178_ ) );
NAND3_X1 _19546_ ( .A1(_03178_ ), .A2(\CLINT.mtime [61] ), .A3(\CLINT.mtime [60] ), .ZN(_03179_ ) );
INV_X1 _19547_ ( .A(\CLINT.mtime [62] ), .ZN(_03180_ ) );
OR3_X1 _19548_ ( .A1(_03179_ ), .A2(_03180_ ), .A3(\CLINT.mtime [63] ), .ZN(_03181_ ) );
OAI21_X1 _19549_ ( .A(\CLINT.mtime [63] ), .B1(_03179_ ), .B2(_03180_ ), .ZN(_03182_ ) );
AOI21_X1 _19550_ ( .A(fanout_net_11 ), .B1(_03181_ ), .B2(_03182_ ), .ZN(_00133_ ) );
NAND2_X1 _19551_ ( .A1(_03179_ ), .A2(\CLINT.mtime [62] ), .ZN(_03183_ ) );
NAND4_X1 _19552_ ( .A1(_03178_ ), .A2(_03180_ ), .A3(\CLINT.mtime [61] ), .A4(\CLINT.mtime [60] ), .ZN(_03184_ ) );
AOI21_X1 _19553_ ( .A(fanout_net_11 ), .B1(_03183_ ), .B2(_03184_ ), .ZN(_00134_ ) );
INV_X1 _19554_ ( .A(_03170_ ), .ZN(_03185_ ) );
INV_X1 _19555_ ( .A(\CLINT.mtime [52] ), .ZN(_03186_ ) );
OR3_X1 _19556_ ( .A1(_03185_ ), .A2(_03186_ ), .A3(_03172_ ), .ZN(_03187_ ) );
NAND2_X1 _19557_ ( .A1(_03187_ ), .A2(\CLINT.mtime [53] ), .ZN(_03188_ ) );
OR4_X1 _19558_ ( .A1(\CLINT.mtime [53] ), .A2(_03185_ ), .A3(_03186_ ), .A4(_03172_ ), .ZN(_03189_ ) );
AOI21_X1 _19559_ ( .A(fanout_net_11 ), .B1(_03188_ ), .B2(_03189_ ), .ZN(_00135_ ) );
INV_X1 _19560_ ( .A(_03159_ ), .ZN(_03190_ ) );
INV_X1 _19561_ ( .A(_03169_ ), .ZN(_03191_ ) );
OR4_X1 _19562_ ( .A1(\CLINT.mtime [52] ), .A2(_03190_ ), .A3(_03191_ ), .A4(_03172_ ), .ZN(_03192_ ) );
OAI21_X1 _19563_ ( .A(\CLINT.mtime [52] ), .B1(_03185_ ), .B2(_03172_ ), .ZN(_03193_ ) );
AOI21_X1 _19564_ ( .A(fanout_net_11 ), .B1(_03192_ ), .B2(_03193_ ), .ZN(_00136_ ) );
NAND3_X1 _19565_ ( .A1(_03170_ ), .A2(\CLINT.mtime [49] ), .A3(\CLINT.mtime [48] ), .ZN(_03194_ ) );
INV_X1 _19566_ ( .A(\CLINT.mtime [50] ), .ZN(_03195_ ) );
OR3_X1 _19567_ ( .A1(_03194_ ), .A2(\CLINT.mtime [51] ), .A3(_03195_ ), .ZN(_03196_ ) );
OAI21_X1 _19568_ ( .A(\CLINT.mtime [51] ), .B1(_03194_ ), .B2(_03195_ ), .ZN(_03197_ ) );
AOI21_X1 _19569_ ( .A(fanout_net_11 ), .B1(_03196_ ), .B2(_03197_ ), .ZN(_00137_ ) );
NAND2_X1 _19570_ ( .A1(_03194_ ), .A2(\CLINT.mtime [50] ), .ZN(_03198_ ) );
NAND4_X1 _19571_ ( .A1(_03170_ ), .A2(_03195_ ), .A3(\CLINT.mtime [49] ), .A4(\CLINT.mtime [48] ), .ZN(_03199_ ) );
AOI21_X1 _19572_ ( .A(fanout_net_11 ), .B1(_03198_ ), .B2(_03199_ ), .ZN(_00138_ ) );
INV_X1 _19573_ ( .A(\CLINT.mtime [48] ), .ZN(_03200_ ) );
OR4_X1 _19574_ ( .A1(\CLINT.mtime [49] ), .A2(_03190_ ), .A3(_03200_ ), .A4(_03191_ ), .ZN(_03201_ ) );
NAND3_X1 _19575_ ( .A1(_03159_ ), .A2(\CLINT.mtime [48] ), .A3(_03169_ ), .ZN(_03202_ ) );
NAND2_X1 _19576_ ( .A1(_03202_ ), .A2(\CLINT.mtime [49] ), .ZN(_03203_ ) );
AOI21_X1 _19577_ ( .A(fanout_net_11 ), .B1(_03201_ ), .B2(_03203_ ), .ZN(_00139_ ) );
OAI21_X1 _19578_ ( .A(\CLINT.mtime [48] ), .B1(_03190_ ), .B2(_03191_ ), .ZN(_03204_ ) );
BUF_X2 _19579_ ( .A(_03148_ ), .Z(_03205_ ) );
NAND4_X1 _19580_ ( .A1(_03205_ ), .A2(_03200_ ), .A3(_03158_ ), .A4(_03169_ ), .ZN(_03206_ ) );
AOI21_X1 _19581_ ( .A(fanout_net_11 ), .B1(_03204_ ), .B2(_03206_ ), .ZN(_00140_ ) );
AND2_X1 _19582_ ( .A1(_03168_ ), .A2(_03164_ ), .ZN(_03207_ ) );
AND2_X2 _19583_ ( .A1(_03159_ ), .A2(_03207_ ), .ZN(_03208_ ) );
NAND3_X1 _19584_ ( .A1(_03208_ ), .A2(_03160_ ), .A3(_03163_ ), .ZN(_03209_ ) );
INV_X1 _19585_ ( .A(\CLINT.mtime [46] ), .ZN(_03210_ ) );
OR3_X1 _19586_ ( .A1(_03209_ ), .A2(\CLINT.mtime [47] ), .A3(_03210_ ), .ZN(_03211_ ) );
OAI21_X1 _19587_ ( .A(\CLINT.mtime [47] ), .B1(_03209_ ), .B2(_03210_ ), .ZN(_03212_ ) );
AOI21_X1 _19588_ ( .A(fanout_net_11 ), .B1(_03211_ ), .B2(_03212_ ), .ZN(_00141_ ) );
NAND2_X1 _19589_ ( .A1(_03209_ ), .A2(\CLINT.mtime [46] ), .ZN(_03213_ ) );
NAND4_X1 _19590_ ( .A1(_03208_ ), .A2(_03210_ ), .A3(_03160_ ), .A4(_03163_ ), .ZN(_03214_ ) );
AOI21_X1 _19591_ ( .A(fanout_net_11 ), .B1(_03213_ ), .B2(_03214_ ), .ZN(_00142_ ) );
NAND3_X1 _19592_ ( .A1(_03208_ ), .A2(\CLINT.mtime [44] ), .A3(_03163_ ), .ZN(_03215_ ) );
OR2_X1 _19593_ ( .A1(_03215_ ), .A2(\CLINT.mtime [45] ), .ZN(_03216_ ) );
NAND2_X1 _19594_ ( .A1(_03215_ ), .A2(\CLINT.mtime [45] ), .ZN(_03217_ ) );
AOI21_X1 _19595_ ( .A(fanout_net_11 ), .B1(_03216_ ), .B2(_03217_ ), .ZN(_00143_ ) );
NAND2_X1 _19596_ ( .A1(_03208_ ), .A2(_03163_ ), .ZN(_03218_ ) );
OR2_X1 _19597_ ( .A1(_03218_ ), .A2(\CLINT.mtime [44] ), .ZN(_03219_ ) );
NAND2_X1 _19598_ ( .A1(_03218_ ), .A2(\CLINT.mtime [44] ), .ZN(_03220_ ) );
AOI21_X1 _19599_ ( .A(fanout_net_11 ), .B1(_03219_ ), .B2(_03220_ ), .ZN(_00144_ ) );
AND3_X1 _19600_ ( .A1(_03146_ ), .A2(\CLINT.mtime [11] ), .A3(\CLINT.mtime [10] ), .ZN(_03221_ ) );
AND2_X4 _19601_ ( .A1(_03144_ ), .A2(_03221_ ), .ZN(_03222_ ) );
AND2_X4 _19602_ ( .A1(_03222_ ), .A2(\CLINT.mtime [12] ), .ZN(_03223_ ) );
AND2_X4 _19603_ ( .A1(_03223_ ), .A2(\CLINT.mtime [13] ), .ZN(_03224_ ) );
AND3_X4 _19604_ ( .A1(_03224_ ), .A2(\CLINT.mtime [15] ), .A3(\CLINT.mtime [14] ), .ZN(_03225_ ) );
AND3_X4 _19605_ ( .A1(_03225_ ), .A2(\CLINT.mtime [17] ), .A3(\CLINT.mtime [16] ), .ZN(_03226_ ) );
AND3_X4 _19606_ ( .A1(_03226_ ), .A2(\CLINT.mtime [19] ), .A3(\CLINT.mtime [18] ), .ZN(_03227_ ) );
AND2_X4 _19607_ ( .A1(_03227_ ), .A2(\CLINT.mtime [20] ), .ZN(_03228_ ) );
AND2_X2 _19608_ ( .A1(_03228_ ), .A2(\CLINT.mtime [21] ), .ZN(_03229_ ) );
AND3_X2 _19609_ ( .A1(_03229_ ), .A2(\CLINT.mtime [23] ), .A3(\CLINT.mtime [22] ), .ZN(_03230_ ) );
AND3_X2 _19610_ ( .A1(_03230_ ), .A2(\CLINT.mtime [25] ), .A3(\CLINT.mtime [24] ), .ZN(_03231_ ) );
AND2_X2 _19611_ ( .A1(_03231_ ), .A2(\CLINT.mtime [26] ), .ZN(_03232_ ) );
NAND3_X1 _19612_ ( .A1(_03232_ ), .A2(\CLINT.mtime [27] ), .A3(_03150_ ), .ZN(_03233_ ) );
INV_X1 _19613_ ( .A(\CLINT.mtime [32] ), .ZN(_03234_ ) );
NOR2_X1 _19614_ ( .A1(_03233_ ), .A2(_03234_ ), .ZN(_03235_ ) );
AND3_X2 _19615_ ( .A1(_03235_ ), .A2(\CLINT.mtime [34] ), .A3(\CLINT.mtime [33] ), .ZN(_03236_ ) );
AND3_X2 _19616_ ( .A1(_03236_ ), .A2(\CLINT.mtime [36] ), .A3(\CLINT.mtime [35] ), .ZN(_03237_ ) );
AND2_X2 _19617_ ( .A1(_03237_ ), .A2(\CLINT.mtime [37] ), .ZN(_03238_ ) );
AND3_X2 _19618_ ( .A1(_03238_ ), .A2(\CLINT.mtime [39] ), .A3(\CLINT.mtime [38] ), .ZN(_03239_ ) );
AND3_X2 _19619_ ( .A1(_03239_ ), .A2(\CLINT.mtime [41] ), .A3(\CLINT.mtime [40] ), .ZN(_03240_ ) );
AND2_X2 _19620_ ( .A1(_03240_ ), .A2(\CLINT.mtime [42] ), .ZN(_03241_ ) );
NAND3_X1 _19621_ ( .A1(_03241_ ), .A2(\CLINT.mtime [43] ), .A3(_03161_ ), .ZN(_03242_ ) );
NOR2_X1 _19622_ ( .A1(_03242_ ), .A2(_03200_ ), .ZN(_03243_ ) );
AND3_X2 _19623_ ( .A1(_03243_ ), .A2(\CLINT.mtime [50] ), .A3(\CLINT.mtime [49] ), .ZN(_03244_ ) );
AND2_X1 _19624_ ( .A1(\CLINT.mtime [53] ), .A2(\CLINT.mtime [52] ), .ZN(_03245_ ) );
AND3_X4 _19625_ ( .A1(_03244_ ), .A2(\CLINT.mtime [51] ), .A3(_03245_ ), .ZN(_03246_ ) );
AND3_X4 _19626_ ( .A1(_03246_ ), .A2(\CLINT.mtime [55] ), .A3(\CLINT.mtime [54] ), .ZN(_03247_ ) );
AND3_X4 _19627_ ( .A1(_03247_ ), .A2(\CLINT.mtime [57] ), .A3(\CLINT.mtime [56] ), .ZN(_03248_ ) );
AND3_X4 _19628_ ( .A1(_03248_ ), .A2(\CLINT.mtime [59] ), .A3(\CLINT.mtime [58] ), .ZN(_03249_ ) );
AND3_X2 _19629_ ( .A1(_03249_ ), .A2(\CLINT.mtime [61] ), .A3(\CLINT.mtime [60] ), .ZN(_03250_ ) );
AOI21_X1 _19630_ ( .A(\CLINT.mtime [61] ), .B1(_03249_ ), .B2(\CLINT.mtime [60] ), .ZN(_03251_ ) );
NOR3_X1 _19631_ ( .A1(_03250_ ), .A2(_03251_ ), .A3(fanout_net_11 ), .ZN(_00145_ ) );
NAND3_X1 _19632_ ( .A1(_03159_ ), .A2(_03162_ ), .A3(_03207_ ), .ZN(_03252_ ) );
INV_X1 _19633_ ( .A(\CLINT.mtime [42] ), .ZN(_03253_ ) );
NOR2_X1 _19634_ ( .A1(_03252_ ), .A2(_03253_ ), .ZN(_03254_ ) );
XNOR2_X1 _19635_ ( .A(_03254_ ), .B(\CLINT.mtime [43] ), .ZN(_03255_ ) );
NOR2_X1 _19636_ ( .A1(_03255_ ), .A2(fanout_net_11 ), .ZN(_00146_ ) );
NAND2_X1 _19637_ ( .A1(_03252_ ), .A2(\CLINT.mtime [42] ), .ZN(_03256_ ) );
NAND4_X1 _19638_ ( .A1(_03159_ ), .A2(_03253_ ), .A3(_03162_ ), .A4(_03207_ ), .ZN(_03257_ ) );
AOI21_X1 _19639_ ( .A(fanout_net_11 ), .B1(_03256_ ), .B2(_03257_ ), .ZN(_00147_ ) );
NAND3_X1 _19640_ ( .A1(_03159_ ), .A2(\CLINT.mtime [40] ), .A3(_03207_ ), .ZN(_03258_ ) );
XNOR2_X1 _19641_ ( .A(_03258_ ), .B(\CLINT.mtime [41] ), .ZN(_03259_ ) );
AND2_X1 _19642_ ( .A1(_03259_ ), .A2(\CLINT.c_axi_arready_$_DFF_P__Q_D ), .ZN(_00148_ ) );
XNOR2_X1 _19643_ ( .A(_03208_ ), .B(\CLINT.mtime [40] ), .ZN(_03260_ ) );
NOR2_X1 _19644_ ( .A1(_03260_ ), .A2(fanout_net_11 ), .ZN(_00149_ ) );
AND2_X1 _19645_ ( .A1(_03159_ ), .A2(_03168_ ), .ZN(_03261_ ) );
NAND3_X1 _19646_ ( .A1(_03261_ ), .A2(\CLINT.mtime [37] ), .A3(\CLINT.mtime [36] ), .ZN(_03262_ ) );
INV_X1 _19647_ ( .A(\CLINT.mtime [38] ), .ZN(_03263_ ) );
OR3_X1 _19648_ ( .A1(_03262_ ), .A2(\CLINT.mtime [39] ), .A3(_03263_ ), .ZN(_03264_ ) );
OAI21_X1 _19649_ ( .A(\CLINT.mtime [39] ), .B1(_03262_ ), .B2(_03263_ ), .ZN(_03265_ ) );
AOI21_X1 _19650_ ( .A(fanout_net_11 ), .B1(_03264_ ), .B2(_03265_ ), .ZN(_00150_ ) );
NAND2_X1 _19651_ ( .A1(_03262_ ), .A2(\CLINT.mtime [38] ), .ZN(_03266_ ) );
NAND4_X1 _19652_ ( .A1(_03261_ ), .A2(_03263_ ), .A3(\CLINT.mtime [37] ), .A4(\CLINT.mtime [36] ), .ZN(_03267_ ) );
AOI21_X1 _19653_ ( .A(fanout_net_11 ), .B1(_03266_ ), .B2(_03267_ ), .ZN(_00151_ ) );
NAND3_X1 _19654_ ( .A1(_03159_ ), .A2(\CLINT.mtime [36] ), .A3(_03168_ ), .ZN(_03268_ ) );
XNOR2_X1 _19655_ ( .A(_03268_ ), .B(\CLINT.mtime [37] ), .ZN(_03269_ ) );
AND2_X1 _19656_ ( .A1(_03269_ ), .A2(\CLINT.c_axi_arready_$_DFF_P__Q_D ), .ZN(_00152_ ) );
XNOR2_X1 _19657_ ( .A(_03261_ ), .B(\CLINT.mtime [36] ), .ZN(_03270_ ) );
NOR2_X1 _19658_ ( .A1(_03270_ ), .A2(fanout_net_11 ), .ZN(_00153_ ) );
INV_X1 _19659_ ( .A(_03205_ ), .ZN(_03271_ ) );
INV_X1 _19660_ ( .A(_03158_ ), .ZN(_03272_ ) );
NOR3_X1 _19661_ ( .A1(_03271_ ), .A2(_03272_ ), .A3(_03165_ ), .ZN(_03273_ ) );
NAND2_X1 _19662_ ( .A1(_03273_ ), .A2(\CLINT.mtime [34] ), .ZN(_03274_ ) );
NAND2_X1 _19663_ ( .A1(_03274_ ), .A2(\CLINT.mtime [35] ), .ZN(_03275_ ) );
NAND3_X1 _19664_ ( .A1(_03273_ ), .A2(_03166_ ), .A3(\CLINT.mtime [34] ), .ZN(_03276_ ) );
AOI21_X1 _19665_ ( .A(fanout_net_11 ), .B1(_03275_ ), .B2(_03276_ ), .ZN(_00154_ ) );
OAI21_X1 _19666_ ( .A(\CLINT.mtime [34] ), .B1(_03190_ ), .B2(_03165_ ), .ZN(_03277_ ) );
NAND4_X1 _19667_ ( .A1(_03159_ ), .A2(_03167_ ), .A3(\CLINT.mtime [33] ), .A4(\CLINT.mtime [32] ), .ZN(_03278_ ) );
AOI21_X1 _19668_ ( .A(fanout_net_12 ), .B1(_03277_ ), .B2(_03278_ ), .ZN(_00155_ ) );
OR3_X1 _19669_ ( .A1(_03176_ ), .A2(\CLINT.mtime [60] ), .A3(_03177_ ), .ZN(_03279_ ) );
OAI21_X1 _19670_ ( .A(\CLINT.mtime [60] ), .B1(_03176_ ), .B2(_03177_ ), .ZN(_03280_ ) );
AOI21_X1 _19671_ ( .A(fanout_net_12 ), .B1(_03279_ ), .B2(_03280_ ), .ZN(_00156_ ) );
OR4_X1 _19672_ ( .A1(\CLINT.mtime [33] ), .A2(_03271_ ), .A3(_03234_ ), .A4(_03272_ ), .ZN(_03281_ ) );
NAND3_X1 _19673_ ( .A1(_03205_ ), .A2(\CLINT.mtime [32] ), .A3(_03158_ ), .ZN(_03282_ ) );
NAND2_X1 _19674_ ( .A1(_03282_ ), .A2(\CLINT.mtime [33] ), .ZN(_03283_ ) );
AOI21_X1 _19675_ ( .A(fanout_net_12 ), .B1(_03281_ ), .B2(_03283_ ), .ZN(_00157_ ) );
OAI21_X1 _19676_ ( .A(\CLINT.mtime [32] ), .B1(_03271_ ), .B2(_03272_ ), .ZN(_03284_ ) );
NAND4_X1 _19677_ ( .A1(_03144_ ), .A2(_03234_ ), .A3(_03147_ ), .A4(_03158_ ), .ZN(_03285_ ) );
AOI21_X1 _19678_ ( .A(fanout_net_12 ), .B1(_03284_ ), .B2(_03285_ ), .ZN(_00158_ ) );
AND2_X1 _19679_ ( .A1(_03157_ ), .A2(_03153_ ), .ZN(_03286_ ) );
AND2_X2 _19680_ ( .A1(_03148_ ), .A2(_03286_ ), .ZN(_03287_ ) );
NAND3_X1 _19681_ ( .A1(_03287_ ), .A2(_03149_ ), .A3(_03152_ ), .ZN(_03288_ ) );
INV_X1 _19682_ ( .A(\CLINT.mtime [30] ), .ZN(_03289_ ) );
OR3_X1 _19683_ ( .A1(_03288_ ), .A2(_03289_ ), .A3(\CLINT.mtime [31] ), .ZN(_03290_ ) );
OAI21_X1 _19684_ ( .A(\CLINT.mtime [31] ), .B1(_03288_ ), .B2(_03289_ ), .ZN(_03291_ ) );
AOI21_X1 _19685_ ( .A(fanout_net_12 ), .B1(_03290_ ), .B2(_03291_ ), .ZN(_00159_ ) );
NAND2_X1 _19686_ ( .A1(_03288_ ), .A2(\CLINT.mtime [30] ), .ZN(_03292_ ) );
NAND4_X1 _19687_ ( .A1(_03287_ ), .A2(_03289_ ), .A3(_03149_ ), .A4(_03152_ ), .ZN(_03293_ ) );
AOI21_X1 _19688_ ( .A(fanout_net_12 ), .B1(_03292_ ), .B2(_03293_ ), .ZN(_00160_ ) );
NAND3_X1 _19689_ ( .A1(_03287_ ), .A2(\CLINT.mtime [28] ), .A3(_03152_ ), .ZN(_03294_ ) );
OR2_X1 _19690_ ( .A1(_03294_ ), .A2(\CLINT.mtime [29] ), .ZN(_03295_ ) );
NAND2_X1 _19691_ ( .A1(_03294_ ), .A2(\CLINT.mtime [29] ), .ZN(_03296_ ) );
AOI21_X1 _19692_ ( .A(fanout_net_12 ), .B1(_03295_ ), .B2(_03296_ ), .ZN(_00161_ ) );
NAND2_X1 _19693_ ( .A1(_03287_ ), .A2(_03152_ ), .ZN(_03297_ ) );
OR2_X1 _19694_ ( .A1(_03297_ ), .A2(\CLINT.mtime [28] ), .ZN(_03298_ ) );
NAND2_X1 _19695_ ( .A1(_03297_ ), .A2(\CLINT.mtime [28] ), .ZN(_03299_ ) );
AOI21_X1 _19696_ ( .A(fanout_net_12 ), .B1(_03298_ ), .B2(_03299_ ), .ZN(_00162_ ) );
NAND3_X1 _19697_ ( .A1(_03205_ ), .A2(_03151_ ), .A3(_03286_ ), .ZN(_03300_ ) );
INV_X1 _19698_ ( .A(\CLINT.mtime [26] ), .ZN(_03301_ ) );
NOR2_X1 _19699_ ( .A1(_03300_ ), .A2(_03301_ ), .ZN(_03302_ ) );
XNOR2_X1 _19700_ ( .A(_03302_ ), .B(\CLINT.mtime [27] ), .ZN(_03303_ ) );
NOR2_X1 _19701_ ( .A1(_03303_ ), .A2(fanout_net_12 ), .ZN(_00163_ ) );
NAND2_X1 _19702_ ( .A1(_03300_ ), .A2(\CLINT.mtime [26] ), .ZN(_03304_ ) );
NAND4_X1 _19703_ ( .A1(_03205_ ), .A2(_03301_ ), .A3(_03151_ ), .A4(_03286_ ), .ZN(_03305_ ) );
AOI21_X1 _19704_ ( .A(fanout_net_12 ), .B1(_03304_ ), .B2(_03305_ ), .ZN(_00164_ ) );
NAND3_X1 _19705_ ( .A1(_03205_ ), .A2(\CLINT.mtime [24] ), .A3(_03286_ ), .ZN(_03306_ ) );
XNOR2_X1 _19706_ ( .A(_03306_ ), .B(\CLINT.mtime [25] ), .ZN(_03307_ ) );
AND2_X1 _19707_ ( .A1(_03307_ ), .A2(\CLINT.c_axi_arready_$_DFF_P__Q_D ), .ZN(_00165_ ) );
XNOR2_X1 _19708_ ( .A(_03287_ ), .B(\CLINT.mtime [24] ), .ZN(_03308_ ) );
NOR2_X1 _19709_ ( .A1(_03308_ ), .A2(fanout_net_12 ), .ZN(_00166_ ) );
NAND3_X1 _19710_ ( .A1(_03175_ ), .A2(\CLINT.mtime [57] ), .A3(\CLINT.mtime [56] ), .ZN(_03309_ ) );
INV_X1 _19711_ ( .A(\CLINT.mtime [58] ), .ZN(_03310_ ) );
OR3_X1 _19712_ ( .A1(_03309_ ), .A2(\CLINT.mtime [59] ), .A3(_03310_ ), .ZN(_03311_ ) );
OAI21_X1 _19713_ ( .A(\CLINT.mtime [59] ), .B1(_03309_ ), .B2(_03310_ ), .ZN(_03312_ ) );
AOI21_X1 _19714_ ( .A(fanout_net_12 ), .B1(_03311_ ), .B2(_03312_ ), .ZN(_00167_ ) );
AND2_X1 _19715_ ( .A1(_03148_ ), .A2(_03157_ ), .ZN(_03313_ ) );
NAND3_X1 _19716_ ( .A1(_03313_ ), .A2(\CLINT.mtime [21] ), .A3(\CLINT.mtime [20] ), .ZN(_03314_ ) );
INV_X1 _19717_ ( .A(\CLINT.mtime [22] ), .ZN(_03315_ ) );
OR3_X1 _19718_ ( .A1(_03314_ ), .A2(\CLINT.mtime [23] ), .A3(_03315_ ), .ZN(_03316_ ) );
OAI21_X1 _19719_ ( .A(\CLINT.mtime [23] ), .B1(_03314_ ), .B2(_03315_ ), .ZN(_03317_ ) );
AOI21_X1 _19720_ ( .A(fanout_net_12 ), .B1(_03316_ ), .B2(_03317_ ), .ZN(_00168_ ) );
NAND2_X1 _19721_ ( .A1(_03314_ ), .A2(\CLINT.mtime [22] ), .ZN(_03318_ ) );
NAND4_X1 _19722_ ( .A1(_03313_ ), .A2(\CLINT.mtime [21] ), .A3(\CLINT.mtime [20] ), .A4(_03315_ ), .ZN(_03319_ ) );
AOI21_X1 _19723_ ( .A(fanout_net_12 ), .B1(_03318_ ), .B2(_03319_ ), .ZN(_00169_ ) );
NAND3_X1 _19724_ ( .A1(_03205_ ), .A2(\CLINT.mtime [20] ), .A3(_03157_ ), .ZN(_03320_ ) );
XNOR2_X1 _19725_ ( .A(_03320_ ), .B(\CLINT.mtime [21] ), .ZN(_03321_ ) );
AND2_X1 _19726_ ( .A1(_03321_ ), .A2(_03806_ ), .ZN(_00170_ ) );
XNOR2_X1 _19727_ ( .A(_03313_ ), .B(\CLINT.mtime [20] ), .ZN(_03322_ ) );
NOR2_X1 _19728_ ( .A1(_03322_ ), .A2(fanout_net_12 ), .ZN(_00171_ ) );
NAND3_X1 _19729_ ( .A1(_03205_ ), .A2(\CLINT.mtime [17] ), .A3(\CLINT.mtime [16] ), .ZN(_03323_ ) );
INV_X1 _19730_ ( .A(\CLINT.mtime [18] ), .ZN(_03324_ ) );
OR3_X1 _19731_ ( .A1(_03323_ ), .A2(\CLINT.mtime [19] ), .A3(_03324_ ), .ZN(_03325_ ) );
OAI21_X1 _19732_ ( .A(\CLINT.mtime [19] ), .B1(_03323_ ), .B2(_03324_ ), .ZN(_03326_ ) );
AOI21_X1 _19733_ ( .A(fanout_net_12 ), .B1(_03325_ ), .B2(_03326_ ), .ZN(_00172_ ) );
NAND2_X1 _19734_ ( .A1(_03323_ ), .A2(\CLINT.mtime [18] ), .ZN(_03327_ ) );
NAND4_X1 _19735_ ( .A1(_03205_ ), .A2(_03324_ ), .A3(\CLINT.mtime [17] ), .A4(\CLINT.mtime [16] ), .ZN(_03328_ ) );
AOI21_X1 _19736_ ( .A(fanout_net_12 ), .B1(_03327_ ), .B2(_03328_ ), .ZN(_00173_ ) );
NAND3_X1 _19737_ ( .A1(_03144_ ), .A2(\CLINT.mtime [16] ), .A3(_03147_ ), .ZN(_03329_ ) );
NAND2_X1 _19738_ ( .A1(_03329_ ), .A2(\CLINT.mtime [17] ), .ZN(_03330_ ) );
NAND4_X1 _19739_ ( .A1(_03144_ ), .A2(_03155_ ), .A3(\CLINT.mtime [16] ), .A4(_03147_ ), .ZN(_03331_ ) );
AOI21_X1 _19740_ ( .A(fanout_net_12 ), .B1(_03330_ ), .B2(_03331_ ), .ZN(_00174_ ) );
OR2_X1 _19741_ ( .A1(_03205_ ), .A2(_03156_ ), .ZN(_03332_ ) );
NAND4_X1 _19742_ ( .A1(_03143_ ), .A2(_03156_ ), .A3(\CLINT.mtime [7] ), .A4(_03147_ ), .ZN(_03333_ ) );
AOI21_X1 _19743_ ( .A(fanout_net_12 ), .B1(_03332_ ), .B2(_03333_ ), .ZN(_00175_ ) );
NAND3_X1 _19744_ ( .A1(_03222_ ), .A2(\CLINT.mtime [13] ), .A3(\CLINT.mtime [12] ), .ZN(_03334_ ) );
INV_X1 _19745_ ( .A(\CLINT.mtime [14] ), .ZN(_03335_ ) );
OR3_X1 _19746_ ( .A1(_03334_ ), .A2(\CLINT.mtime [15] ), .A3(_03335_ ), .ZN(_03336_ ) );
OAI21_X1 _19747_ ( .A(\CLINT.mtime [15] ), .B1(_03334_ ), .B2(_03335_ ), .ZN(_03337_ ) );
AOI21_X1 _19748_ ( .A(fanout_net_12 ), .B1(_03336_ ), .B2(_03337_ ), .ZN(_00176_ ) );
NAND2_X1 _19749_ ( .A1(_03334_ ), .A2(\CLINT.mtime [14] ), .ZN(_03338_ ) );
NAND4_X1 _19750_ ( .A1(_03222_ ), .A2(_03335_ ), .A3(\CLINT.mtime [13] ), .A4(\CLINT.mtime [12] ), .ZN(_03339_ ) );
AOI21_X1 _19751_ ( .A(fanout_net_12 ), .B1(_03338_ ), .B2(_03339_ ), .ZN(_00177_ ) );
NAND2_X1 _19752_ ( .A1(_03309_ ), .A2(\CLINT.mtime [58] ), .ZN(_03340_ ) );
NAND4_X1 _19753_ ( .A1(_03175_ ), .A2(_03310_ ), .A3(\CLINT.mtime [57] ), .A4(\CLINT.mtime [56] ), .ZN(_03341_ ) );
AOI21_X1 _19754_ ( .A(fanout_net_12 ), .B1(_03340_ ), .B2(_03341_ ), .ZN(_00178_ ) );
AOI21_X1 _19755_ ( .A(\CLINT.mtime [13] ), .B1(_03222_ ), .B2(\CLINT.mtime [12] ), .ZN(_03342_ ) );
NOR3_X1 _19756_ ( .A1(_03224_ ), .A2(fanout_net_12 ), .A3(_03342_ ), .ZN(_00179_ ) );
AOI21_X1 _19757_ ( .A(\CLINT.mtime [12] ), .B1(_03144_ ), .B2(_03221_ ), .ZN(_03343_ ) );
NOR3_X1 _19758_ ( .A1(_03223_ ), .A2(fanout_net_12 ), .A3(_03343_ ), .ZN(_00180_ ) );
AND2_X1 _19759_ ( .A1(_03144_ ), .A2(_03146_ ), .ZN(_03344_ ) );
AOI21_X1 _19760_ ( .A(\CLINT.mtime [11] ), .B1(_03344_ ), .B2(\CLINT.mtime [10] ), .ZN(_03345_ ) );
NOR3_X1 _19761_ ( .A1(_03345_ ), .A2(fanout_net_12 ), .A3(_03222_ ), .ZN(_00181_ ) );
XNOR2_X1 _19762_ ( .A(_03344_ ), .B(\CLINT.mtime [10] ), .ZN(_03346_ ) );
NOR2_X1 _19763_ ( .A1(_03346_ ), .A2(fanout_net_12 ), .ZN(_00182_ ) );
AND3_X1 _19764_ ( .A1(_03143_ ), .A2(\CLINT.mtime [8] ), .A3(\CLINT.mtime [7] ), .ZN(_03347_ ) );
XNOR2_X1 _19765_ ( .A(_03347_ ), .B(\CLINT.mtime [9] ), .ZN(_03348_ ) );
NOR2_X1 _19766_ ( .A1(_03348_ ), .A2(fanout_net_12 ), .ZN(_00183_ ) );
AOI21_X1 _19767_ ( .A(\CLINT.mtime [8] ), .B1(_03143_ ), .B2(\CLINT.mtime [7] ), .ZN(_03349_ ) );
NOR3_X1 _19768_ ( .A1(_03347_ ), .A2(_03349_ ), .A3(fanout_net_12 ), .ZN(_00184_ ) );
AOI21_X1 _19769_ ( .A(\CLINT.mtime [7] ), .B1(_03142_ ), .B2(\CLINT.mtime [6] ), .ZN(_03350_ ) );
NOR3_X1 _19770_ ( .A1(_03144_ ), .A2(fanout_net_12 ), .A3(_03350_ ), .ZN(_00185_ ) );
AOI21_X1 _19771_ ( .A(\CLINT.mtime [6] ), .B1(_03140_ ), .B2(_03141_ ), .ZN(_03351_ ) );
NOR3_X1 _19772_ ( .A1(_03143_ ), .A2(fanout_net_12 ), .A3(_03351_ ), .ZN(_00186_ ) );
AND3_X1 _19773_ ( .A1(_03139_ ), .A2(\CLINT.mtime [4] ), .A3(\CLINT.mtime [3] ), .ZN(_03352_ ) );
XNOR2_X1 _19774_ ( .A(_03352_ ), .B(\CLINT.mtime [5] ), .ZN(_03353_ ) );
NOR2_X1 _19775_ ( .A1(_03353_ ), .A2(fanout_net_13 ), .ZN(_00187_ ) );
AOI21_X1 _19776_ ( .A(\CLINT.mtime [4] ), .B1(_03139_ ), .B2(\CLINT.mtime [3] ), .ZN(_03354_ ) );
NOR3_X1 _19777_ ( .A1(_03352_ ), .A2(_03354_ ), .A3(fanout_net_13 ), .ZN(_00188_ ) );
NAND3_X1 _19778_ ( .A1(_03170_ ), .A2(\CLINT.mtime [56] ), .A3(_03174_ ), .ZN(_03355_ ) );
XNOR2_X1 _19779_ ( .A(_03355_ ), .B(\CLINT.mtime [57] ), .ZN(_03356_ ) );
AND2_X1 _19780_ ( .A1(_03356_ ), .A2(_03806_ ), .ZN(_00189_ ) );
AOI21_X1 _19781_ ( .A(\CLINT.mtime [3] ), .B1(_03138_ ), .B2(\CLINT.mtime [2] ), .ZN(_03357_ ) );
NOR3_X1 _19782_ ( .A1(_03140_ ), .A2(fanout_net_13 ), .A3(_03357_ ), .ZN(_00190_ ) );
AOI21_X1 _19783_ ( .A(\CLINT.mtime [2] ), .B1(\CLINT.mtime [1] ), .B2(\CLINT.mtime [0] ), .ZN(_03358_ ) );
NOR3_X1 _19784_ ( .A1(_03139_ ), .A2(fanout_net_13 ), .A3(_03358_ ), .ZN(_00191_ ) );
NOR2_X1 _19785_ ( .A1(\CLINT.mtime [1] ), .A2(\CLINT.mtime [0] ), .ZN(_03359_ ) );
NOR3_X1 _19786_ ( .A1(_03138_ ), .A2(_03359_ ), .A3(fanout_net_13 ), .ZN(_00192_ ) );
AND2_X1 _19787_ ( .A1(\CLINT.c_axi_arready_$_DFF_P__Q_D ), .A2(\CLINT.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_00193_ ) );
OR4_X1 _19788_ ( .A1(\CLINT.mtime [56] ), .A2(_03185_ ), .A3(_03173_ ), .A4(_03172_ ), .ZN(_03360_ ) );
NAND2_X1 _19789_ ( .A1(_03176_ ), .A2(\CLINT.mtime [56] ), .ZN(_03361_ ) );
AOI21_X1 _19790_ ( .A(fanout_net_13 ), .B1(_03360_ ), .B2(_03361_ ), .ZN(_00194_ ) );
NOR2_X1 _19791_ ( .A1(_03185_ ), .A2(_03172_ ), .ZN(_03362_ ) );
NAND3_X1 _19792_ ( .A1(_03362_ ), .A2(\CLINT.mtime [54] ), .A3(_03245_ ), .ZN(_03363_ ) );
OR2_X1 _19793_ ( .A1(_03363_ ), .A2(\CLINT.mtime [55] ), .ZN(_03364_ ) );
NAND2_X1 _19794_ ( .A1(_03363_ ), .A2(\CLINT.mtime [55] ), .ZN(_03365_ ) );
AOI21_X1 _19795_ ( .A(fanout_net_13 ), .B1(_03364_ ), .B2(_03365_ ), .ZN(_00195_ ) );
NAND2_X1 _19796_ ( .A1(_03362_ ), .A2(_03245_ ), .ZN(_03366_ ) );
OR2_X1 _19797_ ( .A1(_03366_ ), .A2(\CLINT.mtime [54] ), .ZN(_03367_ ) );
NAND2_X1 _19798_ ( .A1(_03366_ ), .A2(\CLINT.mtime [54] ), .ZN(_03368_ ) );
AOI21_X1 _19799_ ( .A(fanout_net_13 ), .B1(_03367_ ), .B2(_03368_ ), .ZN(_00196_ ) );
AOI21_X1 _19800_ ( .A(_04367_ ), .B1(_04372_ ), .B2(_04365_ ), .ZN(_03369_ ) );
XNOR2_X1 _19801_ ( .A(_03369_ ), .B(\EXU.counter [1] ), .ZN(_03370_ ) );
NOR2_X1 _19802_ ( .A1(\IDU.updata ), .A2(_03370_ ), .ZN(_00197_ ) );
OAI21_X1 _19803_ ( .A(\EXU.counter_$_SDFFE_PP0N__Q_1_D [0] ), .B1(_04361_ ), .B2(_04364_ ), .ZN(_03371_ ) );
NAND3_X1 _19804_ ( .A1(_04372_ ), .A2(\EXU.counter [0] ), .A3(_04365_ ), .ZN(_03372_ ) );
AOI21_X1 _19805_ ( .A(\IDU.updata ), .B1(_03371_ ), .B2(_03372_ ), .ZN(_00198_ ) );
NAND3_X1 _19806_ ( .A1(_05253_ ), .A2(\EXU.gpr_wen_o ), .A3(_04397_ ), .ZN(_03373_ ) );
OR4_X1 _19807_ ( .A1(\EXU.rd_i [3] ), .A2(\EXU.rd_i [2] ), .A3(\EXU.rd_i [1] ), .A4(\EXU.rd_i [0] ), .ZN(_03374_ ) );
OAI211_X1 _19808_ ( .A(\EXU.state ), .B(_03374_ ), .C1(_04393_ ), .C2(\LSU.ls_read_done_$_OR__B_Y_$_ORNOT__A_Y_$_ANDNOT__A_Y_$_OR__A_1_B ), .ZN(_03375_ ) );
AOI21_X1 _19809_ ( .A(_04331_ ), .B1(_03373_ ), .B2(_03375_ ), .ZN(_00235_ ) );
MUX2_X1 _19810_ ( .A(_05511_ ), .B(_05253_ ), .S(\EXU.state ), .Z(_03376_ ) );
AND2_X1 _19811_ ( .A1(_03376_ ), .A2(_05252_ ), .ZN(_00240_ ) );
AND3_X1 _19812_ ( .A1(_07887_ ), .A2(_07888_ ), .A3(_07890_ ), .ZN(_03377_ ) );
AND2_X1 _19813_ ( .A1(_07880_ ), .A2(_07660_ ), .ZN(_03378_ ) );
NOR3_X1 _19814_ ( .A1(_07622_ ), .A2(_07658_ ), .A3(_03378_ ), .ZN(_03379_ ) );
AND2_X1 _19815_ ( .A1(_03379_ ), .A2(\ICACHE.m_axi_arready ), .ZN(_03380_ ) );
INV_X1 _19816_ ( .A(_03380_ ), .ZN(_03381_ ) );
AOI21_X1 _19817_ ( .A(_03377_ ), .B1(_03381_ ), .B2(_07843_ ), .ZN(_03382_ ) );
MUX2_X1 _19818_ ( .A(_07690_ ), .B(_07889_ ), .S(_03382_ ), .Z(_03383_ ) );
NOR2_X1 _19819_ ( .A1(_03383_ ), .A2(fanout_net_13 ), .ZN(_00550_ ) );
AND2_X1 _19820_ ( .A1(_01589_ ), .A2(\ICACHE.m_axi_rready ), .ZN(_03384_ ) );
INV_X1 _19821_ ( .A(_03384_ ), .ZN(_03385_ ) );
INV_X1 _19822_ ( .A(_03379_ ), .ZN(_03386_ ) );
AOI22_X1 _19823_ ( .A1(_03385_ ), .A2(\ICACHE.s_axi_rready ), .B1(_07844_ ), .B2(_03386_ ), .ZN(_03387_ ) );
NOR2_X1 _19824_ ( .A1(_03387_ ), .A2(fanout_net_13 ), .ZN(_00551_ ) );
OAI21_X1 _19825_ ( .A(\IDU.state ), .B1(_05509_ ), .B2(\EXU.state ), .ZN(_03388_ ) );
AOI21_X1 _19826_ ( .A(_05086_ ), .B1(_02306_ ), .B2(_03388_ ), .ZN(_00739_ ) );
INV_X1 _19827_ ( .A(_04331_ ), .ZN(_03389_ ) );
AND3_X1 _19828_ ( .A1(_01582_ ), .A2(\ICACHE.m_axi_arvalid ), .A3(\ICACHE.s_axi_rready ), .ZN(_03390_ ) );
OAI211_X1 _19829_ ( .A(_03389_ ), .B(_03806_ ), .C1(\IFU.state_$_NOT__A_Y ), .C2(_03390_ ), .ZN(_03391_ ) );
INV_X1 _19830_ ( .A(_03391_ ), .ZN(_00740_ ) );
AND3_X1 _19831_ ( .A1(_01589_ ), .A2(\ICACHE.m_axi_rready ), .A3(\IFU.state ), .ZN(_03392_ ) );
OR2_X1 _19832_ ( .A1(_07660_ ), .A2(\IFU.state_$_NOT__A_Y ), .ZN(_03393_ ) );
AOI21_X1 _19833_ ( .A(\ICACHE.m_axi_rready ), .B1(_03393_ ), .B2(\IFU.state ), .ZN(_03394_ ) );
OR2_X1 _19834_ ( .A1(_03392_ ), .A2(_03394_ ), .ZN(_03395_ ) );
AOI21_X1 _19835_ ( .A(fanout_net_13 ), .B1(_03395_ ), .B2(_03389_ ), .ZN(_00741_ ) );
AOI21_X1 _19836_ ( .A(_05086_ ), .B1(\IFU.updata ), .B2(\IFU.state ), .ZN(_00836_ ) );
NOR2_X1 _19837_ ( .A1(_02642_ ), .A2(_02643_ ), .ZN(_03396_ ) );
OAI21_X1 _19838_ ( .A(_02508_ ), .B1(_03396_ ), .B2(_02498_ ), .ZN(_03397_ ) );
MUX2_X1 _19839_ ( .A(_02503_ ), .B(_02643_ ), .S(_03397_ ), .Z(_03398_ ) );
NOR2_X1 _19840_ ( .A1(_03398_ ), .A2(fanout_net_13 ), .ZN(_00869_ ) );
MUX2_X1 _19841_ ( .A(\LSU.axi_state [0] ), .B(_02639_ ), .S(\LSU.axi_state [1] ), .Z(_03399_ ) );
OAI21_X1 _19842_ ( .A(_03399_ ), .B1(_02553_ ), .B2(_02554_ ), .ZN(_03400_ ) );
MUX2_X1 _19843_ ( .A(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ), .B(\LSU.ls_axi_awvalid ), .S(_03400_ ), .Z(_03401_ ) );
AND2_X1 _19844_ ( .A1(_03401_ ), .A2(_03806_ ), .ZN(_00902_ ) );
NAND2_X1 _19845_ ( .A1(_04402_ ), .A2(\EXU.mcause_i [31] ), .ZN(_03402_ ) );
NAND2_X1 _19846_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [31] ), .ZN(_03403_ ) );
AOI21_X1 _19847_ ( .A(fanout_net_13 ), .B1(_03402_ ), .B2(_03403_ ), .ZN(_01451_ ) );
NAND2_X1 _19848_ ( .A1(_04402_ ), .A2(\EXU.mcause_i [30] ), .ZN(_03404_ ) );
NAND2_X1 _19849_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [30] ), .ZN(_03405_ ) );
AOI21_X1 _19850_ ( .A(fanout_net_13 ), .B1(_03404_ ), .B2(_03405_ ), .ZN(_01452_ ) );
NAND2_X1 _19851_ ( .A1(_04402_ ), .A2(\EXU.mcause_i [21] ), .ZN(_03406_ ) );
NAND2_X1 _19852_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [21] ), .ZN(_03407_ ) );
AOI21_X1 _19853_ ( .A(fanout_net_13 ), .B1(_03406_ ), .B2(_03407_ ), .ZN(_01453_ ) );
NAND2_X1 _19854_ ( .A1(_04402_ ), .A2(\EXU.mcause_i [20] ), .ZN(_03408_ ) );
NAND2_X1 _19855_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [20] ), .ZN(_03409_ ) );
AOI21_X1 _19856_ ( .A(fanout_net_13 ), .B1(_03408_ ), .B2(_03409_ ), .ZN(_01454_ ) );
NAND2_X1 _19857_ ( .A1(_04402_ ), .A2(\EXU.mcause_i [19] ), .ZN(_03410_ ) );
NAND2_X1 _19858_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [19] ), .ZN(_03411_ ) );
AOI21_X1 _19859_ ( .A(fanout_net_13 ), .B1(_03410_ ), .B2(_03411_ ), .ZN(_01455_ ) );
NAND2_X1 _19860_ ( .A1(_04402_ ), .A2(\EXU.mcause_i [18] ), .ZN(_03412_ ) );
NAND2_X1 _19861_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [18] ), .ZN(_03413_ ) );
AOI21_X1 _19862_ ( .A(fanout_net_13 ), .B1(_03412_ ), .B2(_03413_ ), .ZN(_01456_ ) );
NAND2_X1 _19863_ ( .A1(_04402_ ), .A2(\EXU.mcause_i [17] ), .ZN(_03414_ ) );
NAND2_X1 _19864_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [17] ), .ZN(_03415_ ) );
AOI21_X1 _19865_ ( .A(fanout_net_13 ), .B1(_03414_ ), .B2(_03415_ ), .ZN(_01457_ ) );
NAND2_X1 _19866_ ( .A1(_04402_ ), .A2(\EXU.mcause_i [16] ), .ZN(_03416_ ) );
NAND2_X1 _19867_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [16] ), .ZN(_03417_ ) );
AOI21_X1 _19868_ ( .A(fanout_net_13 ), .B1(_03416_ ), .B2(_03417_ ), .ZN(_01458_ ) );
NAND2_X1 _19869_ ( .A1(_04402_ ), .A2(\EXU.mcause_i [15] ), .ZN(_03418_ ) );
NAND2_X1 _19870_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [15] ), .ZN(_03419_ ) );
AOI21_X1 _19871_ ( .A(fanout_net_13 ), .B1(_03418_ ), .B2(_03419_ ), .ZN(_01459_ ) );
BUF_X4 _19872_ ( .A(_04401_ ), .Z(_03420_ ) );
NAND2_X1 _19873_ ( .A1(_03420_ ), .A2(\EXU.mcause_i [14] ), .ZN(_03421_ ) );
NAND2_X1 _19874_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [14] ), .ZN(_03422_ ) );
AOI21_X1 _19875_ ( .A(fanout_net_13 ), .B1(_03421_ ), .B2(_03422_ ), .ZN(_01460_ ) );
NAND2_X1 _19876_ ( .A1(_03420_ ), .A2(\EXU.mcause_i [13] ), .ZN(_03423_ ) );
NAND2_X1 _19877_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [13] ), .ZN(_03424_ ) );
AOI21_X1 _19878_ ( .A(fanout_net_13 ), .B1(_03423_ ), .B2(_03424_ ), .ZN(_01461_ ) );
NAND2_X1 _19879_ ( .A1(_03420_ ), .A2(\EXU.mcause_i [12] ), .ZN(_03425_ ) );
NAND2_X1 _19880_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [12] ), .ZN(_03426_ ) );
AOI21_X1 _19881_ ( .A(fanout_net_13 ), .B1(_03425_ ), .B2(_03426_ ), .ZN(_01462_ ) );
NAND2_X1 _19882_ ( .A1(_03420_ ), .A2(\EXU.mcause_i [29] ), .ZN(_03427_ ) );
NAND2_X1 _19883_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [29] ), .ZN(_03428_ ) );
AOI21_X1 _19884_ ( .A(fanout_net_13 ), .B1(_03427_ ), .B2(_03428_ ), .ZN(_01463_ ) );
NAND2_X1 _19885_ ( .A1(_03420_ ), .A2(\EXU.mcause_i [11] ), .ZN(_03429_ ) );
NAND2_X1 _19886_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [11] ), .ZN(_03430_ ) );
AOI21_X1 _19887_ ( .A(fanout_net_13 ), .B1(_03429_ ), .B2(_03430_ ), .ZN(_01464_ ) );
NAND2_X1 _19888_ ( .A1(_03420_ ), .A2(\EXU.mcause_i [10] ), .ZN(_03431_ ) );
NAND2_X1 _19889_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [10] ), .ZN(_03432_ ) );
AOI21_X1 _19890_ ( .A(fanout_net_13 ), .B1(_03431_ ), .B2(_03432_ ), .ZN(_01465_ ) );
NAND2_X1 _19891_ ( .A1(_03420_ ), .A2(\EXU.mcause_i [9] ), .ZN(_03433_ ) );
NAND2_X1 _19892_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [9] ), .ZN(_03434_ ) );
AOI21_X1 _19893_ ( .A(fanout_net_13 ), .B1(_03433_ ), .B2(_03434_ ), .ZN(_01466_ ) );
NAND2_X1 _19894_ ( .A1(_03420_ ), .A2(\EXU.mcause_i [8] ), .ZN(_03435_ ) );
NAND2_X1 _19895_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [8] ), .ZN(_03436_ ) );
AOI21_X1 _19896_ ( .A(fanout_net_13 ), .B1(_03435_ ), .B2(_03436_ ), .ZN(_01467_ ) );
NAND2_X1 _19897_ ( .A1(_03420_ ), .A2(\EXU.mcause_i [7] ), .ZN(_03437_ ) );
NAND2_X1 _19898_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [7] ), .ZN(_03438_ ) );
AOI21_X1 _19899_ ( .A(fanout_net_13 ), .B1(_03437_ ), .B2(_03438_ ), .ZN(_01468_ ) );
NAND2_X1 _19900_ ( .A1(_03420_ ), .A2(\EXU.mcause_i [6] ), .ZN(_03439_ ) );
NAND2_X1 _19901_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [6] ), .ZN(_03440_ ) );
AOI21_X1 _19902_ ( .A(fanout_net_14 ), .B1(_03439_ ), .B2(_03440_ ), .ZN(_01469_ ) );
BUF_X4 _19903_ ( .A(_04401_ ), .Z(_03441_ ) );
NAND2_X1 _19904_ ( .A1(_03441_ ), .A2(\EXU.mcause_i [5] ), .ZN(_03442_ ) );
NAND2_X1 _19905_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [5] ), .ZN(_03443_ ) );
AOI21_X1 _19906_ ( .A(fanout_net_14 ), .B1(_03442_ ), .B2(_03443_ ), .ZN(_01470_ ) );
NAND2_X1 _19907_ ( .A1(_03441_ ), .A2(\EXU.mcause_i [4] ), .ZN(_03444_ ) );
NAND2_X1 _19908_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [4] ), .ZN(_03445_ ) );
AOI21_X1 _19909_ ( .A(fanout_net_14 ), .B1(_03444_ ), .B2(_03445_ ), .ZN(_01471_ ) );
NAND2_X1 _19910_ ( .A1(_03441_ ), .A2(\EXU.mcause_i [3] ), .ZN(_03446_ ) );
NAND2_X1 _19911_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [3] ), .ZN(_03447_ ) );
AOI21_X1 _19912_ ( .A(fanout_net_14 ), .B1(_03446_ ), .B2(_03447_ ), .ZN(_01472_ ) );
NAND2_X1 _19913_ ( .A1(_03441_ ), .A2(\EXU.mcause_i [2] ), .ZN(_03448_ ) );
NAND2_X1 _19914_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [2] ), .ZN(_03449_ ) );
AOI21_X1 _19915_ ( .A(fanout_net_14 ), .B1(_03448_ ), .B2(_03449_ ), .ZN(_01473_ ) );
NAND2_X1 _19916_ ( .A1(_03441_ ), .A2(\EXU.mcause_i [28] ), .ZN(_03450_ ) );
NAND2_X1 _19917_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [28] ), .ZN(_03451_ ) );
AOI21_X1 _19918_ ( .A(fanout_net_14 ), .B1(_03450_ ), .B2(_03451_ ), .ZN(_01474_ ) );
NAND2_X1 _19919_ ( .A1(_03441_ ), .A2(\EXU.mcause_i [1] ), .ZN(_03452_ ) );
NAND2_X1 _19920_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [1] ), .ZN(_03453_ ) );
AOI21_X1 _19921_ ( .A(fanout_net_14 ), .B1(_03452_ ), .B2(_03453_ ), .ZN(_01475_ ) );
NAND2_X1 _19922_ ( .A1(_03441_ ), .A2(\EXU.mcause_i [0] ), .ZN(_03454_ ) );
NAND2_X1 _19923_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [0] ), .ZN(_03455_ ) );
AOI21_X1 _19924_ ( .A(fanout_net_14 ), .B1(_03454_ ), .B2(_03455_ ), .ZN(_01476_ ) );
NAND2_X1 _19925_ ( .A1(_03441_ ), .A2(\EXU.mcause_i [27] ), .ZN(_03456_ ) );
NAND2_X1 _19926_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [27] ), .ZN(_03457_ ) );
AOI21_X1 _19927_ ( .A(fanout_net_14 ), .B1(_03456_ ), .B2(_03457_ ), .ZN(_01477_ ) );
NAND2_X1 _19928_ ( .A1(_03441_ ), .A2(\EXU.mcause_i [26] ), .ZN(_03458_ ) );
NAND2_X1 _19929_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [26] ), .ZN(_03459_ ) );
AOI21_X1 _19930_ ( .A(fanout_net_14 ), .B1(_03458_ ), .B2(_03459_ ), .ZN(_01478_ ) );
NAND2_X1 _19931_ ( .A1(_03441_ ), .A2(\EXU.mcause_i [25] ), .ZN(_03460_ ) );
NAND2_X1 _19932_ ( .A1(fanout_net_3 ), .A2(\EXU.xrd_o [25] ), .ZN(_03461_ ) );
AOI21_X1 _19933_ ( .A(fanout_net_14 ), .B1(_03460_ ), .B2(_03461_ ), .ZN(_01479_ ) );
NAND2_X1 _19934_ ( .A1(_04401_ ), .A2(\EXU.mcause_i [24] ), .ZN(_03462_ ) );
NAND2_X1 _19935_ ( .A1(\EXU.csrs_wen_o [2] ), .A2(\EXU.xrd_o [24] ), .ZN(_03463_ ) );
AOI21_X1 _19936_ ( .A(fanout_net_14 ), .B1(_03462_ ), .B2(_03463_ ), .ZN(_01480_ ) );
NAND2_X1 _19937_ ( .A1(_04401_ ), .A2(\EXU.mcause_i [23] ), .ZN(_03464_ ) );
NAND2_X1 _19938_ ( .A1(\EXU.csrs_wen_o [2] ), .A2(\EXU.xrd_o [23] ), .ZN(_03465_ ) );
AOI21_X1 _19939_ ( .A(fanout_net_14 ), .B1(_03464_ ), .B2(_03465_ ), .ZN(_01481_ ) );
NAND2_X1 _19940_ ( .A1(_04401_ ), .A2(\EXU.mcause_i [22] ), .ZN(_03466_ ) );
NAND2_X1 _19941_ ( .A1(\EXU.csrs_wen_o [2] ), .A2(\EXU.xrd_o [22] ), .ZN(_03467_ ) );
AOI21_X1 _19942_ ( .A(fanout_net_14 ), .B1(_03466_ ), .B2(_03467_ ), .ZN(_01482_ ) );
NAND2_X1 _19943_ ( .A1(_04412_ ), .A2(\EXU.mepc_i [31] ), .ZN(_03468_ ) );
NAND2_X1 _19944_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [31] ), .ZN(_03469_ ) );
AOI21_X1 _19945_ ( .A(fanout_net_14 ), .B1(_03468_ ), .B2(_03469_ ), .ZN(_01483_ ) );
NAND2_X1 _19946_ ( .A1(_04412_ ), .A2(\EXU.mepc_i [30] ), .ZN(_03470_ ) );
NAND2_X1 _19947_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [30] ), .ZN(_03471_ ) );
AOI21_X1 _19948_ ( .A(fanout_net_14 ), .B1(_03470_ ), .B2(_03471_ ), .ZN(_01484_ ) );
NAND2_X1 _19949_ ( .A1(_04412_ ), .A2(\EXU.mepc_i [21] ), .ZN(_03472_ ) );
NAND2_X1 _19950_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [21] ), .ZN(_03473_ ) );
AOI21_X1 _19951_ ( .A(fanout_net_14 ), .B1(_03472_ ), .B2(_03473_ ), .ZN(_01485_ ) );
NAND2_X1 _19952_ ( .A1(_04412_ ), .A2(\EXU.mepc_i [20] ), .ZN(_03474_ ) );
NAND2_X1 _19953_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [20] ), .ZN(_03475_ ) );
AOI21_X1 _19954_ ( .A(fanout_net_14 ), .B1(_03474_ ), .B2(_03475_ ), .ZN(_01486_ ) );
NAND2_X1 _19955_ ( .A1(_04412_ ), .A2(\EXU.mepc_i [19] ), .ZN(_03476_ ) );
NAND2_X1 _19956_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [19] ), .ZN(_03477_ ) );
AOI21_X1 _19957_ ( .A(fanout_net_14 ), .B1(_03476_ ), .B2(_03477_ ), .ZN(_01487_ ) );
NAND2_X1 _19958_ ( .A1(_04412_ ), .A2(\EXU.mepc_i [18] ), .ZN(_03478_ ) );
NAND2_X1 _19959_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [18] ), .ZN(_03479_ ) );
AOI21_X1 _19960_ ( .A(fanout_net_14 ), .B1(_03478_ ), .B2(_03479_ ), .ZN(_01488_ ) );
NAND2_X1 _19961_ ( .A1(_04412_ ), .A2(\EXU.mepc_i [17] ), .ZN(_03480_ ) );
NAND2_X1 _19962_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [17] ), .ZN(_03481_ ) );
AOI21_X1 _19963_ ( .A(fanout_net_14 ), .B1(_03480_ ), .B2(_03481_ ), .ZN(_01489_ ) );
NAND2_X1 _19964_ ( .A1(_04412_ ), .A2(\EXU.mepc_i [16] ), .ZN(_03482_ ) );
NAND2_X1 _19965_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [16] ), .ZN(_03483_ ) );
AOI21_X1 _19966_ ( .A(fanout_net_14 ), .B1(_03482_ ), .B2(_03483_ ), .ZN(_01490_ ) );
NAND2_X1 _19967_ ( .A1(_04412_ ), .A2(\EXU.mepc_i [15] ), .ZN(_03484_ ) );
NAND2_X1 _19968_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [15] ), .ZN(_03485_ ) );
AOI21_X1 _19969_ ( .A(fanout_net_14 ), .B1(_03484_ ), .B2(_03485_ ), .ZN(_01491_ ) );
BUF_X4 _19970_ ( .A(_04411_ ), .Z(_03486_ ) );
NAND2_X1 _19971_ ( .A1(_03486_ ), .A2(\EXU.mepc_i [14] ), .ZN(_03487_ ) );
NAND2_X1 _19972_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [14] ), .ZN(_03488_ ) );
AOI21_X1 _19973_ ( .A(fanout_net_14 ), .B1(_03487_ ), .B2(_03488_ ), .ZN(_01492_ ) );
NAND2_X1 _19974_ ( .A1(_03486_ ), .A2(\EXU.mepc_i [13] ), .ZN(_03489_ ) );
NAND2_X1 _19975_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [13] ), .ZN(_03490_ ) );
AOI21_X1 _19976_ ( .A(fanout_net_14 ), .B1(_03489_ ), .B2(_03490_ ), .ZN(_01493_ ) );
NAND2_X1 _19977_ ( .A1(_03486_ ), .A2(\EXU.mepc_i [12] ), .ZN(_03491_ ) );
NAND2_X1 _19978_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [12] ), .ZN(_03492_ ) );
AOI21_X1 _19979_ ( .A(fanout_net_14 ), .B1(_03491_ ), .B2(_03492_ ), .ZN(_01494_ ) );
NAND2_X1 _19980_ ( .A1(_03486_ ), .A2(\EXU.mepc_i [29] ), .ZN(_03493_ ) );
NAND2_X1 _19981_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [29] ), .ZN(_03494_ ) );
AOI21_X1 _19982_ ( .A(fanout_net_14 ), .B1(_03493_ ), .B2(_03494_ ), .ZN(_01495_ ) );
NAND2_X1 _19983_ ( .A1(_03486_ ), .A2(\EXU.mepc_i [11] ), .ZN(_03495_ ) );
NAND2_X1 _19984_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [11] ), .ZN(_03496_ ) );
AOI21_X1 _19985_ ( .A(fanout_net_14 ), .B1(_03495_ ), .B2(_03496_ ), .ZN(_01496_ ) );
NAND2_X1 _19986_ ( .A1(_03486_ ), .A2(\EXU.mepc_i [10] ), .ZN(_03497_ ) );
NAND2_X1 _19987_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [10] ), .ZN(_03498_ ) );
AOI21_X1 _19988_ ( .A(fanout_net_14 ), .B1(_03497_ ), .B2(_03498_ ), .ZN(_01497_ ) );
NAND2_X1 _19989_ ( .A1(_03486_ ), .A2(\EXU.mepc_i [9] ), .ZN(_03499_ ) );
NAND2_X1 _19990_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [9] ), .ZN(_03500_ ) );
AOI21_X1 _19991_ ( .A(fanout_net_14 ), .B1(_03499_ ), .B2(_03500_ ), .ZN(_01498_ ) );
NAND2_X1 _19992_ ( .A1(_03486_ ), .A2(\EXU.mepc_i [8] ), .ZN(_03501_ ) );
NAND2_X1 _19993_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [8] ), .ZN(_03502_ ) );
AOI21_X1 _19994_ ( .A(fanout_net_15 ), .B1(_03501_ ), .B2(_03502_ ), .ZN(_01499_ ) );
NAND2_X1 _19995_ ( .A1(_03486_ ), .A2(\EXU.mepc_i [7] ), .ZN(_03503_ ) );
NAND2_X1 _19996_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [7] ), .ZN(_03504_ ) );
AOI21_X1 _19997_ ( .A(fanout_net_15 ), .B1(_03503_ ), .B2(_03504_ ), .ZN(_01500_ ) );
NAND2_X1 _19998_ ( .A1(_03486_ ), .A2(\EXU.mepc_i [6] ), .ZN(_03505_ ) );
NAND2_X1 _19999_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [6] ), .ZN(_03506_ ) );
AOI21_X1 _20000_ ( .A(fanout_net_15 ), .B1(_03505_ ), .B2(_03506_ ), .ZN(_01501_ ) );
BUF_X4 _20001_ ( .A(_04411_ ), .Z(_03507_ ) );
NAND2_X1 _20002_ ( .A1(_03507_ ), .A2(\EXU.mepc_i [5] ), .ZN(_03508_ ) );
NAND2_X1 _20003_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [5] ), .ZN(_03509_ ) );
AOI21_X1 _20004_ ( .A(fanout_net_15 ), .B1(_03508_ ), .B2(_03509_ ), .ZN(_01502_ ) );
NAND2_X1 _20005_ ( .A1(_03507_ ), .A2(\EXU.mepc_i [4] ), .ZN(_03510_ ) );
NAND2_X1 _20006_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [4] ), .ZN(_03511_ ) );
AOI21_X1 _20007_ ( .A(fanout_net_15 ), .B1(_03510_ ), .B2(_03511_ ), .ZN(_01503_ ) );
NAND2_X1 _20008_ ( .A1(_03507_ ), .A2(\EXU.mepc_i [3] ), .ZN(_03512_ ) );
NAND2_X1 _20009_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [3] ), .ZN(_03513_ ) );
AOI21_X1 _20010_ ( .A(fanout_net_15 ), .B1(_03512_ ), .B2(_03513_ ), .ZN(_01504_ ) );
NAND2_X1 _20011_ ( .A1(_03507_ ), .A2(\EXU.mepc_i [2] ), .ZN(_03514_ ) );
NAND2_X1 _20012_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [2] ), .ZN(_03515_ ) );
AOI21_X1 _20013_ ( .A(fanout_net_15 ), .B1(_03514_ ), .B2(_03515_ ), .ZN(_01505_ ) );
NAND2_X1 _20014_ ( .A1(_03507_ ), .A2(\EXU.mepc_i [28] ), .ZN(_03516_ ) );
NAND2_X1 _20015_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [28] ), .ZN(_03517_ ) );
AOI21_X1 _20016_ ( .A(fanout_net_15 ), .B1(_03516_ ), .B2(_03517_ ), .ZN(_01506_ ) );
NAND2_X1 _20017_ ( .A1(_03507_ ), .A2(\EXU.mepc_i [1] ), .ZN(_03518_ ) );
NAND2_X1 _20018_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [1] ), .ZN(_03519_ ) );
AOI21_X1 _20019_ ( .A(fanout_net_15 ), .B1(_03518_ ), .B2(_03519_ ), .ZN(_01507_ ) );
NAND2_X1 _20020_ ( .A1(_03507_ ), .A2(\EXU.mepc_i [0] ), .ZN(_03520_ ) );
NAND2_X1 _20021_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [0] ), .ZN(_03521_ ) );
AOI21_X1 _20022_ ( .A(fanout_net_15 ), .B1(_03520_ ), .B2(_03521_ ), .ZN(_01508_ ) );
NAND2_X1 _20023_ ( .A1(_03507_ ), .A2(\EXU.mepc_i [27] ), .ZN(_03522_ ) );
NAND2_X1 _20024_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [27] ), .ZN(_03523_ ) );
AOI21_X1 _20025_ ( .A(fanout_net_15 ), .B1(_03522_ ), .B2(_03523_ ), .ZN(_01509_ ) );
NAND2_X1 _20026_ ( .A1(_03507_ ), .A2(\EXU.mepc_i [26] ), .ZN(_03524_ ) );
NAND2_X1 _20027_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [26] ), .ZN(_03525_ ) );
AOI21_X1 _20028_ ( .A(fanout_net_15 ), .B1(_03524_ ), .B2(_03525_ ), .ZN(_01510_ ) );
NAND2_X1 _20029_ ( .A1(_03507_ ), .A2(\EXU.mepc_i [25] ), .ZN(_03526_ ) );
NAND2_X1 _20030_ ( .A1(fanout_net_1 ), .A2(\EXU.xrd_o [25] ), .ZN(_03527_ ) );
AOI21_X1 _20031_ ( .A(fanout_net_15 ), .B1(_03526_ ), .B2(_03527_ ), .ZN(_01511_ ) );
NAND2_X1 _20032_ ( .A1(_04411_ ), .A2(\EXU.mepc_i [24] ), .ZN(_03528_ ) );
NAND2_X1 _20033_ ( .A1(\EXU.csrs_wen_o [0] ), .A2(\EXU.xrd_o [24] ), .ZN(_03529_ ) );
AOI21_X1 _20034_ ( .A(fanout_net_15 ), .B1(_03528_ ), .B2(_03529_ ), .ZN(_01512_ ) );
NAND2_X1 _20035_ ( .A1(_04411_ ), .A2(\EXU.mepc_i [23] ), .ZN(_03530_ ) );
NAND2_X1 _20036_ ( .A1(\EXU.csrs_wen_o [0] ), .A2(\EXU.xrd_o [23] ), .ZN(_03531_ ) );
AOI21_X1 _20037_ ( .A(fanout_net_15 ), .B1(_03530_ ), .B2(_03531_ ), .ZN(_01513_ ) );
NAND2_X1 _20038_ ( .A1(_04411_ ), .A2(\EXU.mepc_i [22] ), .ZN(_03532_ ) );
NAND2_X1 _20039_ ( .A1(\EXU.csrs_wen_o [0] ), .A2(\EXU.xrd_o [22] ), .ZN(_03533_ ) );
AOI21_X1 _20040_ ( .A(fanout_net_15 ), .B1(_03532_ ), .B2(_03533_ ), .ZN(_01514_ ) );
NAND2_X1 _20041_ ( .A1(_04409_ ), .A2(\EXU.mstatus_i [31] ), .ZN(_03534_ ) );
NAND2_X1 _20042_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [31] ), .ZN(_03535_ ) );
AOI21_X1 _20043_ ( .A(fanout_net_15 ), .B1(_03534_ ), .B2(_03535_ ), .ZN(_01515_ ) );
NAND2_X1 _20044_ ( .A1(_04409_ ), .A2(\EXU.mstatus_i [30] ), .ZN(_03536_ ) );
NAND2_X1 _20045_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [30] ), .ZN(_03537_ ) );
AOI21_X1 _20046_ ( .A(fanout_net_15 ), .B1(_03536_ ), .B2(_03537_ ), .ZN(_01516_ ) );
NAND2_X1 _20047_ ( .A1(_04409_ ), .A2(\EXU.mstatus_i [21] ), .ZN(_03538_ ) );
NAND2_X1 _20048_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [21] ), .ZN(_03539_ ) );
AOI21_X1 _20049_ ( .A(fanout_net_15 ), .B1(_03538_ ), .B2(_03539_ ), .ZN(_01517_ ) );
NAND2_X1 _20050_ ( .A1(_04409_ ), .A2(\EXU.mstatus_i [20] ), .ZN(_03540_ ) );
NAND2_X1 _20051_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [20] ), .ZN(_03541_ ) );
AOI21_X1 _20052_ ( .A(fanout_net_15 ), .B1(_03540_ ), .B2(_03541_ ), .ZN(_01518_ ) );
NAND2_X1 _20053_ ( .A1(_04409_ ), .A2(\EXU.mstatus_i [19] ), .ZN(_03542_ ) );
NAND2_X1 _20054_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [19] ), .ZN(_03543_ ) );
AOI21_X1 _20055_ ( .A(fanout_net_15 ), .B1(_03542_ ), .B2(_03543_ ), .ZN(_01519_ ) );
NAND2_X1 _20056_ ( .A1(_04409_ ), .A2(\EXU.mstatus_i [18] ), .ZN(_03544_ ) );
NAND2_X1 _20057_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [18] ), .ZN(_03545_ ) );
AOI21_X1 _20058_ ( .A(fanout_net_15 ), .B1(_03544_ ), .B2(_03545_ ), .ZN(_01520_ ) );
NAND2_X1 _20059_ ( .A1(_04409_ ), .A2(\EXU.mstatus_i [17] ), .ZN(_03546_ ) );
NAND2_X1 _20060_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [17] ), .ZN(_03547_ ) );
AOI21_X1 _20061_ ( .A(fanout_net_15 ), .B1(_03546_ ), .B2(_03547_ ), .ZN(_01521_ ) );
NAND2_X1 _20062_ ( .A1(_04409_ ), .A2(\EXU.mstatus_i [16] ), .ZN(_03548_ ) );
NAND2_X1 _20063_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [16] ), .ZN(_03549_ ) );
AOI21_X1 _20064_ ( .A(fanout_net_15 ), .B1(_03548_ ), .B2(_03549_ ), .ZN(_01522_ ) );
NAND2_X1 _20065_ ( .A1(_04409_ ), .A2(\EXU.mstatus_i [15] ), .ZN(_03550_ ) );
NAND2_X1 _20066_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [15] ), .ZN(_03551_ ) );
AOI21_X1 _20067_ ( .A(fanout_net_15 ), .B1(_03550_ ), .B2(_03551_ ), .ZN(_01523_ ) );
BUF_X4 _20068_ ( .A(_04408_ ), .Z(_03552_ ) );
NAND2_X1 _20069_ ( .A1(_03552_ ), .A2(\EXU.mstatus_i [14] ), .ZN(_03553_ ) );
NAND2_X1 _20070_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [14] ), .ZN(_03554_ ) );
AOI21_X1 _20071_ ( .A(fanout_net_15 ), .B1(_03553_ ), .B2(_03554_ ), .ZN(_01524_ ) );
NAND2_X1 _20072_ ( .A1(_03552_ ), .A2(\EXU.mstatus_i [13] ), .ZN(_03555_ ) );
NAND2_X1 _20073_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [13] ), .ZN(_03556_ ) );
AOI21_X1 _20074_ ( .A(fanout_net_15 ), .B1(_03555_ ), .B2(_03556_ ), .ZN(_01525_ ) );
NAND2_X1 _20075_ ( .A1(_03552_ ), .A2(\EXU.mstatus_i [10] ), .ZN(_03557_ ) );
NAND2_X1 _20076_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [10] ), .ZN(_03558_ ) );
AOI21_X1 _20077_ ( .A(fanout_net_15 ), .B1(_03557_ ), .B2(_03558_ ), .ZN(_01526_ ) );
NAND2_X1 _20078_ ( .A1(_03552_ ), .A2(\EXU.mstatus_i [29] ), .ZN(_03559_ ) );
NAND2_X1 _20079_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [29] ), .ZN(_03560_ ) );
AOI21_X1 _20080_ ( .A(fanout_net_15 ), .B1(_03559_ ), .B2(_03560_ ), .ZN(_01527_ ) );
NAND2_X1 _20081_ ( .A1(_03552_ ), .A2(\EXU.mstatus_i [9] ), .ZN(_03561_ ) );
NAND2_X1 _20082_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [9] ), .ZN(_03562_ ) );
AOI21_X1 _20083_ ( .A(fanout_net_15 ), .B1(_03561_ ), .B2(_03562_ ), .ZN(_01528_ ) );
NAND2_X1 _20084_ ( .A1(_03552_ ), .A2(\EXU.mstatus_i [8] ), .ZN(_03563_ ) );
NAND2_X1 _20085_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [8] ), .ZN(_03564_ ) );
AOI21_X1 _20086_ ( .A(fanout_net_16 ), .B1(_03563_ ), .B2(_03564_ ), .ZN(_01529_ ) );
NAND2_X1 _20087_ ( .A1(_03552_ ), .A2(\EXU.mstatus_i [7] ), .ZN(_03565_ ) );
NAND2_X1 _20088_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [7] ), .ZN(_03566_ ) );
AOI21_X1 _20089_ ( .A(fanout_net_16 ), .B1(_03565_ ), .B2(_03566_ ), .ZN(_01530_ ) );
NAND2_X1 _20090_ ( .A1(_03552_ ), .A2(\EXU.mstatus_i [6] ), .ZN(_03567_ ) );
NAND2_X1 _20091_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [6] ), .ZN(_03568_ ) );
AOI21_X1 _20092_ ( .A(fanout_net_16 ), .B1(_03567_ ), .B2(_03568_ ), .ZN(_01531_ ) );
NAND2_X1 _20093_ ( .A1(_03552_ ), .A2(\EXU.mstatus_i [5] ), .ZN(_03569_ ) );
NAND2_X1 _20094_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [5] ), .ZN(_03570_ ) );
AOI21_X1 _20095_ ( .A(fanout_net_16 ), .B1(_03569_ ), .B2(_03570_ ), .ZN(_01532_ ) );
NAND2_X1 _20096_ ( .A1(_03552_ ), .A2(\EXU.mstatus_i [4] ), .ZN(_03571_ ) );
NAND2_X1 _20097_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [4] ), .ZN(_03572_ ) );
AOI21_X1 _20098_ ( .A(fanout_net_16 ), .B1(_03571_ ), .B2(_03572_ ), .ZN(_01533_ ) );
BUF_X4 _20099_ ( .A(_04408_ ), .Z(_03573_ ) );
NAND2_X1 _20100_ ( .A1(_03573_ ), .A2(\EXU.mstatus_i [3] ), .ZN(_03574_ ) );
NAND2_X1 _20101_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [3] ), .ZN(_03575_ ) );
AOI21_X1 _20102_ ( .A(fanout_net_16 ), .B1(_03574_ ), .B2(_03575_ ), .ZN(_01534_ ) );
NAND2_X1 _20103_ ( .A1(_03573_ ), .A2(\EXU.mstatus_i [2] ), .ZN(_03576_ ) );
NAND2_X1 _20104_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [2] ), .ZN(_03577_ ) );
AOI21_X1 _20105_ ( .A(fanout_net_16 ), .B1(_03576_ ), .B2(_03577_ ), .ZN(_01535_ ) );
NAND2_X1 _20106_ ( .A1(_03573_ ), .A2(\EXU.mstatus_i [1] ), .ZN(_03578_ ) );
NAND2_X1 _20107_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [1] ), .ZN(_03579_ ) );
AOI21_X1 _20108_ ( .A(fanout_net_16 ), .B1(_03578_ ), .B2(_03579_ ), .ZN(_01536_ ) );
NAND2_X1 _20109_ ( .A1(_03573_ ), .A2(\EXU.mstatus_i [0] ), .ZN(_03580_ ) );
NAND2_X1 _20110_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [0] ), .ZN(_03581_ ) );
AOI21_X1 _20111_ ( .A(fanout_net_16 ), .B1(_03580_ ), .B2(_03581_ ), .ZN(_01537_ ) );
NAND2_X1 _20112_ ( .A1(_03573_ ), .A2(\EXU.mstatus_i [28] ), .ZN(_03582_ ) );
NAND2_X1 _20113_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [28] ), .ZN(_03583_ ) );
AOI21_X1 _20114_ ( .A(fanout_net_16 ), .B1(_03582_ ), .B2(_03583_ ), .ZN(_01538_ ) );
NAND2_X1 _20115_ ( .A1(_03573_ ), .A2(\EXU.mstatus_i [27] ), .ZN(_03584_ ) );
NAND2_X1 _20116_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [27] ), .ZN(_03585_ ) );
AOI21_X1 _20117_ ( .A(fanout_net_16 ), .B1(_03584_ ), .B2(_03585_ ), .ZN(_01539_ ) );
NAND2_X1 _20118_ ( .A1(_03573_ ), .A2(\EXU.mstatus_i [26] ), .ZN(_03586_ ) );
NAND2_X1 _20119_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [26] ), .ZN(_03587_ ) );
AOI21_X1 _20120_ ( .A(fanout_net_16 ), .B1(_03586_ ), .B2(_03587_ ), .ZN(_01540_ ) );
NAND2_X1 _20121_ ( .A1(_03573_ ), .A2(\EXU.mstatus_i [25] ), .ZN(_03588_ ) );
NAND2_X1 _20122_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [25] ), .ZN(_03589_ ) );
AOI21_X1 _20123_ ( .A(fanout_net_16 ), .B1(_03588_ ), .B2(_03589_ ), .ZN(_01541_ ) );
NAND2_X1 _20124_ ( .A1(_03573_ ), .A2(\EXU.mstatus_i [24] ), .ZN(_03590_ ) );
NAND2_X1 _20125_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [24] ), .ZN(_03591_ ) );
AOI21_X1 _20126_ ( .A(fanout_net_16 ), .B1(_03590_ ), .B2(_03591_ ), .ZN(_01542_ ) );
NAND2_X1 _20127_ ( .A1(_03573_ ), .A2(\EXU.mstatus_i [23] ), .ZN(_03592_ ) );
NAND2_X1 _20128_ ( .A1(fanout_net_2 ), .A2(\EXU.xrd_o [23] ), .ZN(_03593_ ) );
AOI21_X1 _20129_ ( .A(fanout_net_16 ), .B1(_03592_ ), .B2(_03593_ ), .ZN(_01543_ ) );
NAND2_X1 _20130_ ( .A1(_04408_ ), .A2(\EXU.mstatus_i [22] ), .ZN(_03594_ ) );
NAND2_X1 _20131_ ( .A1(\EXU.csrs_wen_o [1] ), .A2(\EXU.xrd_o [22] ), .ZN(_03595_ ) );
AOI21_X1 _20132_ ( .A(fanout_net_16 ), .B1(_03594_ ), .B2(_03595_ ), .ZN(_01544_ ) );
NOR2_X1 _20133_ ( .A1(_04408_ ), .A2(\EXU.xrd_o [12] ), .ZN(_03596_ ) );
NOR2_X1 _20134_ ( .A1(\EXU.csrs_wen_o [1] ), .A2(\EXU.mstatus_i [12] ), .ZN(_03597_ ) );
OAI21_X1 _20135_ ( .A(\CLINT.c_axi_arready_$_DFF_P__Q_D ), .B1(_03596_ ), .B2(_03597_ ), .ZN(_01545_ ) );
NOR2_X1 _20136_ ( .A1(_04408_ ), .A2(\EXU.xrd_o [11] ), .ZN(_03598_ ) );
NOR2_X1 _20137_ ( .A1(\EXU.csrs_wen_o [1] ), .A2(\EXU.mstatus_i [11] ), .ZN(_03599_ ) );
OAI21_X1 _20138_ ( .A(\CLINT.c_axi_arready_$_DFF_P__Q_D ), .B1(_03598_ ), .B2(_03599_ ), .ZN(_01546_ ) );
NAND2_X1 _20139_ ( .A1(_04406_ ), .A2(\EXU.mtvec_i [31] ), .ZN(_03600_ ) );
NAND2_X1 _20140_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [31] ), .ZN(_03601_ ) );
AOI21_X1 _20141_ ( .A(fanout_net_16 ), .B1(_03600_ ), .B2(_03601_ ), .ZN(_01547_ ) );
NAND2_X1 _20142_ ( .A1(_04406_ ), .A2(\EXU.mtvec_i [30] ), .ZN(_03602_ ) );
NAND2_X1 _20143_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [30] ), .ZN(_03603_ ) );
AOI21_X1 _20144_ ( .A(fanout_net_16 ), .B1(_03602_ ), .B2(_03603_ ), .ZN(_01548_ ) );
NAND2_X1 _20145_ ( .A1(_04406_ ), .A2(\EXU.mtvec_i [21] ), .ZN(_03604_ ) );
NAND2_X1 _20146_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [21] ), .ZN(_03605_ ) );
AOI21_X1 _20147_ ( .A(fanout_net_16 ), .B1(_03604_ ), .B2(_03605_ ), .ZN(_01549_ ) );
NAND2_X1 _20148_ ( .A1(_04406_ ), .A2(\EXU.mtvec_i [20] ), .ZN(_03606_ ) );
NAND2_X1 _20149_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [20] ), .ZN(_03607_ ) );
AOI21_X1 _20150_ ( .A(fanout_net_16 ), .B1(_03606_ ), .B2(_03607_ ), .ZN(_01550_ ) );
NAND2_X1 _20151_ ( .A1(_04406_ ), .A2(\EXU.mtvec_i [19] ), .ZN(_03608_ ) );
NAND2_X1 _20152_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [19] ), .ZN(_03609_ ) );
AOI21_X1 _20153_ ( .A(fanout_net_16 ), .B1(_03608_ ), .B2(_03609_ ), .ZN(_01551_ ) );
NAND2_X1 _20154_ ( .A1(_04406_ ), .A2(\EXU.mtvec_i [18] ), .ZN(_03610_ ) );
NAND2_X1 _20155_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [18] ), .ZN(_03611_ ) );
AOI21_X1 _20156_ ( .A(fanout_net_16 ), .B1(_03610_ ), .B2(_03611_ ), .ZN(_01552_ ) );
NAND2_X1 _20157_ ( .A1(_04406_ ), .A2(\EXU.mtvec_i [17] ), .ZN(_03612_ ) );
NAND2_X1 _20158_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [17] ), .ZN(_03613_ ) );
AOI21_X1 _20159_ ( .A(fanout_net_16 ), .B1(_03612_ ), .B2(_03613_ ), .ZN(_01553_ ) );
NAND2_X1 _20160_ ( .A1(_04406_ ), .A2(\EXU.mtvec_i [16] ), .ZN(_03614_ ) );
NAND2_X1 _20161_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [16] ), .ZN(_03615_ ) );
AOI21_X1 _20162_ ( .A(fanout_net_16 ), .B1(_03614_ ), .B2(_03615_ ), .ZN(_01554_ ) );
NAND2_X1 _20163_ ( .A1(_04406_ ), .A2(\EXU.mtvec_i [15] ), .ZN(_03616_ ) );
NAND2_X1 _20164_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [15] ), .ZN(_03617_ ) );
AOI21_X1 _20165_ ( .A(fanout_net_16 ), .B1(_03616_ ), .B2(_03617_ ), .ZN(_01555_ ) );
BUF_X4 _20166_ ( .A(_04405_ ), .Z(_03618_ ) );
NAND2_X1 _20167_ ( .A1(_03618_ ), .A2(\EXU.mtvec_i [14] ), .ZN(_03619_ ) );
NAND2_X1 _20168_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [14] ), .ZN(_03620_ ) );
AOI21_X1 _20169_ ( .A(fanout_net_16 ), .B1(_03619_ ), .B2(_03620_ ), .ZN(_01556_ ) );
NAND2_X1 _20170_ ( .A1(_03618_ ), .A2(\EXU.mtvec_i [13] ), .ZN(_03621_ ) );
NAND2_X1 _20171_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [13] ), .ZN(_03622_ ) );
AOI21_X1 _20172_ ( .A(fanout_net_16 ), .B1(_03621_ ), .B2(_03622_ ), .ZN(_01557_ ) );
NAND2_X1 _20173_ ( .A1(_03618_ ), .A2(\EXU.mtvec_i [12] ), .ZN(_03623_ ) );
NAND2_X1 _20174_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [12] ), .ZN(_03624_ ) );
AOI21_X1 _20175_ ( .A(fanout_net_16 ), .B1(_03623_ ), .B2(_03624_ ), .ZN(_01558_ ) );
NAND2_X1 _20176_ ( .A1(_03618_ ), .A2(\EXU.mtvec_i [29] ), .ZN(_03625_ ) );
NAND2_X1 _20177_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [29] ), .ZN(_03626_ ) );
AOI21_X1 _20178_ ( .A(fanout_net_16 ), .B1(_03625_ ), .B2(_03626_ ), .ZN(_01559_ ) );
NAND2_X1 _20179_ ( .A1(_03618_ ), .A2(\EXU.mtvec_i [11] ), .ZN(_03627_ ) );
NAND2_X1 _20180_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [11] ), .ZN(_03628_ ) );
AOI21_X1 _20181_ ( .A(fanout_net_16 ), .B1(_03627_ ), .B2(_03628_ ), .ZN(_01560_ ) );
NAND2_X1 _20182_ ( .A1(_03618_ ), .A2(\EXU.mtvec_i [10] ), .ZN(_03629_ ) );
NAND2_X1 _20183_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [10] ), .ZN(_03630_ ) );
AOI21_X1 _20184_ ( .A(reset ), .B1(_03629_ ), .B2(_03630_ ), .ZN(_01561_ ) );
NAND2_X1 _20185_ ( .A1(_03618_ ), .A2(\EXU.mtvec_i [9] ), .ZN(_03631_ ) );
NAND2_X1 _20186_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [9] ), .ZN(_03632_ ) );
AOI21_X1 _20187_ ( .A(reset ), .B1(_03631_ ), .B2(_03632_ ), .ZN(_01562_ ) );
NAND2_X1 _20188_ ( .A1(_03618_ ), .A2(\EXU.mtvec_i [8] ), .ZN(_03633_ ) );
NAND2_X1 _20189_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [8] ), .ZN(_03634_ ) );
AOI21_X1 _20190_ ( .A(reset ), .B1(_03633_ ), .B2(_03634_ ), .ZN(_01563_ ) );
NAND2_X1 _20191_ ( .A1(_03618_ ), .A2(\EXU.mtvec_i [7] ), .ZN(_03635_ ) );
NAND2_X1 _20192_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [7] ), .ZN(_03636_ ) );
AOI21_X1 _20193_ ( .A(reset ), .B1(_03635_ ), .B2(_03636_ ), .ZN(_01564_ ) );
NAND2_X1 _20194_ ( .A1(_03618_ ), .A2(\EXU.mtvec_i [6] ), .ZN(_03637_ ) );
NAND2_X1 _20195_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [6] ), .ZN(_03638_ ) );
AOI21_X1 _20196_ ( .A(reset ), .B1(_03637_ ), .B2(_03638_ ), .ZN(_01565_ ) );
BUF_X4 _20197_ ( .A(_04405_ ), .Z(_03639_ ) );
NAND2_X1 _20198_ ( .A1(_03639_ ), .A2(\EXU.mtvec_i [5] ), .ZN(_03640_ ) );
NAND2_X1 _20199_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [5] ), .ZN(_03641_ ) );
AOI21_X1 _20200_ ( .A(reset ), .B1(_03640_ ), .B2(_03641_ ), .ZN(_01566_ ) );
NAND2_X1 _20201_ ( .A1(_03639_ ), .A2(\EXU.mtvec_i [4] ), .ZN(_03642_ ) );
NAND2_X1 _20202_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [4] ), .ZN(_03643_ ) );
AOI21_X1 _20203_ ( .A(reset ), .B1(_03642_ ), .B2(_03643_ ), .ZN(_01567_ ) );
NAND2_X1 _20204_ ( .A1(_03639_ ), .A2(\EXU.mtvec_i [3] ), .ZN(_03644_ ) );
NAND2_X1 _20205_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [3] ), .ZN(_03645_ ) );
AOI21_X1 _20206_ ( .A(reset ), .B1(_03644_ ), .B2(_03645_ ), .ZN(_01568_ ) );
NAND2_X1 _20207_ ( .A1(_03639_ ), .A2(\EXU.mtvec_i [2] ), .ZN(_03646_ ) );
NAND2_X1 _20208_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [2] ), .ZN(_03647_ ) );
AOI21_X1 _20209_ ( .A(reset ), .B1(_03646_ ), .B2(_03647_ ), .ZN(_01569_ ) );
NAND2_X1 _20210_ ( .A1(_03639_ ), .A2(\EXU.mtvec_i [28] ), .ZN(_03648_ ) );
NAND2_X1 _20211_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [28] ), .ZN(_03649_ ) );
AOI21_X1 _20212_ ( .A(reset ), .B1(_03648_ ), .B2(_03649_ ), .ZN(_01570_ ) );
NAND2_X1 _20213_ ( .A1(_03639_ ), .A2(\EXU.mtvec_i [1] ), .ZN(_03650_ ) );
NAND2_X1 _20214_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [1] ), .ZN(_03651_ ) );
AOI21_X1 _20215_ ( .A(reset ), .B1(_03650_ ), .B2(_03651_ ), .ZN(_01571_ ) );
NAND2_X1 _20216_ ( .A1(_03639_ ), .A2(\EXU.mtvec_i [0] ), .ZN(_03652_ ) );
NAND2_X1 _20217_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [0] ), .ZN(_03653_ ) );
AOI21_X1 _20218_ ( .A(reset ), .B1(_03652_ ), .B2(_03653_ ), .ZN(_01572_ ) );
NAND2_X1 _20219_ ( .A1(_03639_ ), .A2(\EXU.mtvec_i [27] ), .ZN(_03654_ ) );
NAND2_X1 _20220_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [27] ), .ZN(_03655_ ) );
AOI21_X1 _20221_ ( .A(reset ), .B1(_03654_ ), .B2(_03655_ ), .ZN(_01573_ ) );
NAND2_X1 _20222_ ( .A1(_03639_ ), .A2(\EXU.mtvec_i [26] ), .ZN(_03656_ ) );
NAND2_X1 _20223_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [26] ), .ZN(_03657_ ) );
AOI21_X1 _20224_ ( .A(reset ), .B1(_03656_ ), .B2(_03657_ ), .ZN(_01574_ ) );
NAND2_X1 _20225_ ( .A1(_03639_ ), .A2(\EXU.mtvec_i [25] ), .ZN(_03658_ ) );
NAND2_X1 _20226_ ( .A1(fanout_net_4 ), .A2(\EXU.xrd_o [25] ), .ZN(_03659_ ) );
AOI21_X1 _20227_ ( .A(reset ), .B1(_03658_ ), .B2(_03659_ ), .ZN(_01575_ ) );
NAND2_X1 _20228_ ( .A1(_04405_ ), .A2(\EXU.mtvec_i [24] ), .ZN(_03660_ ) );
NAND2_X1 _20229_ ( .A1(\EXU.csrs_wen_o [3] ), .A2(\EXU.xrd_o [24] ), .ZN(_03661_ ) );
AOI21_X1 _20230_ ( .A(reset ), .B1(_03660_ ), .B2(_03661_ ), .ZN(_01576_ ) );
NAND2_X1 _20231_ ( .A1(_04405_ ), .A2(\EXU.mtvec_i [23] ), .ZN(_03662_ ) );
NAND2_X1 _20232_ ( .A1(\EXU.csrs_wen_o [3] ), .A2(\EXU.xrd_o [23] ), .ZN(_03663_ ) );
AOI21_X1 _20233_ ( .A(reset ), .B1(_03662_ ), .B2(_03663_ ), .ZN(_01577_ ) );
NAND2_X1 _20234_ ( .A1(_04405_ ), .A2(\EXU.mtvec_i [22] ), .ZN(_03664_ ) );
NAND2_X1 _20235_ ( .A1(\EXU.csrs_wen_o [3] ), .A2(\EXU.xrd_o [22] ), .ZN(_03665_ ) );
AOI21_X1 _20236_ ( .A(reset ), .B1(_03664_ ), .B2(_03665_ ), .ZN(_01578_ ) );
OR3_X1 _20237_ ( .A1(_07622_ ), .A2(_07843_ ), .A3(_07658_ ), .ZN(_03666_ ) );
OAI21_X1 _20238_ ( .A(_01588_ ), .B1(_03666_ ), .B2(_01587_ ), .ZN(\ICACHE.axi_rvalid ) );
NOR4_X1 _20239_ ( .A1(\io_master_araddr [29] ), .A2(\io_master_araddr [28] ), .A3(\io_master_araddr [27] ), .A4(\io_master_araddr [24] ), .ZN(_03667_ ) );
NOR2_X1 _20240_ ( .A1(\io_master_araddr [31] ), .A2(\io_master_araddr [30] ), .ZN(_03668_ ) );
AND3_X1 _20241_ ( .A1(_03667_ ), .A2(_03668_ ), .A3(_04086_ ), .ZN(_03669_ ) );
AND4_X1 _20242_ ( .A1(_04087_ ), .A2(_03669_ ), .A3(_04084_ ), .A4(_04085_ ), .ZN(_03670_ ) );
NOR2_X1 _20243_ ( .A1(\io_master_araddr [9] ), .A2(\io_master_araddr [8] ), .ZN(_03671_ ) );
NOR4_X1 _20244_ ( .A1(\io_master_araddr [11] ), .A2(\io_master_araddr [10] ), .A3(\io_master_araddr [13] ), .A4(\io_master_araddr [12] ), .ZN(_03672_ ) );
NOR4_X1 _20245_ ( .A1(\io_master_araddr [15] ), .A2(\io_master_araddr [14] ), .A3(\io_master_araddr [26] ), .A4(_04082_ ), .ZN(_03673_ ) );
AND4_X1 _20246_ ( .A1(_03671_ ), .A2(_03672_ ), .A3(_03673_ ), .A4(_04064_ ), .ZN(_03674_ ) );
NAND2_X1 _20247_ ( .A1(_03670_ ), .A2(_03674_ ), .ZN(_03675_ ) );
NAND3_X1 _20248_ ( .A1(_04065_ ), .A2(_04066_ ), .A3(_04071_ ), .ZN(_03676_ ) );
NOR2_X1 _20249_ ( .A1(_03675_ ), .A2(_03676_ ), .ZN(_03677_ ) );
NAND3_X1 _20250_ ( .A1(_04065_ ), .A2(_04066_ ), .A3(_04095_ ), .ZN(_03678_ ) );
NOR2_X1 _20251_ ( .A1(_03675_ ), .A2(_03678_ ), .ZN(_03679_ ) );
NOR2_X1 _20252_ ( .A1(_03677_ ), .A2(_03679_ ), .ZN(\io_master_arburst [0] ) );
NAND4_X1 _20253_ ( .A1(_02506_ ), .A2(_03806_ ), .A3(\LSU.axi_state [0] ), .A4(_04384_ ), .ZN(_03680_ ) );
OR3_X1 _20254_ ( .A1(_04380_ ), .A2(reset ), .A3(_02608_ ), .ZN(_03681_ ) );
NAND2_X1 _20255_ ( .A1(_03680_ ), .A2(_03681_ ), .ZN(\LSU.axi_state_$_DFF_P__Q_1_D ) );
NOR4_X1 _20256_ ( .A1(_07542_ ), .A2(reset ), .A3(_02498_ ), .A4(_02504_ ), .ZN(_03682_ ) );
NOR4_X1 _20257_ ( .A1(_02507_ ), .A2(_02553_ ), .A3(reset ), .A4(_02554_ ), .ZN(_03683_ ) );
OR4_X1 _20258_ ( .A1(reset ), .A2(_03682_ ), .A3(_02556_ ), .A4(_03683_ ), .ZN(\LSU.axi_state_$_DFF_P__Q_2_D ) );
OAI211_X1 _20259_ ( .A(_03806_ ), .B(\LSU.axi_state [2] ), .C1(_07542_ ), .C2(_02504_ ), .ZN(_03684_ ) );
NAND4_X1 _20260_ ( .A1(_02506_ ), .A2(_03809_ ), .A3(\LSU.axi_state [0] ), .A4(_02847_ ), .ZN(_03685_ ) );
NAND2_X1 _20261_ ( .A1(_03684_ ), .A2(_03685_ ), .ZN(\LSU.axi_state_$_DFF_P__Q_D ) );
NOR2_X1 _20262_ ( .A1(\LSU.ls_axi_arvalid ), .A2(\LSU.ls_axi_awvalid ), .ZN(_03686_ ) );
NAND4_X1 _20263_ ( .A1(_03686_ ), .A2(\ICACHE.s_axi_arvalid ), .A3(_03833_ ), .A4(\Xbar.state [0] ), .ZN(_03687_ ) );
INV_X1 _20264_ ( .A(io_master_rvalid ), .ZN(_03688_ ) );
OAI21_X1 _20265_ ( .A(\ICACHE.s_axi_araddr [31] ), .B1(\ICACHE.s_axi_araddr [30] ), .B2(\ICACHE.s_axi_araddr [29] ), .ZN(_03689_ ) );
AOI21_X1 _20266_ ( .A(_03689_ ), .B1(\ICACHE.s_axi_araddr [31] ), .B2(\ICACHE.s_axi_araddr [30] ), .ZN(_03690_ ) );
NOR4_X1 _20267_ ( .A1(_07706_ ), .A2(_03688_ ), .A3(_03133_ ), .A4(_03690_ ), .ZN(_03691_ ) );
AND2_X1 _20268_ ( .A1(_03690_ ), .A2(io_master_rlast ), .ZN(_03692_ ) );
OR2_X1 _20269_ ( .A1(_03691_ ), .A2(_03692_ ), .ZN(_03693_ ) );
NAND2_X1 _20270_ ( .A1(_03806_ ), .A2(\Xbar.state [1] ), .ZN(_03694_ ) );
OAI21_X1 _20271_ ( .A(_03687_ ), .B1(_03693_ ), .B2(_03694_ ), .ZN(\Xbar.state_$_DFF_P__Q_1_D ) );
NAND3_X1 _20272_ ( .A1(_03693_ ), .A2(_03809_ ), .A3(\Xbar.state [1] ), .ZN(_03695_ ) );
NAND4_X1 _20273_ ( .A1(_03686_ ), .A2(_07889_ ), .A3(_03844_ ), .A4(\Xbar.state [0] ), .ZN(_03696_ ) );
NOR2_X1 _20274_ ( .A1(\CLINT.c_axi_rvalid ), .A2(io_master_bvalid ), .ZN(_03697_ ) );
NAND2_X1 _20275_ ( .A1(_03697_ ), .A2(_03688_ ), .ZN(_03698_ ) );
NAND3_X1 _20276_ ( .A1(_03698_ ), .A2(_03833_ ), .A3(\Xbar.state [2] ), .ZN(_03699_ ) );
NAND4_X1 _20277_ ( .A1(_03695_ ), .A2(\CLINT.c_axi_arready_$_DFF_P__Q_D ), .A3(_03696_ ), .A4(_03699_ ), .ZN(\Xbar.state_$_DFF_P__Q_2_D ) );
NAND3_X1 _20278_ ( .A1(_03697_ ), .A2(\Xbar.state [2] ), .A3(_03688_ ), .ZN(_03700_ ) );
AOI21_X1 _20279_ ( .A(reset ), .B1(_03700_ ), .B2(_04054_ ), .ZN(\Xbar.state_$_DFF_P__Q_D ) );
NOR3_X1 _20280_ ( .A1(_04110_ ), .A2(_04113_ ), .A3(_04082_ ), .ZN(\io_master_araddr [25] ) );
NOR3_X1 _20281_ ( .A1(_04110_ ), .A2(_04113_ ), .A3(_04070_ ), .ZN(\io_master_araddr [2] ) );
NOR4_X1 _20282_ ( .A1(_04110_ ), .A2(_04113_ ), .A3(_07835_ ), .A4(\io_master_awburst [0] ), .ZN(\io_master_arlen [3] ) );
AND4_X1 _20283_ ( .A1(\ICACHE.s_axi_arlen [1] ), .A2(_04111_ ), .A3(_04114_ ), .A4(_07831_ ), .ZN(\io_master_arlen [1] ) );
NOR4_X1 _20284_ ( .A1(_04110_ ), .A2(_04113_ ), .A3(_01584_ ), .A4(\io_master_awburst [0] ), .ZN(\io_master_arlen [0] ) );
OAI221_X1 _20285_ ( .A(_02847_ ), .B1(_04710_ ), .B2(_05026_ ), .C1(_04715_ ), .C2(_04709_ ), .ZN(_03701_ ) );
AOI21_X1 _20286_ ( .A(_07831_ ), .B1(_03701_ ), .B2(\LSU.ls_axi_arvalid ), .ZN(_03702_ ) );
NOR3_X1 _20287_ ( .A1(_04110_ ), .A2(_04113_ ), .A3(_03702_ ), .ZN(\io_master_arsize [1] ) );
AOI211_X1 _20288_ ( .A(\EXU.funct3_i [1] ), .B(_04714_ ), .C1(\EXU.funct3_i [2] ), .C2(io_master_arsize_$_ANDNOT__Y_1_B_$_OR__Y_A_$_OR__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_AND__Y_B_$_OR__Y_B ), .ZN(_03703_ ) );
AND4_X1 _20289_ ( .A1(_04106_ ), .A2(_07540_ ), .A3(_02847_ ), .A4(_03703_ ), .ZN(\io_master_arsize [0] ) );
NOR3_X1 _20290_ ( .A1(_04110_ ), .A2(_04113_ ), .A3(_03135_ ), .ZN(io_master_arvalid ) );
BUF_X4 _20291_ ( .A(_07831_ ), .Z(_03704_ ) );
BUF_X4 _20292_ ( .A(_03704_ ), .Z(_03705_ ) );
NOR2_X1 _20293_ ( .A1(_03705_ ), .A2(_02562_ ), .ZN(\io_master_awaddr [31] ) );
NOR2_X1 _20294_ ( .A1(_03705_ ), .A2(_02565_ ), .ZN(\io_master_awaddr [30] ) );
NOR2_X1 _20295_ ( .A1(_03705_ ), .A2(_02567_ ), .ZN(\io_master_awaddr [21] ) );
NOR2_X1 _20296_ ( .A1(_03705_ ), .A2(_02569_ ), .ZN(\io_master_awaddr [20] ) );
NOR2_X1 _20297_ ( .A1(_03705_ ), .A2(_02571_ ), .ZN(\io_master_awaddr [19] ) );
NOR2_X1 _20298_ ( .A1(_03705_ ), .A2(_02573_ ), .ZN(\io_master_awaddr [18] ) );
NOR2_X1 _20299_ ( .A1(_03705_ ), .A2(_02575_ ), .ZN(\io_master_awaddr [17] ) );
NOR2_X1 _20300_ ( .A1(_03705_ ), .A2(_02577_ ), .ZN(\io_master_awaddr [16] ) );
NOR2_X1 _20301_ ( .A1(_03705_ ), .A2(_02580_ ), .ZN(\io_master_awaddr [15] ) );
NOR2_X1 _20302_ ( .A1(_03705_ ), .A2(_02583_ ), .ZN(\io_master_awaddr [14] ) );
BUF_X4 _20303_ ( .A(_03704_ ), .Z(_03706_ ) );
NOR2_X1 _20304_ ( .A1(_03706_ ), .A2(_02586_ ), .ZN(\io_master_awaddr [13] ) );
NOR2_X1 _20305_ ( .A1(_03706_ ), .A2(_02589_ ), .ZN(\io_master_awaddr [12] ) );
NOR2_X1 _20306_ ( .A1(_03706_ ), .A2(_02591_ ), .ZN(\io_master_awaddr [29] ) );
NOR2_X1 _20307_ ( .A1(_03706_ ), .A2(_02593_ ), .ZN(\io_master_awaddr [11] ) );
NOR2_X1 _20308_ ( .A1(_03706_ ), .A2(_02595_ ), .ZN(\io_master_awaddr [10] ) );
NOR2_X1 _20309_ ( .A1(_03706_ ), .A2(_02597_ ), .ZN(\io_master_awaddr [9] ) );
NOR2_X1 _20310_ ( .A1(_03706_ ), .A2(_02599_ ), .ZN(\io_master_awaddr [8] ) );
NOR2_X1 _20311_ ( .A1(_03706_ ), .A2(_02601_ ), .ZN(\io_master_awaddr [7] ) );
NOR2_X1 _20312_ ( .A1(_03706_ ), .A2(_02604_ ), .ZN(\io_master_awaddr [6] ) );
NOR2_X1 _20313_ ( .A1(_03706_ ), .A2(_02607_ ), .ZN(\io_master_awaddr [5] ) );
BUF_X4 _20314_ ( .A(_03704_ ), .Z(_03707_ ) );
NOR2_X1 _20315_ ( .A1(_03707_ ), .A2(_02610_ ), .ZN(\io_master_awaddr [4] ) );
NOR2_X1 _20316_ ( .A1(_03707_ ), .A2(_02613_ ), .ZN(\io_master_awaddr [3] ) );
NOR2_X1 _20317_ ( .A1(_03707_ ), .A2(_02615_ ), .ZN(\io_master_awaddr [2] ) );
NOR2_X1 _20318_ ( .A1(_03707_ ), .A2(_02617_ ), .ZN(\io_master_awaddr [28] ) );
NOR2_X1 _20319_ ( .A1(_03707_ ), .A2(_02621_ ), .ZN(\io_master_awaddr [1] ) );
NOR2_X1 _20320_ ( .A1(_03707_ ), .A2(_02624_ ), .ZN(\io_master_awaddr [0] ) );
NOR2_X1 _20321_ ( .A1(_03707_ ), .A2(_02626_ ), .ZN(\io_master_awaddr [27] ) );
NOR2_X1 _20322_ ( .A1(_03707_ ), .A2(_02628_ ), .ZN(\io_master_awaddr [26] ) );
NOR2_X1 _20323_ ( .A1(_03707_ ), .A2(_02630_ ), .ZN(\io_master_awaddr [25] ) );
NOR2_X1 _20324_ ( .A1(_03707_ ), .A2(_02632_ ), .ZN(\io_master_awaddr [24] ) );
BUF_X4 _20325_ ( .A(_03704_ ), .Z(_03708_ ) );
NOR2_X1 _20326_ ( .A1(_03708_ ), .A2(_02634_ ), .ZN(\io_master_awaddr [23] ) );
NOR2_X1 _20327_ ( .A1(_03708_ ), .A2(_02636_ ), .ZN(\io_master_awaddr [22] ) );
AND2_X1 _20328_ ( .A1(_04384_ ), .A2(_05528_ ), .ZN(_03709_ ) );
AND3_X1 _20329_ ( .A1(_04382_ ), .A2(_04383_ ), .A3(_02918_ ), .ZN(_03710_ ) );
NOR4_X1 _20330_ ( .A1(_03709_ ), .A2(\LSU.ls_axi_awvalid_$_NOT__A_Y ), .A3(_03704_ ), .A4(_03710_ ), .ZN(\io_master_awsize [1] ) );
AND3_X1 _20331_ ( .A1(io_master_awvalid ), .A2(_04384_ ), .A3(_05528_ ), .ZN(\io_master_awsize [0] ) );
NOR3_X1 _20332_ ( .A1(_04110_ ), .A2(_04113_ ), .A3(_03133_ ), .ZN(io_master_rready ) );
NOR2_X1 _20333_ ( .A1(_03708_ ), .A2(_02666_ ), .ZN(\io_master_wdata [31] ) );
NOR2_X1 _20334_ ( .A1(_03708_ ), .A2(_02671_ ), .ZN(\io_master_wdata [30] ) );
NOR2_X1 _20335_ ( .A1(_03708_ ), .A2(_02675_ ), .ZN(\io_master_wdata [21] ) );
NOR2_X1 _20336_ ( .A1(_03708_ ), .A2(_02680_ ), .ZN(\io_master_wdata [20] ) );
NOR2_X1 _20337_ ( .A1(_03708_ ), .A2(_02685_ ), .ZN(\io_master_wdata [19] ) );
NOR2_X1 _20338_ ( .A1(_03708_ ), .A2(_02689_ ), .ZN(\io_master_wdata [18] ) );
NOR2_X1 _20339_ ( .A1(_03708_ ), .A2(_02692_ ), .ZN(\io_master_wdata [17] ) );
NOR2_X1 _20340_ ( .A1(_03708_ ), .A2(_02696_ ), .ZN(\io_master_wdata [16] ) );
BUF_X4 _20341_ ( .A(_03704_ ), .Z(_03711_ ) );
NOR2_X1 _20342_ ( .A1(_03711_ ), .A2(_02700_ ), .ZN(\io_master_wdata [15] ) );
NOR2_X1 _20343_ ( .A1(_03711_ ), .A2(_02703_ ), .ZN(\io_master_wdata [14] ) );
NOR2_X1 _20344_ ( .A1(_03711_ ), .A2(_02707_ ), .ZN(\io_master_wdata [13] ) );
NOR2_X1 _20345_ ( .A1(_03711_ ), .A2(_02710_ ), .ZN(\io_master_wdata [12] ) );
NOR2_X1 _20346_ ( .A1(_03711_ ), .A2(_02714_ ), .ZN(\io_master_wdata [29] ) );
NOR2_X1 _20347_ ( .A1(_03711_ ), .A2(_02718_ ), .ZN(\io_master_wdata [11] ) );
NOR2_X1 _20348_ ( .A1(_03711_ ), .A2(_02721_ ), .ZN(\io_master_wdata [10] ) );
NOR2_X1 _20349_ ( .A1(_03711_ ), .A2(_02724_ ), .ZN(\io_master_wdata [9] ) );
NOR2_X1 _20350_ ( .A1(_03711_ ), .A2(_02727_ ), .ZN(\io_master_wdata [8] ) );
NOR2_X1 _20351_ ( .A1(_03711_ ), .A2(_02730_ ), .ZN(\io_master_wdata [7] ) );
BUF_X4 _20352_ ( .A(_07831_ ), .Z(_03712_ ) );
NOR2_X1 _20353_ ( .A1(_03712_ ), .A2(_02732_ ), .ZN(\io_master_wdata [6] ) );
NOR2_X1 _20354_ ( .A1(_03712_ ), .A2(_02734_ ), .ZN(\io_master_wdata [5] ) );
NOR2_X1 _20355_ ( .A1(_03712_ ), .A2(_02736_ ), .ZN(\io_master_wdata [4] ) );
NOR2_X1 _20356_ ( .A1(_03712_ ), .A2(_02738_ ), .ZN(\io_master_wdata [3] ) );
NOR2_X1 _20357_ ( .A1(_03712_ ), .A2(_02740_ ), .ZN(\io_master_wdata [2] ) );
NOR2_X1 _20358_ ( .A1(_03712_ ), .A2(_02745_ ), .ZN(\io_master_wdata [28] ) );
NOR2_X1 _20359_ ( .A1(_03712_ ), .A2(_02747_ ), .ZN(\io_master_wdata [1] ) );
NOR2_X1 _20360_ ( .A1(_03712_ ), .A2(_02749_ ), .ZN(\io_master_wdata [0] ) );
NOR2_X1 _20361_ ( .A1(_03712_ ), .A2(_02753_ ), .ZN(\io_master_wdata [27] ) );
NOR2_X1 _20362_ ( .A1(_03712_ ), .A2(_02758_ ), .ZN(\io_master_wdata [26] ) );
NOR2_X1 _20363_ ( .A1(_03704_ ), .A2(_02762_ ), .ZN(\io_master_wdata [25] ) );
NOR2_X1 _20364_ ( .A1(_03704_ ), .A2(_02767_ ), .ZN(\io_master_wdata [24] ) );
NOR2_X1 _20365_ ( .A1(_03704_ ), .A2(_02770_ ), .ZN(\io_master_wdata [23] ) );
NOR2_X1 _20366_ ( .A1(_03704_ ), .A2(_02773_ ), .ZN(\io_master_wdata [22] ) );
AND2_X1 _20367_ ( .A1(\io_master_awburst [0] ), .A2(\LSU.ls_axi_wlast ), .ZN(io_master_wlast ) );
INV_X1 _20368_ ( .A(io_master_wvalid ), .ZN(_03713_ ) );
AOI22_X1 _20369_ ( .A1(_02955_ ), .A2(_03710_ ), .B1(_02655_ ), .B2(_03709_ ), .ZN(_03714_ ) );
NOR3_X1 _20370_ ( .A1(_02649_ ), .A2(_04413_ ), .A3(_02650_ ), .ZN(_03715_ ) );
NAND2_X1 _20371_ ( .A1(_03715_ ), .A2(_02800_ ), .ZN(_03716_ ) );
AOI21_X1 _20372_ ( .A(_03713_ ), .B1(_03714_ ), .B2(_03716_ ), .ZN(\io_master_wstrb [3] ) );
OAI211_X1 _20373_ ( .A(_02649_ ), .B(_02623_ ), .C1(_03710_ ), .C2(_03709_ ), .ZN(_03717_ ) );
AOI21_X1 _20374_ ( .A(_03713_ ), .B1(_03716_ ), .B2(_03717_ ), .ZN(\io_master_wstrb [2] ) );
OAI21_X1 _20375_ ( .A(_03715_ ), .B1(_05528_ ), .B2(_02800_ ), .ZN(_03718_ ) );
NAND4_X1 _20376_ ( .A1(_05354_ ), .A2(_02552_ ), .A3(_05359_ ), .A4(_03710_ ), .ZN(_03719_ ) );
AOI21_X1 _20377_ ( .A(_03713_ ), .B1(_03718_ ), .B2(_03719_ ), .ZN(\io_master_wstrb [1] ) );
NAND4_X1 _20378_ ( .A1(_02619_ ), .A2(_04384_ ), .A3(_02918_ ), .A4(_02623_ ), .ZN(_03720_ ) );
AOI21_X1 _20379_ ( .A(_03713_ ), .B1(_03718_ ), .B2(_03720_ ), .ZN(\io_master_wstrb [0] ) );
LOGIC0_X1 _20380_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \BTB.bsnpc_reg[0]_$_SDFFCE_PN0P__Q ( .D(_00000_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[0][7] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_Y ) );
DFF_X1 \BTB.bsnpc_reg[0]_$_SDFFCE_PN0P__Q_1 ( .D(_00001_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[0][6] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_1_Y ) );
DFF_X1 \BTB.bsnpc_reg[0]_$_SDFFCE_PN0P__Q_2 ( .D(_00002_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[0][5] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_2_Y ) );
DFF_X1 \BTB.bsnpc_reg[0]_$_SDFFCE_PN0P__Q_3 ( .D(_00003_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[0][4] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_3_Y ) );
DFF_X1 \BTB.bsnpc_reg[0]_$_SDFFCE_PN0P__Q_4 ( .D(_00004_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[0][3] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_4_Y ) );
DFF_X1 \BTB.bsnpc_reg[0]_$_SDFFCE_PN0P__Q_5 ( .D(_00005_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[0][2] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_5_Y ) );
DFF_X1 \BTB.bsnpc_reg[0]_$_SDFFCE_PN0P__Q_6 ( .D(_00006_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[0][1] ), .QN(_10790_ ) );
DFF_X1 \BTB.bsnpc_reg[0]_$_SDFFCE_PN0P__Q_7 ( .D(_00007_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[0][0] ), .QN(_10789_ ) );
DFF_X1 \BTB.bsnpc_reg[1]_$_SDFFCE_PN0P__Q ( .D(_00008_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[1][7] ), .QN(\BTB.bsnpc_reg[1]_$_NOT__A_Y ) );
DFF_X1 \BTB.bsnpc_reg[1]_$_SDFFCE_PN0P__Q_1 ( .D(_00009_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[1][6] ), .QN(\BTB.bsnpc_reg[1]_$_NOT__A_1_Y ) );
DFF_X1 \BTB.bsnpc_reg[1]_$_SDFFCE_PN0P__Q_2 ( .D(_00010_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[1][5] ), .QN(\BTB.bsnpc_reg[1]_$_NOT__A_2_Y ) );
DFF_X1 \BTB.bsnpc_reg[1]_$_SDFFCE_PN0P__Q_3 ( .D(_00011_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[1][4] ), .QN(\BTB.bsnpc_reg[1]_$_NOT__A_3_Y ) );
DFF_X1 \BTB.bsnpc_reg[1]_$_SDFFCE_PN0P__Q_4 ( .D(_00012_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[1][3] ), .QN(\BTB.bsnpc_reg[1]_$_NOT__A_4_Y ) );
DFF_X1 \BTB.bsnpc_reg[1]_$_SDFFCE_PN0P__Q_5 ( .D(_00013_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[1][2] ), .QN(\BTB.bsnpc_reg[1]_$_NOT__A_5_Y ) );
DFF_X1 \BTB.bsnpc_reg[1]_$_SDFFCE_PN0P__Q_6 ( .D(_00014_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[1][1] ), .QN(_10788_ ) );
DFF_X1 \BTB.bsnpc_reg[1]_$_SDFFCE_PN0P__Q_7 ( .D(_00015_ ), .CK(clock ), .Q(\BTB.bsnpc_reg[1][0] ), .QN(_10787_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q ( .D(_00016_ ), .CK(clock ), .Q(\BTB.btag_reg[0][12] ), .QN(_10786_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q_1 ( .D(_00017_ ), .CK(clock ), .Q(\BTB.btag_reg[0][11] ), .QN(_10785_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q_10 ( .D(_00018_ ), .CK(clock ), .Q(\BTB.btag_reg[0][2] ), .QN(_10784_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q_11 ( .D(_00019_ ), .CK(clock ), .Q(\BTB.btag_reg[0][1] ), .QN(_10783_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q_12 ( .D(_00020_ ), .CK(clock ), .Q(\BTB.btag_reg[0][0] ), .QN(_10782_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q_2 ( .D(_00021_ ), .CK(clock ), .Q(\BTB.btag_reg[0][10] ), .QN(_10781_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q_3 ( .D(_00022_ ), .CK(clock ), .Q(\BTB.btag_reg[0][9] ), .QN(_10780_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q_4 ( .D(_00023_ ), .CK(clock ), .Q(\BTB.btag_reg[0][8] ), .QN(_10779_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q_5 ( .D(_00024_ ), .CK(clock ), .Q(\BTB.btag_reg[0][7] ), .QN(_10778_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q_6 ( .D(_00025_ ), .CK(clock ), .Q(\BTB.btag_reg[0][6] ), .QN(_10777_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q_7 ( .D(_00026_ ), .CK(clock ), .Q(\BTB.btag_reg[0][5] ), .QN(_10776_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q_8 ( .D(_00027_ ), .CK(clock ), .Q(\BTB.btag_reg[0][4] ), .QN(_10775_ ) );
DFF_X1 \BTB.btag_reg[0]_$_SDFFCE_PN0P__Q_9 ( .D(_00028_ ), .CK(clock ), .Q(\BTB.btag_reg[0][3] ), .QN(_10774_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q ( .D(_00029_ ), .CK(clock ), .Q(\BTB.btag_reg[1][12] ), .QN(_10773_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q_1 ( .D(_00030_ ), .CK(clock ), .Q(\BTB.btag_reg[1][11] ), .QN(_10772_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q_10 ( .D(_00031_ ), .CK(clock ), .Q(\BTB.btag_reg[1][2] ), .QN(_10771_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q_11 ( .D(_00032_ ), .CK(clock ), .Q(\BTB.btag_reg[1][1] ), .QN(_10770_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q_12 ( .D(_00033_ ), .CK(clock ), .Q(\BTB.btag_reg[1][0] ), .QN(_10769_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q_2 ( .D(_00034_ ), .CK(clock ), .Q(\BTB.btag_reg[1][10] ), .QN(_10768_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q_3 ( .D(_00035_ ), .CK(clock ), .Q(\BTB.btag_reg[1][9] ), .QN(_10767_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q_4 ( .D(_00036_ ), .CK(clock ), .Q(\BTB.btag_reg[1][8] ), .QN(_10766_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q_5 ( .D(_00037_ ), .CK(clock ), .Q(\BTB.btag_reg[1][7] ), .QN(_10765_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q_6 ( .D(_00038_ ), .CK(clock ), .Q(\BTB.btag_reg[1][6] ), .QN(_10764_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q_7 ( .D(_00039_ ), .CK(clock ), .Q(\BTB.btag_reg[1][5] ), .QN(_10763_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q_8 ( .D(_00040_ ), .CK(clock ), .Q(\BTB.btag_reg[1][4] ), .QN(_10762_ ) );
DFF_X1 \BTB.btag_reg[1]_$_SDFFCE_PN0P__Q_9 ( .D(_00041_ ), .CK(clock ), .Q(\BTB.btag_reg[1][3] ), .QN(_10761_ ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q ( .D(_00042_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][15] ), .QN(_10760_ ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_1 ( .D(_00043_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][14] ), .QN(_10759_ ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_10 ( .D(_00044_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][5] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_2_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_11 ( .D(_00045_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][4] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_3_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_12 ( .D(_00046_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][3] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_4_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_13 ( .D(_00047_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][2] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_5_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_14 ( .D(_00048_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][1] ), .QN(_10758_ ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_15 ( .D(_00049_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][0] ), .QN(_10757_ ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_2 ( .D(_00050_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][13] ), .QN(_10756_ ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_3 ( .D(_00051_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][12] ), .QN(_10755_ ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_4 ( .D(_00052_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][11] ), .QN(_10754_ ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_5 ( .D(_00053_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][10] ), .QN(_10753_ ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_6 ( .D(_00054_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][9] ), .QN(_10752_ ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_7 ( .D(_00055_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][8] ), .QN(_10751_ ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_8 ( .D(_00056_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][7] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ) );
DFF_X1 \BTB.jsnpc_reg[0]_$_SDFFCE_PN0P__Q_9 ( .D(_00057_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[0][6] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_1_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_A ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q ( .D(_00058_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][15] ), .QN(_10750_ ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_1 ( .D(_00059_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][14] ), .QN(_10749_ ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_10 ( .D(_00060_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][5] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_2_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_11 ( .D(_00061_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][4] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_3_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_12 ( .D(_00062_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][3] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_4_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_13 ( .D(_00063_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][2] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_5_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_14 ( .D(_00064_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][1] ), .QN(_10748_ ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_15 ( .D(_00065_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][0] ), .QN(_10747_ ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_2 ( .D(_00066_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][13] ), .QN(_10746_ ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_3 ( .D(_00067_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][12] ), .QN(_10745_ ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_4 ( .D(_00068_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][11] ), .QN(_10744_ ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_5 ( .D(_00069_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][10] ), .QN(_10743_ ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_6 ( .D(_00070_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][9] ), .QN(_10742_ ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_7 ( .D(_00071_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][8] ), .QN(_10741_ ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_8 ( .D(_00072_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][7] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \BTB.jsnpc_reg[1]_$_SDFFCE_PN0P__Q_9 ( .D(_00073_ ), .CK(clock ), .Q(\BTB.jsnpc_reg[1][6] ), .QN(\BTB.bsnpc_reg[0]_$_NOT__A_1_Y_$_MUX__A_Y_$_MUX__B_Y_$_MUX__A_B_$_MUX__Y_B ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q ( .D(_00074_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][12] ), .QN(_10740_ ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q_1 ( .D(_00075_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][11] ), .QN(_10739_ ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q_10 ( .D(_00076_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][2] ), .QN(_10738_ ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q_11 ( .D(_00077_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][1] ), .QN(_10737_ ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q_12 ( .D(_00078_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][0] ), .QN(_10736_ ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q_2 ( .D(_00079_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][10] ), .QN(_10735_ ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q_3 ( .D(_00080_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][9] ), .QN(_10734_ ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q_4 ( .D(_00081_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][8] ), .QN(_10733_ ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q_5 ( .D(_00082_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][7] ), .QN(_10732_ ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q_6 ( .D(_00083_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][6] ), .QN(_10731_ ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q_7 ( .D(_00084_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][5] ), .QN(_10730_ ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q_8 ( .D(_00085_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][4] ), .QN(_10729_ ) );
DFF_X1 \BTB.jtag_reg[0]_$_SDFFCE_PN0P__Q_9 ( .D(_00086_ ), .CK(clock ), .Q(\BTB.jtag_reg[0][3] ), .QN(_10728_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q ( .D(_00087_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][12] ), .QN(_10727_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q_1 ( .D(_00088_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][11] ), .QN(_10726_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q_10 ( .D(_00089_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][2] ), .QN(_10725_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q_11 ( .D(_00090_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][1] ), .QN(_10724_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q_12 ( .D(_00091_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][0] ), .QN(_10723_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q_2 ( .D(_00092_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][10] ), .QN(_10722_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q_3 ( .D(_00093_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][9] ), .QN(_10721_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q_4 ( .D(_00094_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][8] ), .QN(_10720_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q_5 ( .D(_00095_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][7] ), .QN(_10719_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q_6 ( .D(_00096_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][6] ), .QN(_10718_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q_7 ( .D(_00097_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][5] ), .QN(_10717_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q_8 ( .D(_00098_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][4] ), .QN(_10716_ ) );
DFF_X1 \BTB.jtag_reg[1]_$_SDFFCE_PN0P__Q_9 ( .D(_00099_ ), .CK(clock ), .Q(\BTB.jtag_reg[1][3] ), .QN(_10791_ ) );
DFF_X1 CHazarden_$_DFF_P__Q ( .D(\IDU.updata ), .CK(clock ), .Q(CHazarden ), .QN(_10792_ ) );
DFF_X1 \CLINT.c_axi_arready_$_DFF_P__Q ( .D(\CLINT.c_axi_arready_$_DFF_P__Q_D ), .CK(clock ), .Q(\CLINT.c_axi_arready ), .QN(\CLINT.c_axi_arready_$_NOT__A_Y ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q ( .D(_00100_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [31] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_1 ( .D(_00101_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [30] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_1_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_10 ( .D(_00102_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [21] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_10_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_11 ( .D(_00103_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [20] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_11_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_12 ( .D(_00104_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [19] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_12_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_13 ( .D(_00105_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [18] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_13_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_14 ( .D(_00106_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [17] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_14_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_15 ( .D(_00107_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [16] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_15_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_16 ( .D(_00108_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [15] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_16_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_17 ( .D(_00109_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [14] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_17_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_18 ( .D(_00110_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [13] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_18_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_19 ( .D(_00111_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [12] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_19_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_2 ( .D(_00112_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [29] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_2_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_20 ( .D(_00113_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [11] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_20_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_21 ( .D(_00114_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [10] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_21_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_22 ( .D(_00115_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [9] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_22_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_23 ( .D(_00116_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [8] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_23_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_24 ( .D(_00117_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [7] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_24_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_25 ( .D(_00118_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [6] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_25_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_26 ( .D(_00119_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [5] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_26_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_27 ( .D(_00120_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [4] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_27_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_28 ( .D(_00121_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [3] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_28_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_29 ( .D(_00122_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [2] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_29_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_3 ( .D(_00123_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [28] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_3_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_30 ( .D(_00124_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [1] ), .QN(_10715_ ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_31 ( .D(_00125_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [0] ), .QN(_10714_ ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_4 ( .D(_00126_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [27] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_4_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_5 ( .D(_00127_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [26] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_5_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_6 ( .D(_00128_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [25] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_6_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_7 ( .D(_00129_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [24] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_7_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_8 ( .D(_00130_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [23] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_8_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rdata_$_DFFE_PP__Q_9 ( .D(_00131_ ), .CK(clock ), .Q(\CLINT.c_axi_rdata [22] ), .QN(\ICACHE.s_axi_rdata_$_ANDNOT__Y_9_B_$_MUX__Y_A ) );
DFF_X1 \CLINT.c_axi_rvalid_$_SDFFE_PP0P__Q ( .D(_00132_ ), .CK(clock ), .Q(\CLINT.c_axi_rvalid ), .QN(\CLINT.c_axi_rvalid_$_NOT__A_Y ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q ( .D(_00133_ ), .CK(clock ), .Q(\CLINT.mtime [63] ), .QN(_10713_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_1 ( .D(_00134_ ), .CK(clock ), .Q(\CLINT.mtime [62] ), .QN(_10712_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_10 ( .D(_00135_ ), .CK(clock ), .Q(\CLINT.mtime [53] ), .QN(_10711_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_11 ( .D(_00136_ ), .CK(clock ), .Q(\CLINT.mtime [52] ), .QN(_10710_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_12 ( .D(_00137_ ), .CK(clock ), .Q(\CLINT.mtime [51] ), .QN(_10709_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_13 ( .D(_00138_ ), .CK(clock ), .Q(\CLINT.mtime [50] ), .QN(_10708_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_14 ( .D(_00139_ ), .CK(clock ), .Q(\CLINT.mtime [49] ), .QN(_10707_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_15 ( .D(_00140_ ), .CK(clock ), .Q(\CLINT.mtime [48] ), .QN(_10706_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_16 ( .D(_00141_ ), .CK(clock ), .Q(\CLINT.mtime [47] ), .QN(_10705_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_17 ( .D(_00142_ ), .CK(clock ), .Q(\CLINT.mtime [46] ), .QN(_10704_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_18 ( .D(_00143_ ), .CK(clock ), .Q(\CLINT.mtime [45] ), .QN(_10703_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_19 ( .D(_00144_ ), .CK(clock ), .Q(\CLINT.mtime [44] ), .QN(_10702_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_2 ( .D(_00145_ ), .CK(clock ), .Q(\CLINT.mtime [61] ), .QN(_10701_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_20 ( .D(_00146_ ), .CK(clock ), .Q(\CLINT.mtime [43] ), .QN(_10700_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_21 ( .D(_00147_ ), .CK(clock ), .Q(\CLINT.mtime [42] ), .QN(_10699_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_22 ( .D(_00148_ ), .CK(clock ), .Q(\CLINT.mtime [41] ), .QN(_10698_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_23 ( .D(_00149_ ), .CK(clock ), .Q(\CLINT.mtime [40] ), .QN(_10697_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_24 ( .D(_00150_ ), .CK(clock ), .Q(\CLINT.mtime [39] ), .QN(_10696_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_25 ( .D(_00151_ ), .CK(clock ), .Q(\CLINT.mtime [38] ), .QN(_10695_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_26 ( .D(_00152_ ), .CK(clock ), .Q(\CLINT.mtime [37] ), .QN(_10694_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_27 ( .D(_00153_ ), .CK(clock ), .Q(\CLINT.mtime [36] ), .QN(_10693_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_28 ( .D(_00154_ ), .CK(clock ), .Q(\CLINT.mtime [35] ), .QN(_10692_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_29 ( .D(_00155_ ), .CK(clock ), .Q(\CLINT.mtime [34] ), .QN(_10691_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_3 ( .D(_00156_ ), .CK(clock ), .Q(\CLINT.mtime [60] ), .QN(_10690_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_30 ( .D(_00157_ ), .CK(clock ), .Q(\CLINT.mtime [33] ), .QN(_10689_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_31 ( .D(_00158_ ), .CK(clock ), .Q(\CLINT.mtime [32] ), .QN(_10688_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_32 ( .D(_00159_ ), .CK(clock ), .Q(\CLINT.mtime [31] ), .QN(_10687_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_33 ( .D(_00160_ ), .CK(clock ), .Q(\CLINT.mtime [30] ), .QN(_10686_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_34 ( .D(_00161_ ), .CK(clock ), .Q(\CLINT.mtime [29] ), .QN(_10685_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_35 ( .D(_00162_ ), .CK(clock ), .Q(\CLINT.mtime [28] ), .QN(_10684_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_36 ( .D(_00163_ ), .CK(clock ), .Q(\CLINT.mtime [27] ), .QN(_10683_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_37 ( .D(_00164_ ), .CK(clock ), .Q(\CLINT.mtime [26] ), .QN(_10682_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_38 ( .D(_00165_ ), .CK(clock ), .Q(\CLINT.mtime [25] ), .QN(_10681_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_39 ( .D(_00166_ ), .CK(clock ), .Q(\CLINT.mtime [24] ), .QN(_10680_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_4 ( .D(_00167_ ), .CK(clock ), .Q(\CLINT.mtime [59] ), .QN(_10679_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_40 ( .D(_00168_ ), .CK(clock ), .Q(\CLINT.mtime [23] ), .QN(_10678_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_41 ( .D(_00169_ ), .CK(clock ), .Q(\CLINT.mtime [22] ), .QN(_10677_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_42 ( .D(_00170_ ), .CK(clock ), .Q(\CLINT.mtime [21] ), .QN(_10676_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_43 ( .D(_00171_ ), .CK(clock ), .Q(\CLINT.mtime [20] ), .QN(_10675_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_44 ( .D(_00172_ ), .CK(clock ), .Q(\CLINT.mtime [19] ), .QN(_10674_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_45 ( .D(_00173_ ), .CK(clock ), .Q(\CLINT.mtime [18] ), .QN(_10673_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_46 ( .D(_00174_ ), .CK(clock ), .Q(\CLINT.mtime [17] ), .QN(_10672_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_47 ( .D(_00175_ ), .CK(clock ), .Q(\CLINT.mtime [16] ), .QN(_10671_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_48 ( .D(_00176_ ), .CK(clock ), .Q(\CLINT.mtime [15] ), .QN(_10670_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_49 ( .D(_00177_ ), .CK(clock ), .Q(\CLINT.mtime [14] ), .QN(_10669_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_5 ( .D(_00178_ ), .CK(clock ), .Q(\CLINT.mtime [58] ), .QN(_10668_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_50 ( .D(_00179_ ), .CK(clock ), .Q(\CLINT.mtime [13] ), .QN(_10667_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_51 ( .D(_00180_ ), .CK(clock ), .Q(\CLINT.mtime [12] ), .QN(_10666_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_52 ( .D(_00181_ ), .CK(clock ), .Q(\CLINT.mtime [11] ), .QN(_10665_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_53 ( .D(_00182_ ), .CK(clock ), .Q(\CLINT.mtime [10] ), .QN(_10664_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_54 ( .D(_00183_ ), .CK(clock ), .Q(\CLINT.mtime [9] ), .QN(_10663_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_55 ( .D(_00184_ ), .CK(clock ), .Q(\CLINT.mtime [8] ), .QN(_10662_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_56 ( .D(_00185_ ), .CK(clock ), .Q(\CLINT.mtime [7] ), .QN(_10661_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_57 ( .D(_00186_ ), .CK(clock ), .Q(\CLINT.mtime [6] ), .QN(_10660_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_58 ( .D(_00187_ ), .CK(clock ), .Q(\CLINT.mtime [5] ), .QN(_10659_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_59 ( .D(_00188_ ), .CK(clock ), .Q(\CLINT.mtime [4] ), .QN(_10658_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_6 ( .D(_00189_ ), .CK(clock ), .Q(\CLINT.mtime [57] ), .QN(_10657_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_60 ( .D(_00190_ ), .CK(clock ), .Q(\CLINT.mtime [3] ), .QN(_10656_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_61 ( .D(_00191_ ), .CK(clock ), .Q(\CLINT.mtime [2] ), .QN(_10655_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_62 ( .D(_00192_ ), .CK(clock ), .Q(\CLINT.mtime [1] ), .QN(_10654_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_63 ( .D(_00193_ ), .CK(clock ), .Q(\CLINT.mtime [0] ), .QN(\CLINT.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_7 ( .D(_00194_ ), .CK(clock ), .Q(\CLINT.mtime [56] ), .QN(_10653_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_8 ( .D(_00195_ ), .CK(clock ), .Q(\CLINT.mtime [55] ), .QN(_10652_ ) );
DFF_X1 \CLINT.mtime_$_SDFF_PP0__Q_9 ( .D(_00196_ ), .CK(clock ), .Q(\CLINT.mtime [54] ), .QN(_10651_ ) );
DFF_X1 \EXU.counter_$_SDFFE_PP0N__Q ( .D(_00197_ ), .CK(clock ), .Q(\EXU.counter [1] ), .QN(_10650_ ) );
DFF_X1 \EXU.counter_$_SDFFE_PP0N__Q_1 ( .D(_00198_ ), .CK(clock ), .Q(\EXU.counter [0] ), .QN(\EXU.counter_$_SDFFE_PP0N__Q_1_D [0] ) );
DFF_X1 \EXU.csrs_wen_o_$_SDFFCE_PP0P__Q ( .D(_00199_ ), .CK(clock ), .Q(\EXU.csrs_wen_o [2] ), .QN(_10649_ ) );
DFF_X1 \EXU.csrs_wen_o_$_SDFFCE_PP0P__Q_1 ( .D(_00200_ ), .CK(clock ), .Q(\EXU.csrs_wen_o [3] ), .QN(_10648_ ) );
DFF_X1 \EXU.csrs_wen_o_$_SDFFCE_PP0P__Q_2 ( .D(_00201_ ), .CK(clock ), .Q(\EXU.csrs_wen_o [1] ), .QN(_10647_ ) );
DFF_X1 \EXU.csrs_wen_o_$_SDFFCE_PP0P__Q_3 ( .D(_00202_ ), .CK(clock ), .Q(\EXU.csrs_wen_o [0] ), .QN(_10646_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q ( .D(_00203_ ), .CK(clock ), .Q(\EXU.dnpc_o [31] ), .QN(_10645_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_1 ( .D(_00204_ ), .CK(clock ), .Q(\EXU.dnpc_o [30] ), .QN(_10644_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_10 ( .D(_00205_ ), .CK(clock ), .Q(\EXU.dnpc_o [21] ), .QN(_10643_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_11 ( .D(_00206_ ), .CK(clock ), .Q(\EXU.dnpc_o [20] ), .QN(_10642_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_12 ( .D(_00207_ ), .CK(clock ), .Q(\EXU.dnpc_o [19] ), .QN(_10641_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_13 ( .D(_00208_ ), .CK(clock ), .Q(\EXU.dnpc_o [18] ), .QN(_10640_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_14 ( .D(_00209_ ), .CK(clock ), .Q(\EXU.dnpc_o [17] ), .QN(_10639_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_15 ( .D(_00210_ ), .CK(clock ), .Q(\EXU.dnpc_o [16] ), .QN(_10638_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_16 ( .D(_00211_ ), .CK(clock ), .Q(\EXU.dnpc_o [15] ), .QN(_10637_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_17 ( .D(_00212_ ), .CK(clock ), .Q(\EXU.dnpc_o [14] ), .QN(_10636_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_18 ( .D(_00213_ ), .CK(clock ), .Q(\EXU.dnpc_o [13] ), .QN(_10635_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_19 ( .D(_00214_ ), .CK(clock ), .Q(\EXU.dnpc_o [12] ), .QN(_10634_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_2 ( .D(_00215_ ), .CK(clock ), .Q(\EXU.dnpc_o [29] ), .QN(_10633_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_20 ( .D(_00216_ ), .CK(clock ), .Q(\EXU.dnpc_o [11] ), .QN(_10632_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_21 ( .D(_00217_ ), .CK(clock ), .Q(\EXU.dnpc_o [10] ), .QN(_10631_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_22 ( .D(_00218_ ), .CK(clock ), .Q(\EXU.dnpc_o [9] ), .QN(_10630_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_23 ( .D(_00219_ ), .CK(clock ), .Q(\EXU.dnpc_o [8] ), .QN(_10629_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_24 ( .D(_00220_ ), .CK(clock ), .Q(\EXU.dnpc_o [7] ), .QN(_10628_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_25 ( .D(_00221_ ), .CK(clock ), .Q(\EXU.dnpc_o [6] ), .QN(_10627_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_26 ( .D(_00222_ ), .CK(clock ), .Q(\EXU.dnpc_o [5] ), .QN(_10626_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_27 ( .D(_00223_ ), .CK(clock ), .Q(\EXU.dnpc_o [4] ), .QN(_10625_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_28 ( .D(_00224_ ), .CK(clock ), .Q(\EXU.dnpc_o [3] ), .QN(_10624_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_29 ( .D(_00225_ ), .CK(clock ), .Q(\EXU.dnpc_o [2] ), .QN(_10623_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_3 ( .D(_00226_ ), .CK(clock ), .Q(\EXU.dnpc_o [28] ), .QN(_10622_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_30 ( .D(_00227_ ), .CK(clock ), .Q(\EXU.dnpc_o [1] ), .QN(_10621_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_31 ( .D(_00228_ ), .CK(clock ), .Q(\EXU.dnpc_o [0] ), .QN(_10620_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_4 ( .D(_00229_ ), .CK(clock ), .Q(\EXU.dnpc_o [27] ), .QN(_10619_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_5 ( .D(_00230_ ), .CK(clock ), .Q(\EXU.dnpc_o [26] ), .QN(_10618_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_6 ( .D(_00231_ ), .CK(clock ), .Q(\EXU.dnpc_o [25] ), .QN(_10617_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_7 ( .D(_00232_ ), .CK(clock ), .Q(\EXU.dnpc_o [24] ), .QN(_10616_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_8 ( .D(_00233_ ), .CK(clock ), .Q(\EXU.dnpc_o [23] ), .QN(_10615_ ) );
DFF_X1 \EXU.dnpc_o_$_SDFFCE_PP0P__Q_9 ( .D(_00234_ ), .CK(clock ), .Q(\EXU.dnpc_o [22] ), .QN(_10614_ ) );
DFF_X1 \EXU.gpr_wen_o_$_SDFFE_PP0P__Q ( .D(_00235_ ), .CK(clock ), .Q(\EXU.gpr_wen_o ), .QN(_10613_ ) );
DFF_X1 \EXU.rd_o_$_SDFFCE_PN0P__Q ( .D(_00236_ ), .CK(clock ), .Q(\EXU.rd_o [3] ), .QN(_10612_ ) );
DFF_X1 \EXU.rd_o_$_SDFFCE_PN0P__Q_1 ( .D(_00237_ ), .CK(clock ), .Q(\EXU.rd_o [2] ), .QN(_10611_ ) );
DFF_X1 \EXU.rd_o_$_SDFFCE_PN0P__Q_2 ( .D(_00238_ ), .CK(clock ), .Q(\EXU.rd_o [1] ), .QN(_10610_ ) );
DFF_X1 \EXU.rd_o_$_SDFFCE_PN0P__Q_3 ( .D(_00239_ ), .CK(clock ), .Q(\EXU.rd_o [0] ), .QN(_10609_ ) );
DFF_X1 \EXU.state_$_SDFFE_PP0P__Q ( .D(_00240_ ), .CK(clock ), .Q(\EXU.state ), .QN(\LSU.ls_read_done_$_OR__B_Y_$_ORNOT__A_Y_$_ANDNOT__A_Y_$_OR__A_1_B ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q ( .D(_00241_ ), .CK(clock ), .Q(\EXU.xrd_o [31] ), .QN(_10608_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_1 ( .D(_00242_ ), .CK(clock ), .Q(\EXU.xrd_o [30] ), .QN(_10607_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_10 ( .D(_00243_ ), .CK(clock ), .Q(\EXU.xrd_o [21] ), .QN(_10606_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_11 ( .D(_00244_ ), .CK(clock ), .Q(\EXU.xrd_o [20] ), .QN(_10605_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_12 ( .D(_00245_ ), .CK(clock ), .Q(\EXU.xrd_o [19] ), .QN(_10604_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_13 ( .D(_00246_ ), .CK(clock ), .Q(\EXU.xrd_o [18] ), .QN(_10603_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_14 ( .D(_00247_ ), .CK(clock ), .Q(\EXU.xrd_o [17] ), .QN(_10602_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_15 ( .D(_00248_ ), .CK(clock ), .Q(\EXU.xrd_o [16] ), .QN(_10601_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_16 ( .D(_00249_ ), .CK(clock ), .Q(\EXU.xrd_o [15] ), .QN(_10600_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_17 ( .D(_00250_ ), .CK(clock ), .Q(\EXU.xrd_o [14] ), .QN(_10599_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_18 ( .D(_00251_ ), .CK(clock ), .Q(\EXU.xrd_o [13] ), .QN(_10598_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_19 ( .D(_00252_ ), .CK(clock ), .Q(\EXU.xrd_o [12] ), .QN(_10597_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_2 ( .D(_00253_ ), .CK(clock ), .Q(\EXU.xrd_o [29] ), .QN(_10596_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_20 ( .D(_00254_ ), .CK(clock ), .Q(\EXU.xrd_o [11] ), .QN(_10595_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_21 ( .D(_00255_ ), .CK(clock ), .Q(\EXU.xrd_o [10] ), .QN(_10594_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_22 ( .D(_00256_ ), .CK(clock ), .Q(\EXU.xrd_o [9] ), .QN(_10593_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_23 ( .D(_00257_ ), .CK(clock ), .Q(\EXU.xrd_o [8] ), .QN(_10592_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_24 ( .D(_00258_ ), .CK(clock ), .Q(\EXU.xrd_o [7] ), .QN(_10591_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_25 ( .D(_00259_ ), .CK(clock ), .Q(\EXU.xrd_o [6] ), .QN(_10590_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_26 ( .D(_00260_ ), .CK(clock ), .Q(\EXU.xrd_o [5] ), .QN(_10589_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_27 ( .D(_00261_ ), .CK(clock ), .Q(\EXU.xrd_o [4] ), .QN(_10588_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_28 ( .D(_00262_ ), .CK(clock ), .Q(\EXU.xrd_o [3] ), .QN(_10587_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_29 ( .D(_00263_ ), .CK(clock ), .Q(\EXU.xrd_o [2] ), .QN(_10586_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_3 ( .D(_00264_ ), .CK(clock ), .Q(\EXU.xrd_o [28] ), .QN(_10585_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_30 ( .D(_00265_ ), .CK(clock ), .Q(\EXU.xrd_o [1] ), .QN(_10584_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_31 ( .D(_00266_ ), .CK(clock ), .Q(\EXU.xrd_o [0] ), .QN(_10583_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_4 ( .D(_00267_ ), .CK(clock ), .Q(\EXU.xrd_o [27] ), .QN(_10582_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_5 ( .D(_00268_ ), .CK(clock ), .Q(\EXU.xrd_o [26] ), .QN(_10581_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_6 ( .D(_00269_ ), .CK(clock ), .Q(\EXU.xrd_o [25] ), .QN(_10580_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_7 ( .D(_00270_ ), .CK(clock ), .Q(\EXU.xrd_o [24] ), .QN(_10579_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_8 ( .D(_00271_ ), .CK(clock ), .Q(\EXU.xrd_o [23] ), .QN(_10578_ ) );
DFF_X1 \EXU.xrd_o_$_SDFFCE_PP0P__Q_9 ( .D(_00272_ ), .CK(clock ), .Q(\EXU.xrd_o [22] ), .QN(_10793_ ) );
DFF_X1 \ICACHE.axi_rvalid_enable_$_DFF_P__Q ( .D(\ICACHE.axi_rvalid ), .CK(clock ), .Q(\ICACHE.axi_rvalid_enable ), .QN(_10577_ ) );
DFF_X1 \ICACHE.burst_counter_$_DFFE_PP__Q ( .D(_00273_ ), .CK(clock ), .Q(\ICACHE.burst_counter [1] ), .QN(_10576_ ) );
DFF_X1 \ICACHE.burst_counter_$_DFFE_PP__Q_1 ( .D(_00274_ ), .CK(clock ), .Q(\ICACHE.burst_counter [0] ), .QN(\ICACHE.burst_counter_$_DFFE_PP__Q_1_D_$_MUX__Y_B ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q ( .D(_00275_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][31] ), .QN(_10575_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_1 ( .D(_00276_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][30] ), .QN(_10574_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_10 ( .D(_00277_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][21] ), .QN(_10573_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_11 ( .D(_00278_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][20] ), .QN(_10572_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_12 ( .D(_00279_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][19] ), .QN(_10571_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_13 ( .D(_00280_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][18] ), .QN(_10570_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_14 ( .D(_00281_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][17] ), .QN(_10569_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_15 ( .D(_00282_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][16] ), .QN(_10568_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_16 ( .D(_00283_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][15] ), .QN(_10567_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_17 ( .D(_00284_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][14] ), .QN(_10566_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_18 ( .D(_00285_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][13] ), .QN(_10565_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_19 ( .D(_00286_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][12] ), .QN(_10564_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_2 ( .D(_00287_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][29] ), .QN(_10563_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_20 ( .D(_00288_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][11] ), .QN(_10562_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_21 ( .D(_00289_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][10] ), .QN(_10561_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_22 ( .D(_00290_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][9] ), .QN(_10560_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_23 ( .D(_00291_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][8] ), .QN(_10559_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_24 ( .D(_00292_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][7] ), .QN(_10558_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_25 ( .D(_00293_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][6] ), .QN(_10557_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_26 ( .D(_00294_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][5] ), .QN(_10556_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_27 ( .D(_00295_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][4] ), .QN(_10555_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_28 ( .D(_00296_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][3] ), .QN(_10554_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_29 ( .D(_00297_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][2] ), .QN(_10553_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_3 ( .D(_00298_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][28] ), .QN(_10552_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_4 ( .D(_00299_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][27] ), .QN(_10551_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_5 ( .D(_00300_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][26] ), .QN(_10550_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_6 ( .D(_00301_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][25] ), .QN(_10549_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_7 ( .D(_00302_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][24] ), .QN(_10548_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_8 ( .D(_00303_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][23] ), .QN(_10547_ ) );
DFF_X1 \ICACHE.cache_reg[0]_$_DFFE_PP__Q_9 ( .D(_00304_ ), .CK(clock ), .Q(\ICACHE.cache_reg[0][22] ), .QN(_10546_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q ( .D(_00305_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][31] ), .QN(_10545_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_1 ( .D(_00306_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][30] ), .QN(_10544_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_10 ( .D(_00307_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][21] ), .QN(_10543_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_11 ( .D(_00308_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][20] ), .QN(_10542_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_12 ( .D(_00309_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][19] ), .QN(_10541_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_13 ( .D(_00310_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][18] ), .QN(_10540_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_14 ( .D(_00311_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][17] ), .QN(_10539_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_15 ( .D(_00312_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][16] ), .QN(_10538_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_16 ( .D(_00313_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][15] ), .QN(_10537_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_17 ( .D(_00314_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][14] ), .QN(_10536_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_18 ( .D(_00315_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][13] ), .QN(_10535_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_19 ( .D(_00316_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][12] ), .QN(_10534_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_2 ( .D(_00317_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][29] ), .QN(_10533_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_20 ( .D(_00318_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][11] ), .QN(_10532_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_21 ( .D(_00319_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][10] ), .QN(_10531_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_22 ( .D(_00320_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][9] ), .QN(_10530_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_23 ( .D(_00321_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][8] ), .QN(_10529_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_24 ( .D(_00322_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][7] ), .QN(_10528_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_25 ( .D(_00323_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][6] ), .QN(_10527_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_26 ( .D(_00324_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][5] ), .QN(_10526_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_27 ( .D(_00325_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][4] ), .QN(_10525_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_28 ( .D(_00326_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][3] ), .QN(_10524_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_29 ( .D(_00327_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][2] ), .QN(_10523_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_3 ( .D(_00328_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][28] ), .QN(_10522_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_4 ( .D(_00329_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][27] ), .QN(_10521_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_5 ( .D(_00330_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][26] ), .QN(_10520_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_6 ( .D(_00331_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][25] ), .QN(_10519_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_7 ( .D(_00332_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][24] ), .QN(_10518_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_8 ( .D(_00333_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][23] ), .QN(_10517_ ) );
DFF_X1 \ICACHE.cache_reg[1]_$_DFFE_PP__Q_9 ( .D(_00334_ ), .CK(clock ), .Q(\ICACHE.cache_reg[1][22] ), .QN(_10516_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q ( .D(_00335_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][31] ), .QN(_10515_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_1 ( .D(_00336_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][30] ), .QN(_10514_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_10 ( .D(_00337_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][21] ), .QN(_10513_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_11 ( .D(_00338_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][20] ), .QN(_10512_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_12 ( .D(_00339_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][19] ), .QN(_10511_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_13 ( .D(_00340_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][18] ), .QN(_10510_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_14 ( .D(_00341_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][17] ), .QN(_10509_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_15 ( .D(_00342_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][16] ), .QN(_10508_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_16 ( .D(_00343_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][15] ), .QN(_10507_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_17 ( .D(_00344_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][14] ), .QN(_10506_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_18 ( .D(_00345_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][13] ), .QN(_10505_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_19 ( .D(_00346_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][12] ), .QN(_10504_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_2 ( .D(_00347_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][29] ), .QN(_10503_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_20 ( .D(_00348_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][11] ), .QN(_10502_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_21 ( .D(_00349_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][10] ), .QN(_10501_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_22 ( .D(_00350_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][9] ), .QN(_10500_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_23 ( .D(_00351_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][8] ), .QN(_10499_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_24 ( .D(_00352_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][7] ), .QN(_10498_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_25 ( .D(_00353_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][6] ), .QN(_10497_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_26 ( .D(_00354_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][5] ), .QN(_10496_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_27 ( .D(_00355_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][4] ), .QN(_10495_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_28 ( .D(_00356_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][3] ), .QN(_10494_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_29 ( .D(_00357_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][2] ), .QN(_10493_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_3 ( .D(_00358_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][28] ), .QN(_10492_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_4 ( .D(_00359_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][27] ), .QN(_10491_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_5 ( .D(_00360_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][26] ), .QN(_10490_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_6 ( .D(_00361_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][25] ), .QN(_10489_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_7 ( .D(_00362_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][24] ), .QN(_10488_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_8 ( .D(_00363_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][23] ), .QN(_10487_ ) );
DFF_X1 \ICACHE.cache_reg[2]_$_DFFE_PP__Q_9 ( .D(_00364_ ), .CK(clock ), .Q(\ICACHE.cache_reg[2][22] ), .QN(_10486_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q ( .D(_00365_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][31] ), .QN(_10485_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_1 ( .D(_00366_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][30] ), .QN(_10484_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_10 ( .D(_00367_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][21] ), .QN(_10483_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_11 ( .D(_00368_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][20] ), .QN(_10482_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_12 ( .D(_00369_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][19] ), .QN(_10481_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_13 ( .D(_00370_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][18] ), .QN(_10480_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_14 ( .D(_00371_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][17] ), .QN(_10479_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_15 ( .D(_00372_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][16] ), .QN(_10478_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_16 ( .D(_00373_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][15] ), .QN(_10477_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_17 ( .D(_00374_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][14] ), .QN(_10476_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_18 ( .D(_00375_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][13] ), .QN(_10475_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_19 ( .D(_00376_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][12] ), .QN(_10474_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_2 ( .D(_00377_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][29] ), .QN(_10473_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_20 ( .D(_00378_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][11] ), .QN(_10472_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_21 ( .D(_00379_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][10] ), .QN(_10471_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_22 ( .D(_00380_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][9] ), .QN(_10470_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_23 ( .D(_00381_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][8] ), .QN(_10469_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_24 ( .D(_00382_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][7] ), .QN(_10468_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_25 ( .D(_00383_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][6] ), .QN(_10467_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_26 ( .D(_00384_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][5] ), .QN(_10466_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_27 ( .D(_00385_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][4] ), .QN(_10465_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_28 ( .D(_00386_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][3] ), .QN(_10464_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_29 ( .D(_00387_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][2] ), .QN(_10463_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_3 ( .D(_00388_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][28] ), .QN(_10462_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_4 ( .D(_00389_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][27] ), .QN(_10461_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_5 ( .D(_00390_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][26] ), .QN(_10460_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_6 ( .D(_00391_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][25] ), .QN(_10459_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_7 ( .D(_00392_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][24] ), .QN(_10458_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_8 ( .D(_00393_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][23] ), .QN(_10457_ ) );
DFF_X1 \ICACHE.cache_reg[3]_$_DFFE_PP__Q_9 ( .D(_00394_ ), .CK(clock ), .Q(\ICACHE.cache_reg[3][22] ), .QN(_10456_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q ( .D(_00395_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][31] ), .QN(_10455_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_1 ( .D(_00396_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][30] ), .QN(_10454_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_10 ( .D(_00397_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][21] ), .QN(_10453_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_11 ( .D(_00398_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][20] ), .QN(_10452_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_12 ( .D(_00399_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][19] ), .QN(_10451_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_13 ( .D(_00400_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][18] ), .QN(_10450_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_14 ( .D(_00401_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][17] ), .QN(_10449_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_15 ( .D(_00402_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][16] ), .QN(_10448_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_16 ( .D(_00403_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][15] ), .QN(_10447_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_17 ( .D(_00404_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][14] ), .QN(_10446_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_18 ( .D(_00405_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][13] ), .QN(_10445_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_19 ( .D(_00406_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][12] ), .QN(_10444_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_2 ( .D(_00407_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][29] ), .QN(_10443_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_20 ( .D(_00408_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][11] ), .QN(_10442_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_21 ( .D(_00409_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][10] ), .QN(_10441_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_22 ( .D(_00410_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][9] ), .QN(_10440_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_23 ( .D(_00411_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][8] ), .QN(_10439_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_24 ( .D(_00412_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][7] ), .QN(_10438_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_25 ( .D(_00413_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][6] ), .QN(_10437_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_26 ( .D(_00414_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][5] ), .QN(_10436_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_27 ( .D(_00415_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][4] ), .QN(_10435_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_28 ( .D(_00416_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][3] ), .QN(_10434_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_29 ( .D(_00417_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][2] ), .QN(_10433_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_3 ( .D(_00418_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][28] ), .QN(_10432_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_4 ( .D(_00419_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][27] ), .QN(_10431_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_5 ( .D(_00420_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][26] ), .QN(_10430_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_6 ( .D(_00421_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][25] ), .QN(_10429_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_7 ( .D(_00422_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][24] ), .QN(_10428_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_8 ( .D(_00423_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][23] ), .QN(_10427_ ) );
DFF_X1 \ICACHE.cache_reg[4]_$_DFFE_PP__Q_9 ( .D(_00424_ ), .CK(clock ), .Q(\ICACHE.cache_reg[4][22] ), .QN(_10426_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q ( .D(_00425_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][31] ), .QN(_10425_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_1 ( .D(_00426_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][30] ), .QN(_10424_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_10 ( .D(_00427_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][21] ), .QN(_10423_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_11 ( .D(_00428_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][20] ), .QN(_10422_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_12 ( .D(_00429_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][19] ), .QN(_10421_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_13 ( .D(_00430_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][18] ), .QN(_10420_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_14 ( .D(_00431_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][17] ), .QN(_10419_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_15 ( .D(_00432_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][16] ), .QN(_10418_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_16 ( .D(_00433_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][15] ), .QN(_10417_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_17 ( .D(_00434_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][14] ), .QN(_10416_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_18 ( .D(_00435_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][13] ), .QN(_10415_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_19 ( .D(_00436_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][12] ), .QN(_10414_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_2 ( .D(_00437_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][29] ), .QN(_10413_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_20 ( .D(_00438_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][11] ), .QN(_10412_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_21 ( .D(_00439_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][10] ), .QN(_10411_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_22 ( .D(_00440_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][9] ), .QN(_10410_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_23 ( .D(_00441_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][8] ), .QN(_10409_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_24 ( .D(_00442_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][7] ), .QN(_10408_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_25 ( .D(_00443_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][6] ), .QN(_10407_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_26 ( .D(_00444_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][5] ), .QN(_10406_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_27 ( .D(_00445_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][4] ), .QN(_10405_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_28 ( .D(_00446_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][3] ), .QN(_10404_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_29 ( .D(_00447_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][2] ), .QN(_10403_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_3 ( .D(_00448_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][28] ), .QN(_10402_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_4 ( .D(_00449_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][27] ), .QN(_10401_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_5 ( .D(_00450_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][26] ), .QN(_10400_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_6 ( .D(_00451_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][25] ), .QN(_10399_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_7 ( .D(_00452_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][24] ), .QN(_10398_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_8 ( .D(_00453_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][23] ), .QN(_10397_ ) );
DFF_X1 \ICACHE.cache_reg[5]_$_DFFE_PP__Q_9 ( .D(_00454_ ), .CK(clock ), .Q(\ICACHE.cache_reg[5][22] ), .QN(_10396_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q ( .D(_00455_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][31] ), .QN(_10395_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_1 ( .D(_00456_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][30] ), .QN(_10394_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_10 ( .D(_00457_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][21] ), .QN(_10393_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_11 ( .D(_00458_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][20] ), .QN(_10392_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_12 ( .D(_00459_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][19] ), .QN(_10391_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_13 ( .D(_00460_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][18] ), .QN(_10390_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_14 ( .D(_00461_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][17] ), .QN(_10389_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_15 ( .D(_00462_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][16] ), .QN(_10388_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_16 ( .D(_00463_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][15] ), .QN(_10387_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_17 ( .D(_00464_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][14] ), .QN(_10386_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_18 ( .D(_00465_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][13] ), .QN(_10385_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_19 ( .D(_00466_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][12] ), .QN(_10384_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_2 ( .D(_00467_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][29] ), .QN(_10383_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_20 ( .D(_00468_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][11] ), .QN(_10382_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_21 ( .D(_00469_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][10] ), .QN(_10381_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_22 ( .D(_00470_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][9] ), .QN(_10380_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_23 ( .D(_00471_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][8] ), .QN(_10379_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_24 ( .D(_00472_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][7] ), .QN(_10378_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_25 ( .D(_00473_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][6] ), .QN(_10377_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_26 ( .D(_00474_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][5] ), .QN(_10376_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_27 ( .D(_00475_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][4] ), .QN(_10375_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_28 ( .D(_00476_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][3] ), .QN(_10374_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_29 ( .D(_00477_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][2] ), .QN(_10373_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_3 ( .D(_00478_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][28] ), .QN(_10372_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_4 ( .D(_00479_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][27] ), .QN(_10371_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_5 ( .D(_00480_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][26] ), .QN(_10370_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_6 ( .D(_00481_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][25] ), .QN(_10369_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_7 ( .D(_00482_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][24] ), .QN(_10368_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_8 ( .D(_00483_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][23] ), .QN(_10367_ ) );
DFF_X1 \ICACHE.cache_reg[6]_$_DFFE_PP__Q_9 ( .D(_00484_ ), .CK(clock ), .Q(\ICACHE.cache_reg[6][22] ), .QN(_10366_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q ( .D(_00485_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][31] ), .QN(_10365_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_1 ( .D(_00486_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][30] ), .QN(_10364_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_10 ( .D(_00487_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][21] ), .QN(_10363_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_11 ( .D(_00488_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][20] ), .QN(_10362_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_12 ( .D(_00489_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][19] ), .QN(_10361_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_13 ( .D(_00490_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][18] ), .QN(_10360_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_14 ( .D(_00491_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][17] ), .QN(_10359_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_15 ( .D(_00492_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][16] ), .QN(_10358_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_16 ( .D(_00493_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][15] ), .QN(_10357_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_17 ( .D(_00494_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][14] ), .QN(_10356_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_18 ( .D(_00495_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][13] ), .QN(_10355_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_19 ( .D(_00496_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][12] ), .QN(_10354_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_2 ( .D(_00497_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][29] ), .QN(_10353_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_20 ( .D(_00498_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][11] ), .QN(_10352_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_21 ( .D(_00499_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][10] ), .QN(_10351_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_22 ( .D(_00500_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][9] ), .QN(_10350_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_23 ( .D(_00501_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][8] ), .QN(_10349_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_24 ( .D(_00502_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][7] ), .QN(_10348_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_25 ( .D(_00503_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][6] ), .QN(_10347_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_26 ( .D(_00504_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][5] ), .QN(_10346_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_27 ( .D(_00505_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][4] ), .QN(_10345_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_28 ( .D(_00506_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][3] ), .QN(_10344_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_29 ( .D(_00507_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][2] ), .QN(_10343_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_3 ( .D(_00508_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][28] ), .QN(_10342_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_4 ( .D(_00509_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][27] ), .QN(_10341_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_5 ( .D(_00510_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][26] ), .QN(_10340_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_6 ( .D(_00511_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][25] ), .QN(_10339_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_7 ( .D(_00512_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][24] ), .QN(_10338_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_8 ( .D(_00513_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][23] ), .QN(_10337_ ) );
DFF_X1 \ICACHE.cache_reg[7]_$_DFFE_PP__Q_9 ( .D(_00514_ ), .CK(clock ), .Q(\ICACHE.cache_reg[7][22] ), .QN(_10336_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q ( .D(_00515_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [15] ), .QN(_10335_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_1 ( .D(_00516_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [14] ), .QN(_10334_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_10 ( .D(_00517_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [5] ), .QN(_10333_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_11 ( .D(_00518_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [4] ), .QN(_10332_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_12 ( .D(_00519_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [3] ), .QN(\ICACHE.state_$_MUX__S_B ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_13 ( .D(_00520_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [2] ), .QN(_10331_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_2 ( .D(_00521_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [13] ), .QN(_10330_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_3 ( .D(_00522_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [12] ), .QN(_10329_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_4 ( .D(_00523_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [11] ), .QN(_10328_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_5 ( .D(_00524_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [10] ), .QN(_10327_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_6 ( .D(_00525_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [9] ), .QN(_10326_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_7 ( .D(_00526_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [8] ), .QN(_10325_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_8 ( .D(_00527_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [7] ), .QN(_10324_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PN__Q_9 ( .D(_00528_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [6] ), .QN(_10323_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q ( .D(_00529_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [31] ), .QN(_10322_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_1 ( .D(_00530_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [30] ), .QN(_10321_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_10 ( .D(_00531_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [21] ), .QN(_10320_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_11 ( .D(_00532_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [20] ), .QN(_10319_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_12 ( .D(_00533_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [19] ), .QN(_10318_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_13 ( .D(_00534_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [18] ), .QN(_10317_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_14 ( .D(_00535_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [17] ), .QN(_10316_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_15 ( .D(_00536_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [16] ), .QN(_10315_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_16 ( .D(_00537_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [1] ), .QN(_10314_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_17 ( .D(_00538_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [0] ), .QN(_10313_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_2 ( .D(_00539_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [29] ), .QN(_10312_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_3 ( .D(_00540_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [28] ), .QN(_10311_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_4 ( .D(_00541_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [27] ), .QN(_10310_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_5 ( .D(_00542_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [26] ), .QN(_10309_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_6 ( .D(_00543_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [25] ), .QN(_10308_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_7 ( .D(_00544_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [24] ), .QN(_10307_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_8 ( .D(_00545_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [23] ), .QN(_10306_ ) );
DFF_X1 \ICACHE.s_axi_araddr_$_DFFE_PP__Q_9 ( .D(_00546_ ), .CK(clock ), .Q(\ICACHE.s_axi_araddr [22] ), .QN(_10305_ ) );
DFF_X1 \ICACHE.s_axi_arlen_$_SDFFCE_PP0P__Q ( .D(_00547_ ), .CK(clock ), .Q(\ICACHE.s_axi_arlen [3] ), .QN(_10304_ ) );
DFF_X1 \ICACHE.s_axi_arlen_$_SDFFCE_PP0P__Q_2 ( .D(_00548_ ), .CK(clock ), .Q(\ICACHE.s_axi_arlen [1] ), .QN(_10303_ ) );
DFF_X1 \ICACHE.s_axi_arlen_$_SDFFCE_PP0P__Q_3 ( .D(_00549_ ), .CK(clock ), .Q(\ICACHE.s_axi_arlen [0] ), .QN(_10302_ ) );
DFF_X1 \ICACHE.s_axi_arvalid_$_SDFFE_PP0P__Q ( .D(_00550_ ), .CK(clock ), .Q(\ICACHE.s_axi_arvalid ), .QN(io_master_arvalid_$_ANDNOT__Y_B_$_MUX__Y_A ) );
DFF_X1 \ICACHE.state_$_SDFF_PP0__Q ( .D(_00551_ ), .CK(clock ), .Q(\ICACHE.s_axi_rready ), .QN(\ICACHE.m_axi_arready ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q ( .D(_00552_ ), .CK(clock ), .Q(\ICACHE.tag_check [15] ), .QN(_10301_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_1 ( .D(_00553_ ), .CK(clock ), .Q(\ICACHE.tag_check [14] ), .QN(_10300_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_10 ( .D(_00554_ ), .CK(clock ), .Q(\ICACHE.tag_check [5] ), .QN(_10299_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_11 ( .D(_00555_ ), .CK(clock ), .Q(\ICACHE.tag_check [4] ), .QN(_10298_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_12 ( .D(_00556_ ), .CK(clock ), .Q(\ICACHE.tag_check [3] ), .QN(_10297_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_13 ( .D(_00557_ ), .CK(clock ), .Q(\ICACHE.tag_check [2] ), .QN(_10296_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_14 ( .D(_00558_ ), .CK(clock ), .Q(\ICACHE.tag_check [1] ), .QN(_10295_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_15 ( .D(_00559_ ), .CK(clock ), .Q(\ICACHE.tag_check [0] ), .QN(_10294_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_2 ( .D(_00560_ ), .CK(clock ), .Q(\ICACHE.tag_check [13] ), .QN(_10293_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_3 ( .D(_00561_ ), .CK(clock ), .Q(\ICACHE.tag_check [12] ), .QN(_10292_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_4 ( .D(_00562_ ), .CK(clock ), .Q(\ICACHE.tag_check [11] ), .QN(_10291_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_5 ( .D(_00563_ ), .CK(clock ), .Q(\ICACHE.tag_check [10] ), .QN(_10290_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_6 ( .D(_00564_ ), .CK(clock ), .Q(\ICACHE.tag_check [9] ), .QN(_10289_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_7 ( .D(_00565_ ), .CK(clock ), .Q(\ICACHE.tag_check [8] ), .QN(_10288_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_8 ( .D(_00566_ ), .CK(clock ), .Q(\ICACHE.tag_check [7] ), .QN(_10287_ ) );
DFF_X1 \ICACHE.tag_check_$_DFFE_PP__Q_9 ( .D(_00567_ ), .CK(clock ), .Q(\ICACHE.tag_check [6] ), .QN(_10286_ ) );
DFF_X1 \ICACHE.tag_reg[0]_$_SDFFCE_PN0P__Q ( .D(_00568_ ), .CK(clock ), .Q(\ICACHE.tag_reg[0][10] ), .QN(_10285_ ) );
DFF_X1 \ICACHE.tag_reg[0]_$_SDFFCE_PN0P__Q_1 ( .D(_00569_ ), .CK(clock ), .Q(\ICACHE.tag_reg[0][9] ), .QN(_10284_ ) );
DFF_X1 \ICACHE.tag_reg[0]_$_SDFFCE_PN0P__Q_10 ( .D(_00570_ ), .CK(clock ), .Q(\ICACHE.tag_reg[0][0] ), .QN(_10283_ ) );
DFF_X1 \ICACHE.tag_reg[0]_$_SDFFCE_PN0P__Q_2 ( .D(_00571_ ), .CK(clock ), .Q(\ICACHE.tag_reg[0][8] ), .QN(_10282_ ) );
DFF_X1 \ICACHE.tag_reg[0]_$_SDFFCE_PN0P__Q_3 ( .D(_00572_ ), .CK(clock ), .Q(\ICACHE.tag_reg[0][7] ), .QN(_10281_ ) );
DFF_X1 \ICACHE.tag_reg[0]_$_SDFFCE_PN0P__Q_4 ( .D(_00573_ ), .CK(clock ), .Q(\ICACHE.tag_reg[0][6] ), .QN(_10280_ ) );
DFF_X1 \ICACHE.tag_reg[0]_$_SDFFCE_PN0P__Q_5 ( .D(_00574_ ), .CK(clock ), .Q(\ICACHE.tag_reg[0][5] ), .QN(_10279_ ) );
DFF_X1 \ICACHE.tag_reg[0]_$_SDFFCE_PN0P__Q_6 ( .D(_00575_ ), .CK(clock ), .Q(\ICACHE.tag_reg[0][4] ), .QN(_10278_ ) );
DFF_X1 \ICACHE.tag_reg[0]_$_SDFFCE_PN0P__Q_7 ( .D(_00576_ ), .CK(clock ), .Q(\ICACHE.tag_reg[0][3] ), .QN(_10277_ ) );
DFF_X1 \ICACHE.tag_reg[0]_$_SDFFCE_PN0P__Q_8 ( .D(_00577_ ), .CK(clock ), .Q(\ICACHE.tag_reg[0][2] ), .QN(_10276_ ) );
DFF_X1 \ICACHE.tag_reg[0]_$_SDFFCE_PN0P__Q_9 ( .D(_00578_ ), .CK(clock ), .Q(\ICACHE.tag_reg[0][1] ), .QN(_10275_ ) );
DFF_X1 \ICACHE.tag_reg[1]_$_SDFFCE_PN0P__Q ( .D(_00579_ ), .CK(clock ), .Q(\ICACHE.tag_reg[1][10] ), .QN(_10274_ ) );
DFF_X1 \ICACHE.tag_reg[1]_$_SDFFCE_PN0P__Q_1 ( .D(_00580_ ), .CK(clock ), .Q(\ICACHE.tag_reg[1][9] ), .QN(_10273_ ) );
DFF_X1 \ICACHE.tag_reg[1]_$_SDFFCE_PN0P__Q_10 ( .D(_00581_ ), .CK(clock ), .Q(\ICACHE.tag_reg[1][0] ), .QN(_10272_ ) );
DFF_X1 \ICACHE.tag_reg[1]_$_SDFFCE_PN0P__Q_2 ( .D(_00582_ ), .CK(clock ), .Q(\ICACHE.tag_reg[1][8] ), .QN(_10271_ ) );
DFF_X1 \ICACHE.tag_reg[1]_$_SDFFCE_PN0P__Q_3 ( .D(_00583_ ), .CK(clock ), .Q(\ICACHE.tag_reg[1][7] ), .QN(_10270_ ) );
DFF_X1 \ICACHE.tag_reg[1]_$_SDFFCE_PN0P__Q_4 ( .D(_00584_ ), .CK(clock ), .Q(\ICACHE.tag_reg[1][6] ), .QN(_10269_ ) );
DFF_X1 \ICACHE.tag_reg[1]_$_SDFFCE_PN0P__Q_5 ( .D(_00585_ ), .CK(clock ), .Q(\ICACHE.tag_reg[1][5] ), .QN(_10268_ ) );
DFF_X1 \ICACHE.tag_reg[1]_$_SDFFCE_PN0P__Q_6 ( .D(_00586_ ), .CK(clock ), .Q(\ICACHE.tag_reg[1][4] ), .QN(_10267_ ) );
DFF_X1 \ICACHE.tag_reg[1]_$_SDFFCE_PN0P__Q_7 ( .D(_00587_ ), .CK(clock ), .Q(\ICACHE.tag_reg[1][3] ), .QN(_10266_ ) );
DFF_X1 \ICACHE.tag_reg[1]_$_SDFFCE_PN0P__Q_8 ( .D(_00588_ ), .CK(clock ), .Q(\ICACHE.tag_reg[1][2] ), .QN(_10265_ ) );
DFF_X1 \ICACHE.tag_reg[1]_$_SDFFCE_PN0P__Q_9 ( .D(_00589_ ), .CK(clock ), .Q(\ICACHE.tag_reg[1][1] ), .QN(_10264_ ) );
DFF_X1 \ICACHE.valid_reg[0]_$_SDFFCE_PN0P__Q ( .D(_00590_ ), .CK(clock ), .Q(\ICACHE.valid_reg[0][0] ), .QN(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \ICACHE.valid_reg[0]_$_SDFFCE_PN0P__Q_1 ( .D(_00591_ ), .CK(clock ), .Q(\ICACHE.valid_reg[0][1] ), .QN(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \ICACHE.valid_reg[0]_$_SDFFCE_PN0P__Q_2 ( .D(_00592_ ), .CK(clock ), .Q(\ICACHE.valid_reg[0][2] ), .QN(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \ICACHE.valid_reg[0]_$_SDFFCE_PN0P__Q_3 ( .D(_00593_ ), .CK(clock ), .Q(\ICACHE.valid_reg[0][3] ), .QN(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \ICACHE.valid_reg[1]_$_SDFFCE_PN0P__Q ( .D(_00594_ ), .CK(clock ), .Q(\ICACHE.valid_reg[1][1] ), .QN(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \ICACHE.valid_reg[1]_$_SDFFCE_PN0P__Q_1 ( .D(_00595_ ), .CK(clock ), .Q(\ICACHE.valid_reg[1][2] ), .QN(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \ICACHE.valid_reg[1]_$_SDFFCE_PN0P__Q_2 ( .D(_00596_ ), .CK(clock ), .Q(\ICACHE.valid_reg[1][0] ), .QN(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \ICACHE.valid_reg[1]_$_SDFFCE_PN0P__Q_3 ( .D(_00597_ ), .CK(clock ), .Q(\ICACHE.valid_reg[1][3] ), .QN(\ICACHE.hit_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \IDU.funct3_o_$_DFFE_PP__Q ( .D(_00598_ ), .CK(clock ), .Q(\EXU.funct3_i [2] ), .QN(io_master_arsize_$_ANDNOT__Y_1_B_$_OR__Y_A_$_OR__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_AND__Y_B_$_OR__Y_B ) );
DFF_X1 \IDU.funct3_o_$_DFFE_PP__Q_1 ( .D(_00599_ ), .CK(clock ), .Q(\EXU.funct3_i [1] ), .QN(_10263_ ) );
DFF_X1 \IDU.funct3_o_$_DFFE_PP__Q_2 ( .D(_00600_ ), .CK(clock ), .Q(\EXU.funct3_i [0] ), .QN(_10262_ ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q ( .D(_00601_ ), .CK(clock ), .Q(\EXU.imm_i [31] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_1 ( .D(_00602_ ), .CK(clock ), .Q(\EXU.imm_i [30] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_10 ( .D(_00603_ ), .CK(clock ), .Q(\EXU.imm_i [21] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_11 ( .D(_00604_ ), .CK(clock ), .Q(\EXU.imm_i [20] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_12 ( .D(_00605_ ), .CK(clock ), .Q(\EXU.imm_i [19] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_7_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_13 ( .D(_00606_ ), .CK(clock ), .Q(\EXU.imm_i [18] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_8_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_14 ( .D(_00607_ ), .CK(clock ), .Q(\EXU.imm_i [17] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_15 ( .D(_00608_ ), .CK(clock ), .Q(\EXU.imm_i [16] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_16 ( .D(_00609_ ), .CK(clock ), .Q(\EXU.imm_i [15] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_10_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_17 ( .D(_00610_ ), .CK(clock ), .Q(\EXU.imm_i [14] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_11_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_18 ( .D(_00611_ ), .CK(clock ), .Q(\EXU.imm_i [13] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_19 ( .D(_00612_ ), .CK(clock ), .Q(\EXU.imm_i [12] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_2 ( .D(_00613_ ), .CK(clock ), .Q(\EXU.imm_i [29] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_20 ( .D(_00614_ ), .CK(clock ), .Q(\EXU.imm_i [11] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_21 ( .D(_00615_ ), .CK(clock ), .Q(\EXU.funct7_i ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_14_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_22 ( .D(_00616_ ), .CK(clock ), .Q(\EXU.imm_i [9] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_15_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_23 ( .D(_00617_ ), .CK(clock ), .Q(\EXU.imm_i [8] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_16_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_24 ( .D(_00618_ ), .CK(clock ), .Q(\EXU.imm_i [7] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_17_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_25 ( .D(_00619_ ), .CK(clock ), .Q(\EXU.imm_i [6] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_18_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_26 ( .D(_00620_ ), .CK(clock ), .Q(\EXU.imm_i [5] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_19_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_27 ( .D(_00621_ ), .CK(clock ), .Q(\EXU.imm_i [4] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_20_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_28 ( .D(_00622_ ), .CK(clock ), .Q(\EXU.imm_i [3] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_21_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_29 ( .D(_00623_ ), .CK(clock ), .Q(\EXU.imm_i [2] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_3 ( .D(_00624_ ), .CK(clock ), .Q(\EXU.imm_i [28] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_30 ( .D(_00625_ ), .CK(clock ), .Q(\EXU.imm_i [1] ), .QN(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_31 ( .D(_00626_ ), .CK(clock ), .Q(\EXU.imm_i [0] ), .QN(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_4 ( .D(_00627_ ), .CK(clock ), .Q(\EXU.imm_i [27] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_2_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_5 ( .D(_00628_ ), .CK(clock ), .Q(\EXU.imm_i [26] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_6 ( .D(_00629_ ), .CK(clock ), .Q(\EXU.imm_i [25] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_7 ( .D(_00630_ ), .CK(clock ), .Q(\EXU.imm_i [24] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_8 ( .D(_00631_ ), .CK(clock ), .Q(\EXU.imm_i [23] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_4_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.imm_o_$_DFFE_PP__Q_9 ( .D(_00632_ ), .CK(clock ), .Q(\EXU.imm_i [22] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_5_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.ls_valid_o_$_DFFE_PP__Q ( .D(_00633_ ), .CK(clock ), .Q(\IDU.ls_valid_o ), .QN(_10261_ ) );
DFF_X1 \IDU.op_o_$_DFFE_PP__Q ( .D(_00634_ ), .CK(clock ), .Q(\EXU.op_i [4] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B ) );
DFF_X1 \IDU.op_o_$_DFFE_PP__Q_1 ( .D(_00635_ ), .CK(clock ), .Q(\EXU.op_i [3] ), .QN(_10260_ ) );
DFF_X1 \IDU.op_o_$_DFFE_PP__Q_2 ( .D(_00636_ ), .CK(clock ), .Q(\EXU.op_i [2] ), .QN(_10259_ ) );
DFF_X1 \IDU.op_o_$_DFFE_PP__Q_3 ( .D(_00637_ ), .CK(clock ), .Q(\EXU.op_i [1] ), .QN(_10258_ ) );
DFF_X1 \IDU.op_o_$_DFFE_PP__Q_4 ( .D(_00638_ ), .CK(clock ), .Q(\EXU.op_i [0] ), .QN(_10257_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q ( .D(_00639_ ), .CK(clock ), .Q(\EXU.pc_i [31] ), .QN(_10256_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_1 ( .D(_00640_ ), .CK(clock ), .Q(\EXU.pc_i [30] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_B ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_10 ( .D(_00641_ ), .CK(clock ), .Q(\EXU.pc_i [21] ), .QN(_10255_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_11 ( .D(_00642_ ), .CK(clock ), .Q(\EXU.pc_i [20] ), .QN(_10254_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_12 ( .D(_00643_ ), .CK(clock ), .Q(\EXU.pc_i [19] ), .QN(_10253_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_13 ( .D(_00644_ ), .CK(clock ), .Q(\EXU.pc_i [18] ), .QN(_10252_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_14 ( .D(_00645_ ), .CK(clock ), .Q(\EXU.pc_i [17] ), .QN(_10251_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_15 ( .D(_00646_ ), .CK(clock ), .Q(\EXU.pc_i [16] ), .QN(_10250_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_16 ( .D(_00647_ ), .CK(clock ), .Q(\EXU.pc_i [15] ), .QN(_10249_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_17 ( .D(_00648_ ), .CK(clock ), .Q(\EXU.pc_i [14] ), .QN(_10248_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_18 ( .D(_00649_ ), .CK(clock ), .Q(\EXU.pc_i [13] ), .QN(_10247_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_19 ( .D(_00650_ ), .CK(clock ), .Q(\EXU.pc_i [12] ), .QN(_10246_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_2 ( .D(_00651_ ), .CK(clock ), .Q(\EXU.pc_i [29] ), .QN(_10245_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_20 ( .D(_00652_ ), .CK(clock ), .Q(\EXU.pc_i [11] ), .QN(_10244_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_21 ( .D(_00653_ ), .CK(clock ), .Q(\EXU.pc_i [10] ), .QN(_10243_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_22 ( .D(_00654_ ), .CK(clock ), .Q(\EXU.pc_i [9] ), .QN(_10242_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_23 ( .D(_00655_ ), .CK(clock ), .Q(\EXU.pc_i [8] ), .QN(_10241_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_24 ( .D(_00656_ ), .CK(clock ), .Q(\EXU.pc_i [7] ), .QN(_10240_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_25 ( .D(_00657_ ), .CK(clock ), .Q(\EXU.pc_i [6] ), .QN(_10239_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_26 ( .D(_00658_ ), .CK(clock ), .Q(\EXU.pc_i [5] ), .QN(_10238_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_27 ( .D(_00659_ ), .CK(clock ), .Q(\EXU.pc_i [4] ), .QN(_10237_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_28 ( .D(_00660_ ), .CK(clock ), .Q(\EXU.pc_i [3] ), .QN(_10236_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_29 ( .D(_00661_ ), .CK(clock ), .Q(\EXU.pc_i [2] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_B_$_MUX__Y_B ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_3 ( .D(_00662_ ), .CK(clock ), .Q(\EXU.pc_i [28] ), .QN(_10235_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_30 ( .D(_00663_ ), .CK(clock ), .Q(\EXU.add_pc_4 [1] ), .QN(_10234_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_31 ( .D(_00664_ ), .CK(clock ), .Q(\EXU.add_pc_4 [0] ), .QN(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_B ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_4 ( .D(_00665_ ), .CK(clock ), .Q(\EXU.pc_i [27] ), .QN(_10233_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_5 ( .D(_00666_ ), .CK(clock ), .Q(\EXU.pc_i [26] ), .QN(_10232_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_6 ( .D(_00667_ ), .CK(clock ), .Q(\EXU.pc_i [25] ), .QN(_10231_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_7 ( .D(_00668_ ), .CK(clock ), .Q(\EXU.pc_i [24] ), .QN(_10230_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_8 ( .D(_00669_ ), .CK(clock ), .Q(\EXU.pc_i [23] ), .QN(_10229_ ) );
DFF_X1 \IDU.pc_o_$_DFFE_PP__Q_9 ( .D(_00670_ ), .CK(clock ), .Q(\EXU.pc_i [22] ), .QN(_10794_ ) );
DFF_X1 \IDU.prevalid_$_DFF_P__Q ( .D(\IFU.updata ), .CK(clock ), .Q(\IDU.prevalid ), .QN(_10228_ ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q ( .D(_00671_ ), .CK(clock ), .Q(\EXU.r1_i [31] ), .QN(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_A_$_MUX__Y_B_$_MUX__B_Y_$_XOR__B_Y_$_OR__A_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_1 ( .D(_00672_ ), .CK(clock ), .Q(\EXU.r1_i [30] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_B_$_MUX__Y_A ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_10 ( .D(_00673_ ), .CK(clock ), .Q(\EXU.r1_i [21] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_11 ( .D(_00674_ ), .CK(clock ), .Q(\EXU.r1_i [20] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_11_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_12 ( .D(_00675_ ), .CK(clock ), .Q(\EXU.r1_i [19] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_12_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_13 ( .D(_00676_ ), .CK(clock ), .Q(\EXU.r1_i [18] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_13_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_14 ( .D(_00677_ ), .CK(clock ), .Q(\EXU.r1_i [17] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_15 ( .D(_00678_ ), .CK(clock ), .Q(\EXU.r1_i [16] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_16 ( .D(_00679_ ), .CK(clock ), .Q(\EXU.r1_i [15] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_16_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_17 ( .D(_00680_ ), .CK(clock ), .Q(\EXU.r1_i [14] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_18 ( .D(_00681_ ), .CK(clock ), .Q(\EXU.r1_i [13] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_19 ( .D(_00682_ ), .CK(clock ), .Q(\EXU.r1_i [12] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_19_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_2 ( .D(_00683_ ), .CK(clock ), .Q(\EXU.r1_i [29] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_2_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_20 ( .D(_00684_ ), .CK(clock ), .Q(\EXU.r1_i [11] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_20_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_21 ( .D(_00685_ ), .CK(clock ), .Q(\EXU.r1_i [10] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_21_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_22 ( .D(_00686_ ), .CK(clock ), .Q(\EXU.r1_i [9] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_22_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_23 ( .D(_00687_ ), .CK(clock ), .Q(\EXU.r1_i [8] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_24 ( .D(_00688_ ), .CK(clock ), .Q(\EXU.r1_i [7] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_24_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_25 ( .D(_00689_ ), .CK(clock ), .Q(\EXU.r1_i [6] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_26 ( .D(_00690_ ), .CK(clock ), .Q(\EXU.r1_i [5] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_26_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_27 ( .D(_00691_ ), .CK(clock ), .Q(\EXU.r1_i [4] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_27_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_28 ( .D(_00692_ ), .CK(clock ), .Q(\EXU.r1_i [3] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_28_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_29 ( .D(_00693_ ), .CK(clock ), .Q(\EXU.r1_i [2] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_22_B_$_XOR__Y_B_$_NOT__Y_A_$_XNOR__Y_B_$_MUX__Y_A ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_3 ( .D(_00694_ ), .CK(clock ), .Q(\EXU.r1_i [28] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_3_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_30 ( .D(_00695_ ), .CK(clock ), .Q(\EXU.r1_i [1] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_B_$_OR__Y_B_$_OR__Y_A_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_31 ( .D(_00696_ ), .CK(clock ), .Q(\EXU.r1_i [0] ), .QN(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_A ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_4 ( .D(_00697_ ), .CK(clock ), .Q(\EXU.r1_i [27] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_4_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_5 ( .D(_00698_ ), .CK(clock ), .Q(\EXU.r1_i [26] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_5_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_6 ( .D(_00699_ ), .CK(clock ), .Q(\EXU.r1_i [25] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_6_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_7 ( .D(_00700_ ), .CK(clock ), .Q(\EXU.r1_i [24] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_8 ( .D(_00701_ ), .CK(clock ), .Q(\EXU.r1_i [23] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_8_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_NAND__Y_B ) );
DFF_X1 \IDU.r1_o_$_DFFE_PP__Q_9 ( .D(_00702_ ), .CK(clock ), .Q(\EXU.r1_i [22] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_OR__Y_A_$_OR__Y_B ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q ( .D(_00703_ ), .CK(clock ), .Q(\EXU.r2_i [31] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_1 ( .D(_00704_ ), .CK(clock ), .Q(\EXU.r2_i [30] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_10 ( .D(_00705_ ), .CK(clock ), .Q(\EXU.r2_i [21] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_11 ( .D(_00706_ ), .CK(clock ), .Q(\EXU.r2_i [20] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_6_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_12 ( .D(_00707_ ), .CK(clock ), .Q(\EXU.r2_i [19] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_7_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_13 ( .D(_00708_ ), .CK(clock ), .Q(\EXU.r2_i [18] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_8_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_14 ( .D(_00709_ ), .CK(clock ), .Q(\EXU.r2_i [17] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_15 ( .D(_00710_ ), .CK(clock ), .Q(\EXU.r2_i [16] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_9_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_16 ( .D(_00711_ ), .CK(clock ), .Q(\EXU.r2_i [15] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_10_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_17 ( .D(_00712_ ), .CK(clock ), .Q(\EXU.r2_i [14] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_11_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_18 ( .D(_00713_ ), .CK(clock ), .Q(\EXU.r2_i [13] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_19 ( .D(_00714_ ), .CK(clock ), .Q(\EXU.r2_i [12] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_12_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_2 ( .D(_00715_ ), .CK(clock ), .Q(\EXU.r2_i [29] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_20 ( .D(_00716_ ), .CK(clock ), .Q(\EXU.r2_i [11] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_21 ( .D(_00717_ ), .CK(clock ), .Q(\EXU.r2_i [10] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_14_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_22 ( .D(_00718_ ), .CK(clock ), .Q(\EXU.r2_i [9] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_15_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_23 ( .D(_00719_ ), .CK(clock ), .Q(\EXU.r2_i [8] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_16_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_24 ( .D(_00720_ ), .CK(clock ), .Q(\EXU.r2_i [7] ), .QN(\LSU.ls_wdata_i_$_MUX__Y_16_A_$_ANDNOT__Y_B ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_25 ( .D(_00721_ ), .CK(clock ), .Q(\EXU.r2_i [6] ), .QN(\LSU.ls_wdata_i_$_MUX__Y_17_A_$_ANDNOT__Y_B ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_26 ( .D(_00722_ ), .CK(clock ), .Q(\EXU.r2_i [5] ), .QN(\LSU.ls_wdata_i_$_MUX__Y_18_A_$_ANDNOT__Y_B ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_27 ( .D(_00723_ ), .CK(clock ), .Q(\EXU.r2_i [4] ), .QN(\LSU.ls_wdata_i_$_MUX__Y_19_A_$_ANDNOT__Y_B ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_28 ( .D(_00724_ ), .CK(clock ), .Q(\EXU.r2_i [3] ), .QN(\LSU.ls_wdata_i_$_MUX__Y_20_A_$_ANDNOT__Y_B ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_29 ( .D(_00725_ ), .CK(clock ), .Q(\EXU.r2_i [2] ), .QN(\LSU.ls_wdata_i_$_MUX__Y_21_A_$_ANDNOT__Y_B ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_3 ( .D(_00726_ ), .CK(clock ), .Q(\EXU.r2_i [28] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_1_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_30 ( .D(_00727_ ), .CK(clock ), .Q(\EXU.r2_i [1] ), .QN(\LSU.ls_wdata_i_$_MUX__Y_22_A_$_ANDNOT__Y_B ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_31 ( .D(_00728_ ), .CK(clock ), .Q(\EXU.r2_i [0] ), .QN(\LSU.ls_wdata_i_$_MUX__Y_23_A_$_ANDNOT__Y_B ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_4 ( .D(_00729_ ), .CK(clock ), .Q(\EXU.r2_i [27] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_2_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_5 ( .D(_00730_ ), .CK(clock ), .Q(\EXU.r2_i [26] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_6 ( .D(_00731_ ), .CK(clock ), .Q(\EXU.r2_i [25] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_7 ( .D(_00732_ ), .CK(clock ), .Q(\EXU.r2_i [24] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_3_B_$_XOR__Y_A_$_ANDNOT__Y_B_$_NOR__Y_A_$_OR__Y_B_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_8 ( .D(_00733_ ), .CK(clock ), .Q(\EXU.r2_i [23] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_4_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.r2_o_$_DFFE_PP__Q_9 ( .D(_00734_ ), .CK(clock ), .Q(\EXU.r2_i [22] ), .QN(\LSU.ls_addr_i_$_ANDNOT__Y_5_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A ) );
DFF_X1 \IDU.rd_o_$_SDFFCE_PN0P__Q ( .D(_00735_ ), .CK(clock ), .Q(\EXU.rd_i [3] ), .QN(_10227_ ) );
DFF_X1 \IDU.rd_o_$_SDFFCE_PN0P__Q_1 ( .D(_00736_ ), .CK(clock ), .Q(\EXU.rd_i [2] ), .QN(_10226_ ) );
DFF_X1 \IDU.rd_o_$_SDFFCE_PN0P__Q_2 ( .D(_00737_ ), .CK(clock ), .Q(\EXU.rd_i [1] ), .QN(_10225_ ) );
DFF_X1 \IDU.rd_o_$_SDFFCE_PN0P__Q_3 ( .D(_00738_ ), .CK(clock ), .Q(\EXU.rd_i [0] ), .QN(_10224_ ) );
DFF_X1 \IDU.state_$_SDFF_PP0__Q ( .D(_00739_ ), .CK(clock ), .Q(\IDU.state ), .QN(\IDU.ls_valid_o_$_DFFE_PP__Q_E_$_OR__Y_B ) );
DFF_X1 \IFU.if_axi_arvalid_o_$_SDFFE_PP0P__Q ( .D(_00740_ ), .CK(clock ), .Q(\ICACHE.m_axi_arvalid ), .QN(\ICACHE.burst_counter_$_DFFE_PP__Q_E_$_ANDNOT__Y_B_$_MUX__Y_A ) );
DFF_X1 \IFU.if_axi_rready_o_$_SDFFE_PP0P__Q ( .D(_00741_ ), .CK(clock ), .Q(\ICACHE.m_axi_rready ), .QN(_10223_ ) );
DFF_X1 \IFU.if_valid_o_$_DFFE_PP__Q ( .D(_00742_ ), .CK(clock ), .Q(\IDU.if_valid_i ), .QN(_10222_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q ( .D(_00743_ ), .CK(clock ), .Q(\IDU.funct7 [6] ), .QN(\IDU.prevalid_$_NAND__B_A_$_ANDNOT__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_1 ( .D(_00744_ ), .CK(clock ), .Q(\IDU.funct7 [5] ), .QN(\IDU.imm_$_NOR__Y_1_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_10 ( .D(_00745_ ), .CK(clock ), .Q(\IDU.immI [1] ), .QN(\IDU.imm_$_NOR__Y_10_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_11 ( .D(_00746_ ), .CK(clock ), .Q(\IDU.immI [0] ), .QN(\IDU.imm_$_NOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_12 ( .D(_00747_ ), .CK(clock ), .Q(\IDU.immJ [19] ), .QN(_10221_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_13 ( .D(_00748_ ), .CK(clock ), .Q(\IDU.immJ [18] ), .QN(_10220_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_14 ( .D(_00749_ ), .CK(clock ), .Q(\IDU.immJ [17] ), .QN(_10219_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_15 ( .D(_00750_ ), .CK(clock ), .Q(\IDU.immJ [16] ), .QN(_10218_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_16 ( .D(_00751_ ), .CK(clock ), .Q(\IDU.immJ [15] ), .QN(_10217_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_17 ( .D(_00752_ ), .CK(clock ), .Q(\IDU.funct3 [2] ), .QN(_10216_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_18 ( .D(_00753_ ), .CK(clock ), .Q(\IDU.funct3 [1] ), .QN(_10215_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_19 ( .D(_00754_ ), .CK(clock ), .Q(\IDU.funct3 [0] ), .QN(_10214_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_2 ( .D(_00755_ ), .CK(clock ), .Q(\IDU.funct7 [4] ), .QN(\IDU.imm_$_NOR__Y_2_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_20 ( .D(_00756_ ), .CK(clock ), .Q(\IDU.immB [4] ), .QN(\IDU.imm_$_NOR__Y_7_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_21 ( .D(_00757_ ), .CK(clock ), .Q(\IDU.immB [3] ), .QN(\IDU.imm_$_NOR__Y_8_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_22 ( .D(_00758_ ), .CK(clock ), .Q(\IDU.immB [2] ), .QN(\IDU.imm_$_NOR__Y_9_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_23 ( .D(_00759_ ), .CK(clock ), .Q(\IDU.immB [1] ), .QN(\IDU.imm_$_NOR__Y_10_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_24 ( .D(_00760_ ), .CK(clock ), .Q(\IDU.immB [11] ), .QN(\IDU.imm_$_NOR__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_25 ( .D(_00761_ ), .CK(clock ), .Q(\IDU.inst_i [6] ), .QN(\IDU.ls_valid_o_$_DFFE_PP__Q_D_$_ANDNOT__Y_B_$_NOR__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_26 ( .D(_00762_ ), .CK(clock ), .Q(\IDU.inst_i [5] ), .QN(_10213_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_27 ( .D(_00763_ ), .CK(clock ), .Q(\IDU.inst_i [4] ), .QN(_10212_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_28 ( .D(_00764_ ), .CK(clock ), .Q(\IDU.inst_i [3] ), .QN(_10211_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_29 ( .D(_00765_ ), .CK(clock ), .Q(\IDU.inst_i [2] ), .QN(_10210_ ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_3 ( .D(_00766_ ), .CK(clock ), .Q(\IDU.funct7 [3] ), .QN(\IDU.imm_$_NOR__Y_3_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_4 ( .D(_00767_ ), .CK(clock ), .Q(\IDU.funct7 [2] ), .QN(\IDU.imm_$_NOR__Y_4_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_5 ( .D(_00768_ ), .CK(clock ), .Q(\IDU.funct7 [1] ), .QN(\IDU.imm_$_NOR__Y_5_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_6 ( .D(_00769_ ), .CK(clock ), .Q(\IDU.funct7 [0] ), .QN(\IDU.imm_$_NOR__Y_6_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_7 ( .D(_00770_ ), .CK(clock ), .Q(\IDU.immI [4] ), .QN(\IDU.imm_$_NOR__Y_7_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_8 ( .D(_00771_ ), .CK(clock ), .Q(\IDU.immI [3] ), .QN(\IDU.imm_$_NOR__Y_8_A_$_MUX__Y_B ) );
DFF_X1 \IFU.inst_o_$_SDFFCE_PN0P__Q_9 ( .D(_00772_ ), .CK(clock ), .Q(\IDU.immI [2] ), .QN(\IDU.imm_$_NOR__Y_9_A_$_MUX__Y_B ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q ( .D(_00773_ ), .CK(clock ), .Q(\BTB.pc_i [31] ), .QN(_10209_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_1 ( .D(_00774_ ), .CK(clock ), .Q(\BTB.pc_i [30] ), .QN(_10208_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_10 ( .D(_00775_ ), .CK(clock ), .Q(\BTB.pc_i [21] ), .QN(_10207_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_11 ( .D(_00776_ ), .CK(clock ), .Q(\BTB.pc_i [20] ), .QN(_10206_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_12 ( .D(_00777_ ), .CK(clock ), .Q(\BTB.pc_i [19] ), .QN(_10205_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_13 ( .D(_00778_ ), .CK(clock ), .Q(\BTB.pc_i [18] ), .QN(_10204_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_14 ( .D(_00779_ ), .CK(clock ), .Q(\BTB.pc_i [17] ), .QN(_10203_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_15 ( .D(_00780_ ), .CK(clock ), .Q(\BTB.pc_i [16] ), .QN(_10202_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_16 ( .D(_00781_ ), .CK(clock ), .Q(\BTB.btag [12] ), .QN(_10201_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_17 ( .D(_00782_ ), .CK(clock ), .Q(\BTB.btag [11] ), .QN(_10200_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_18 ( .D(_00783_ ), .CK(clock ), .Q(\BTB.btag [10] ), .QN(_10199_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_19 ( .D(_00784_ ), .CK(clock ), .Q(\BTB.btag [9] ), .QN(_10198_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_2 ( .D(_00785_ ), .CK(clock ), .Q(\BTB.pc_i [29] ), .QN(_10197_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_20 ( .D(_00786_ ), .CK(clock ), .Q(\BTB.btag [8] ), .QN(_10196_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_21 ( .D(_00787_ ), .CK(clock ), .Q(\BTB.btag [7] ), .QN(_10195_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_22 ( .D(_00788_ ), .CK(clock ), .Q(\BTB.btag [6] ), .QN(_10194_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_23 ( .D(_00789_ ), .CK(clock ), .Q(\BTB.btag [5] ), .QN(_10193_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_24 ( .D(_00790_ ), .CK(clock ), .Q(\BTB.pc_i [1] ), .QN(_10192_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_25 ( .D(_00791_ ), .CK(clock ), .Q(\BTB.pc_i [0] ), .QN(_10191_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_26 ( .D(_00792_ ), .CK(clock ), .Q(\BTB.btag [4] ), .QN(_10190_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_27 ( .D(_00793_ ), .CK(clock ), .Q(\BTB.btag [3] ), .QN(_10189_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_28 ( .D(_00794_ ), .CK(clock ), .Q(\BTB.btag [2] ), .QN(_10188_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_29 ( .D(_00795_ ), .CK(clock ), .Q(\BTB.btag [1] ), .QN(_10187_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_3 ( .D(_00796_ ), .CK(clock ), .Q(\BTB.pc_i [28] ), .QN(_10186_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_30 ( .D(_00797_ ), .CK(clock ), .Q(\BTB.btag [0] ), .QN(\ICACHE.state_$_MUX__S_A ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_31 ( .D(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y ), .CK(clock ), .Q(\BTB.bindex ), .QN(_10795_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D ( .D(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y ), .CK(clock ), .Q(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .QN(_10185_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_4 ( .D(_00798_ ), .CK(clock ), .Q(\BTB.pc_i [27] ), .QN(_10184_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_5 ( .D(_00799_ ), .CK(clock ), .Q(\BTB.pc_i [26] ), .QN(_10183_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_6 ( .D(_00800_ ), .CK(clock ), .Q(\BTB.pc_i [25] ), .QN(_10182_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_7 ( .D(_00801_ ), .CK(clock ), .Q(\BTB.pc_i [24] ), .QN(_10181_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_8 ( .D(_00802_ ), .CK(clock ), .Q(\BTB.pc_i [23] ), .QN(_10180_ ) );
DFF_X1 \IFU.pc_$_DFFE_PP__Q_9 ( .D(_00803_ ), .CK(clock ), .Q(\BTB.pc_i [22] ), .QN(_10179_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q ( .D(_00804_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [31] ), .QN(_10178_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_1 ( .D(_00805_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [30] ), .QN(_10177_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_10 ( .D(_00806_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [21] ), .QN(_10176_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_11 ( .D(_00807_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [20] ), .QN(_10175_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_12 ( .D(_00808_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [19] ), .QN(_10174_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_13 ( .D(_00809_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [18] ), .QN(_10173_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_14 ( .D(_00810_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [17] ), .QN(_10172_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_15 ( .D(_00811_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [16] ), .QN(_10171_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_16 ( .D(_00812_ ), .CK(clock ), .Q(\BTB.btag_pre [12] ), .QN(_10170_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_17 ( .D(_00813_ ), .CK(clock ), .Q(\BTB.btag_pre [11] ), .QN(_10169_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_18 ( .D(_00814_ ), .CK(clock ), .Q(\BTB.btag_pre [10] ), .QN(_10168_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_19 ( .D(_00815_ ), .CK(clock ), .Q(\BTB.btag_pre [9] ), .QN(_10167_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_2 ( .D(_00816_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [29] ), .QN(_10166_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_20 ( .D(_00817_ ), .CK(clock ), .Q(\BTB.btag_pre [8] ), .QN(_10165_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_21 ( .D(_00818_ ), .CK(clock ), .Q(\BTB.btag_pre [7] ), .QN(_10164_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_22 ( .D(_00819_ ), .CK(clock ), .Q(\BTB.btag_pre [6] ), .QN(prepc_$_ANDNOT__Y_6_B_$_XOR__Y_B_$_XOR__Y_B ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_23 ( .D(_00820_ ), .CK(clock ), .Q(\BTB.btag_pre [5] ), .QN(_10163_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_24 ( .D(_00821_ ), .CK(clock ), .Q(\BTB.btag_pre [4] ), .QN(prepc_$_ANDNOT__Y_8_B_$_XOR__Y_B_$_XOR__Y_B ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_25 ( .D(_00822_ ), .CK(clock ), .Q(\BTB.btag_pre [3] ), .QN(_10162_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_26 ( .D(_00823_ ), .CK(clock ), .Q(\BTB.btag_pre [2] ), .QN(prepc_$_ANDNOT__Y_10_B_$_XOR__Y_B_$_XOR__Y_B ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_27 ( .D(_00824_ ), .CK(clock ), .Q(\BTB.btag_pre [1] ), .QN(_10161_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_28 ( .D(_00825_ ), .CK(clock ), .Q(\BTB.btag_pre [0] ), .QN(prepc_$_ANDNOT__Y_12_B_$_XOR__Y_B_$_XOR__Y_B ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_29 ( .D(_00826_ ), .CK(clock ), .Q(\BTB.bindex_pre ), .QN(prepc_$_ANDNOT__Y_13_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_3 ( .D(_00827_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [28] ), .QN(_10160_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_30 ( .D(_00828_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [1] ), .QN(_10159_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_31 ( .D(_00829_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [0] ), .QN(_10158_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_4 ( .D(_00830_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [27] ), .QN(_10157_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_5 ( .D(_00831_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [26] ), .QN(_10156_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_6 ( .D(_00832_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [25] ), .QN(_10155_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_7 ( .D(_00833_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [24] ), .QN(_10154_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_8 ( .D(_00834_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [23] ), .QN(_10153_ ) );
DFF_X1 \IFU.pc_o_$_DFFE_PP__Q_9 ( .D(_00835_ ), .CK(clock ), .Q(\BTB.prepc_tag_i [22] ), .QN(_10152_ ) );
DFF_X1 \IFU.state_$_SDFF_PP0__Q ( .D(_00836_ ), .CK(clock ), .Q(\IFU.state ), .QN(\IFU.state_$_NOT__A_Y ) );
DFF_X1 \LSU.axi_state_$_DFF_P__Q ( .D(\LSU.axi_state_$_DFF_P__Q_D ), .CK(clock ), .Q(\LSU.axi_state [2] ), .QN(\LSU.ls_axi_arvalid_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \LSU.axi_state_$_DFF_P__Q_1 ( .D(\LSU.axi_state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\LSU.axi_state [1] ), .QN(\LSU.ls_axi_wlast_$_DFFE_PP__Q_D ) );
DFF_X1 \LSU.axi_state_$_DFF_P__Q_2 ( .D(\LSU.axi_state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\LSU.axi_state [0] ), .QN(_10151_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q ( .D(_00837_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [31] ), .QN(_10150_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_1 ( .D(_00838_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [30] ), .QN(_10149_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_10 ( .D(_00839_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [21] ), .QN(_10148_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_11 ( .D(_00840_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [20] ), .QN(_10147_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_12 ( .D(_00841_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [19] ), .QN(_10146_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_13 ( .D(_00842_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [18] ), .QN(_10145_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_14 ( .D(_00843_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [17] ), .QN(_10144_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_15 ( .D(_00844_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [16] ), .QN(_10143_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_16 ( .D(_00845_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [15] ), .QN(_10142_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_17 ( .D(_00846_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [14] ), .QN(_10141_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_18 ( .D(_00847_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [13] ), .QN(_10140_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_19 ( .D(_00848_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [12] ), .QN(_10139_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_2 ( .D(_00849_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [29] ), .QN(_10138_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_20 ( .D(_00850_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [11] ), .QN(_10137_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_21 ( .D(_00851_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [10] ), .QN(_10136_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_22 ( .D(_00852_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [9] ), .QN(_10135_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_23 ( .D(_00853_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [8] ), .QN(_10134_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_24 ( .D(_00854_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [7] ), .QN(_10133_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_25 ( .D(_00855_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [6] ), .QN(_10132_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_26 ( .D(_00856_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [5] ), .QN(_10131_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_27 ( .D(_00857_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [4] ), .QN(_10130_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_28 ( .D(_00858_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [3] ), .QN(_10129_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_29 ( .D(_00859_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [2] ), .QN(_10128_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_3 ( .D(_00860_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [28] ), .QN(_10127_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_30 ( .D(_00861_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [1] ), .QN(_10126_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_31 ( .D(_00862_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [0] ), .QN(_10125_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_4 ( .D(_00863_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [27] ), .QN(_10124_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_5 ( .D(_00864_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [26] ), .QN(_10123_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_6 ( .D(_00865_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [25] ), .QN(_10122_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_7 ( .D(_00866_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [24] ), .QN(_10121_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_8 ( .D(_00867_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [23] ), .QN(_10120_ ) );
DFF_X1 \LSU.ls_axi_araddr_$_SDFFCE_PP0P__Q_9 ( .D(_00868_ ), .CK(clock ), .Q(\LSU.ls_axi_araddr [22] ), .QN(_10119_ ) );
DFF_X1 \LSU.ls_axi_arvalid_$_SDFFE_PP0P__Q ( .D(_00869_ ), .CK(clock ), .Q(\LSU.ls_axi_arvalid ), .QN(io_master_arvalid_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q ( .D(_00870_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [31] ), .QN(_10118_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_1 ( .D(_00871_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [30] ), .QN(_10117_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_10 ( .D(_00872_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [21] ), .QN(_10116_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_11 ( .D(_00873_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [20] ), .QN(_10115_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_12 ( .D(_00874_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [19] ), .QN(_10114_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_13 ( .D(_00875_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [18] ), .QN(_10113_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_14 ( .D(_00876_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [17] ), .QN(_10112_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_15 ( .D(_00877_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [16] ), .QN(_10111_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_16 ( .D(_00878_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [15] ), .QN(_10110_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_17 ( .D(_00879_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [14] ), .QN(_10109_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_18 ( .D(_00880_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [13] ), .QN(_10108_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_19 ( .D(_00881_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [12] ), .QN(_10107_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_2 ( .D(_00882_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [29] ), .QN(_10106_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_20 ( .D(_00883_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [11] ), .QN(_10105_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_21 ( .D(_00884_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [10] ), .QN(_10104_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_22 ( .D(_00885_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [9] ), .QN(_10103_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_23 ( .D(_00886_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [8] ), .QN(_10102_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_24 ( .D(_00887_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [7] ), .QN(_10101_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_25 ( .D(_00888_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [6] ), .QN(_10100_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_26 ( .D(_00889_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [5] ), .QN(_10099_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_27 ( .D(_00890_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [4] ), .QN(_10098_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_28 ( .D(_00891_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [3] ), .QN(_10097_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_29 ( .D(_00892_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [2] ), .QN(_10096_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_3 ( .D(_00893_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [28] ), .QN(_10095_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_30 ( .D(_00894_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [1] ), .QN(_10094_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_31 ( .D(_00895_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [0] ), .QN(_10093_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_4 ( .D(_00896_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [27] ), .QN(_10092_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_5 ( .D(_00897_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [26] ), .QN(_10091_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_6 ( .D(_00898_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [25] ), .QN(_10090_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_7 ( .D(_00899_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [24] ), .QN(_10089_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_8 ( .D(_00900_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [23] ), .QN(_10088_ ) );
DFF_X1 \LSU.ls_axi_awaddr_$_SDFFCE_PP0P__Q_9 ( .D(_00901_ ), .CK(clock ), .Q(\LSU.ls_axi_awaddr [22] ), .QN(_10087_ ) );
DFF_X1 \LSU.ls_axi_awvalid_$_SDFFE_PP0P__Q ( .D(_00902_ ), .CK(clock ), .Q(\LSU.ls_axi_awvalid ), .QN(\LSU.ls_axi_awvalid_$_NOT__A_Y ) );
DFF_X1 \LSU.ls_axi_bready_$_SDFFCE_PP0P__Q ( .D(_00903_ ), .CK(clock ), .Q(\LSU.ls_axi_bready ), .QN(_10086_ ) );
DFF_X1 \LSU.ls_axi_rready_$_SDFFCE_PP0P__Q ( .D(_00904_ ), .CK(clock ), .Q(\LSU.ls_axi_rready ), .QN(\LSU.ls_axi_rready_$_NOT__A_Y ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q ( .D(_00905_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [31] ), .QN(_10085_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_1 ( .D(_00906_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [30] ), .QN(_10084_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_10 ( .D(_00907_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [21] ), .QN(_10083_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_11 ( .D(_00908_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [20] ), .QN(_10082_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_12 ( .D(_00909_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [19] ), .QN(_10081_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_13 ( .D(_00910_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [18] ), .QN(_10080_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_14 ( .D(_00911_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [17] ), .QN(_10079_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_15 ( .D(_00912_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [16] ), .QN(_10078_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_16 ( .D(_00913_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [15] ), .QN(_10077_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_17 ( .D(_00914_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [14] ), .QN(_10076_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_18 ( .D(_00915_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [13] ), .QN(_10075_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_19 ( .D(_00916_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [12] ), .QN(_10074_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_2 ( .D(_00917_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [29] ), .QN(_10073_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_20 ( .D(_00918_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [11] ), .QN(_10072_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_21 ( .D(_00919_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [10] ), .QN(_10071_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_22 ( .D(_00920_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [9] ), .QN(_10070_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_23 ( .D(_00921_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [8] ), .QN(_10069_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_24 ( .D(_00922_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [7] ), .QN(_10068_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_25 ( .D(_00923_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [6] ), .QN(_10067_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_26 ( .D(_00924_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [5] ), .QN(_10066_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_27 ( .D(_00925_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [4] ), .QN(_10065_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_28 ( .D(_00926_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [3] ), .QN(_10064_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_29 ( .D(_00927_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [2] ), .QN(_10063_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_3 ( .D(_00928_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [28] ), .QN(_10062_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_30 ( .D(_00929_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [1] ), .QN(_10061_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_31 ( .D(_00930_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [0] ), .QN(_10060_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_4 ( .D(_00931_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [27] ), .QN(_10059_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_5 ( .D(_00932_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [26] ), .QN(_10058_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_6 ( .D(_00933_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [25] ), .QN(_10057_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_7 ( .D(_00934_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [24] ), .QN(_10056_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_8 ( .D(_00935_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [23] ), .QN(_10055_ ) );
DFF_X1 \LSU.ls_axi_wdata_$_SDFFCE_PP0P__Q_9 ( .D(_00936_ ), .CK(clock ), .Q(\LSU.ls_axi_wdata [22] ), .QN(_10054_ ) );
DFF_X1 \LSU.ls_axi_wlast_$_DFFE_PP__Q ( .D(_00937_ ), .CK(clock ), .Q(\LSU.ls_axi_wlast ), .QN(_10053_ ) );
DFF_X1 \LSU.ls_axi_wvalid_$_DFFE_PP__Q ( .D(_00938_ ), .CK(clock ), .Q(\LSU.ls_axi_wvalid ), .QN(\LSU.ls_axi_wvalid_$_NOT__A_Y ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q ( .D(_00939_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [31] ), .QN(_10052_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_1 ( .D(_00940_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [30] ), .QN(_10051_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_10 ( .D(_00941_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [21] ), .QN(_10050_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_11 ( .D(_00942_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [20] ), .QN(_10049_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_12 ( .D(_00943_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [19] ), .QN(_10048_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_13 ( .D(_00944_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [18] ), .QN(_10047_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_14 ( .D(_00945_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [17] ), .QN(_10046_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_15 ( .D(_00946_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [16] ), .QN(_10045_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_16 ( .D(_00947_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [15] ), .QN(_10044_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_17 ( .D(_00948_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [14] ), .QN(_10043_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_18 ( .D(_00949_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [13] ), .QN(_10042_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_19 ( .D(_00950_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [12] ), .QN(_10041_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_2 ( .D(_00951_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [29] ), .QN(_10040_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_20 ( .D(_00952_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [11] ), .QN(_10039_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_21 ( .D(_00953_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [10] ), .QN(_10038_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_22 ( .D(_00954_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [9] ), .QN(_10037_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_23 ( .D(_00955_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [8] ), .QN(_10036_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_24 ( .D(_00956_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [7] ), .QN(_10035_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_25 ( .D(_00957_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [6] ), .QN(_10034_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_26 ( .D(_00958_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [5] ), .QN(_10033_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_27 ( .D(_00959_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [4] ), .QN(_10032_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_28 ( .D(_00960_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [3] ), .QN(_10031_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_29 ( .D(_00961_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [2] ), .QN(_10030_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_3 ( .D(_00962_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [28] ), .QN(_10029_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_30 ( .D(_00963_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [1] ), .QN(_10028_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_31 ( .D(_00964_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [0] ), .QN(_10027_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_4 ( .D(_00965_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [27] ), .QN(_10026_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_5 ( .D(_00966_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [26] ), .QN(_10025_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_6 ( .D(_00967_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [25] ), .QN(_10024_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_7 ( .D(_00968_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [24] ), .QN(_10023_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_8 ( .D(_00969_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [23] ), .QN(_10022_ ) );
DFF_X1 \LSU.ls_rdata_o_$_DFFE_PP__Q_9 ( .D(_00970_ ), .CK(clock ), .Q(\EXU.ls_rdata_i [22] ), .QN(_10796_ ) );
DFF_X1 \LSU.ls_read_done_$_DFF_P__Q ( .D(\LSU.ls_axi_rready_$_ANDNOT__A_Y ), .CK(clock ), .Q(\LSU.ls_read_done ), .QN(_10021_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q ( .D(_00971_ ), .CK(clock ), .Q(\RFU.rf[10][31] ), .QN(_10020_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_1 ( .D(_00972_ ), .CK(clock ), .Q(\RFU.rf[10][30] ), .QN(_10019_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_10 ( .D(_00973_ ), .CK(clock ), .Q(\RFU.rf[10][21] ), .QN(_10018_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_11 ( .D(_00974_ ), .CK(clock ), .Q(\RFU.rf[10][20] ), .QN(_10017_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_12 ( .D(_00975_ ), .CK(clock ), .Q(\RFU.rf[10][19] ), .QN(_10016_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_13 ( .D(_00976_ ), .CK(clock ), .Q(\RFU.rf[10][18] ), .QN(_10015_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_14 ( .D(_00977_ ), .CK(clock ), .Q(\RFU.rf[10][17] ), .QN(_10014_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_15 ( .D(_00978_ ), .CK(clock ), .Q(\RFU.rf[10][16] ), .QN(_10013_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_16 ( .D(_00979_ ), .CK(clock ), .Q(\RFU.rf[10][15] ), .QN(_10012_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_17 ( .D(_00980_ ), .CK(clock ), .Q(\RFU.rf[10][14] ), .QN(_10011_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_18 ( .D(_00981_ ), .CK(clock ), .Q(\RFU.rf[10][13] ), .QN(_10010_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_19 ( .D(_00982_ ), .CK(clock ), .Q(\RFU.rf[10][12] ), .QN(_10009_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_2 ( .D(_00983_ ), .CK(clock ), .Q(\RFU.rf[10][29] ), .QN(_10008_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_20 ( .D(_00984_ ), .CK(clock ), .Q(\RFU.rf[10][11] ), .QN(_10007_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_21 ( .D(_00985_ ), .CK(clock ), .Q(\RFU.rf[10][10] ), .QN(_10006_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_22 ( .D(_00986_ ), .CK(clock ), .Q(\RFU.rf[10][9] ), .QN(_10005_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_23 ( .D(_00987_ ), .CK(clock ), .Q(\RFU.rf[10][8] ), .QN(_10004_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_24 ( .D(_00988_ ), .CK(clock ), .Q(\RFU.rf[10][7] ), .QN(_10003_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_25 ( .D(_00989_ ), .CK(clock ), .Q(\RFU.rf[10][6] ), .QN(_10002_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_26 ( .D(_00990_ ), .CK(clock ), .Q(\RFU.rf[10][5] ), .QN(_10001_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_27 ( .D(_00991_ ), .CK(clock ), .Q(\RFU.rf[10][4] ), .QN(_10000_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_28 ( .D(_00992_ ), .CK(clock ), .Q(\RFU.rf[10][3] ), .QN(_09999_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_29 ( .D(_00993_ ), .CK(clock ), .Q(\RFU.rf[10][2] ), .QN(_09998_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_3 ( .D(_00994_ ), .CK(clock ), .Q(\RFU.rf[10][28] ), .QN(_09997_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_30 ( .D(_00995_ ), .CK(clock ), .Q(\RFU.rf[10][1] ), .QN(_09996_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_31 ( .D(_00996_ ), .CK(clock ), .Q(\RFU.rf[10][0] ), .QN(_09995_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_4 ( .D(_00997_ ), .CK(clock ), .Q(\RFU.rf[10][27] ), .QN(_09994_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_5 ( .D(_00998_ ), .CK(clock ), .Q(\RFU.rf[10][26] ), .QN(_09993_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_6 ( .D(_00999_ ), .CK(clock ), .Q(\RFU.rf[10][25] ), .QN(_09992_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_7 ( .D(_01000_ ), .CK(clock ), .Q(\RFU.rf[10][24] ), .QN(_09991_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_8 ( .D(_01001_ ), .CK(clock ), .Q(\RFU.rf[10][23] ), .QN(_09990_ ) );
DFF_X1 \RFU.rf[10]_$_DFFE_PP__Q_9 ( .D(_01002_ ), .CK(clock ), .Q(\RFU.rf[10][22] ), .QN(_09989_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q ( .D(_01003_ ), .CK(clock ), .Q(\RFU.rf[11][31] ), .QN(_09988_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_1 ( .D(_01004_ ), .CK(clock ), .Q(\RFU.rf[11][30] ), .QN(_09987_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_10 ( .D(_01005_ ), .CK(clock ), .Q(\RFU.rf[11][21] ), .QN(_09986_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_11 ( .D(_01006_ ), .CK(clock ), .Q(\RFU.rf[11][20] ), .QN(_09985_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_12 ( .D(_01007_ ), .CK(clock ), .Q(\RFU.rf[11][19] ), .QN(_09984_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_13 ( .D(_01008_ ), .CK(clock ), .Q(\RFU.rf[11][18] ), .QN(_09983_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_14 ( .D(_01009_ ), .CK(clock ), .Q(\RFU.rf[11][17] ), .QN(_09982_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_15 ( .D(_01010_ ), .CK(clock ), .Q(\RFU.rf[11][16] ), .QN(_09981_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_16 ( .D(_01011_ ), .CK(clock ), .Q(\RFU.rf[11][15] ), .QN(_09980_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_17 ( .D(_01012_ ), .CK(clock ), .Q(\RFU.rf[11][14] ), .QN(_09979_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_18 ( .D(_01013_ ), .CK(clock ), .Q(\RFU.rf[11][13] ), .QN(_09978_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_19 ( .D(_01014_ ), .CK(clock ), .Q(\RFU.rf[11][12] ), .QN(_09977_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_2 ( .D(_01015_ ), .CK(clock ), .Q(\RFU.rf[11][29] ), .QN(_09976_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_20 ( .D(_01016_ ), .CK(clock ), .Q(\RFU.rf[11][11] ), .QN(_09975_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_21 ( .D(_01017_ ), .CK(clock ), .Q(\RFU.rf[11][10] ), .QN(_09974_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_22 ( .D(_01018_ ), .CK(clock ), .Q(\RFU.rf[11][9] ), .QN(_09973_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_23 ( .D(_01019_ ), .CK(clock ), .Q(\RFU.rf[11][8] ), .QN(_09972_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_24 ( .D(_01020_ ), .CK(clock ), .Q(\RFU.rf[11][7] ), .QN(_09971_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_25 ( .D(_01021_ ), .CK(clock ), .Q(\RFU.rf[11][6] ), .QN(_09970_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_26 ( .D(_01022_ ), .CK(clock ), .Q(\RFU.rf[11][5] ), .QN(_09969_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_27 ( .D(_01023_ ), .CK(clock ), .Q(\RFU.rf[11][4] ), .QN(_09968_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_28 ( .D(_01024_ ), .CK(clock ), .Q(\RFU.rf[11][3] ), .QN(_09967_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_29 ( .D(_01025_ ), .CK(clock ), .Q(\RFU.rf[11][2] ), .QN(_09966_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_3 ( .D(_01026_ ), .CK(clock ), .Q(\RFU.rf[11][28] ), .QN(_09965_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_30 ( .D(_01027_ ), .CK(clock ), .Q(\RFU.rf[11][1] ), .QN(_09964_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_31 ( .D(_01028_ ), .CK(clock ), .Q(\RFU.rf[11][0] ), .QN(_09963_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_4 ( .D(_01029_ ), .CK(clock ), .Q(\RFU.rf[11][27] ), .QN(_09962_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_5 ( .D(_01030_ ), .CK(clock ), .Q(\RFU.rf[11][26] ), .QN(_09961_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_6 ( .D(_01031_ ), .CK(clock ), .Q(\RFU.rf[11][25] ), .QN(_09960_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_7 ( .D(_01032_ ), .CK(clock ), .Q(\RFU.rf[11][24] ), .QN(_09959_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_8 ( .D(_01033_ ), .CK(clock ), .Q(\RFU.rf[11][23] ), .QN(_09958_ ) );
DFF_X1 \RFU.rf[11]_$_DFFE_PP__Q_9 ( .D(_01034_ ), .CK(clock ), .Q(\RFU.rf[11][22] ), .QN(_09957_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q ( .D(_01035_ ), .CK(clock ), .Q(\RFU.rf[12][31] ), .QN(_09956_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_1 ( .D(_01036_ ), .CK(clock ), .Q(\RFU.rf[12][30] ), .QN(_09955_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_10 ( .D(_01037_ ), .CK(clock ), .Q(\RFU.rf[12][21] ), .QN(_09954_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_11 ( .D(_01038_ ), .CK(clock ), .Q(\RFU.rf[12][20] ), .QN(_09953_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_12 ( .D(_01039_ ), .CK(clock ), .Q(\RFU.rf[12][19] ), .QN(_09952_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_13 ( .D(_01040_ ), .CK(clock ), .Q(\RFU.rf[12][18] ), .QN(_09951_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_14 ( .D(_01041_ ), .CK(clock ), .Q(\RFU.rf[12][17] ), .QN(_09950_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_15 ( .D(_01042_ ), .CK(clock ), .Q(\RFU.rf[12][16] ), .QN(_09949_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_16 ( .D(_01043_ ), .CK(clock ), .Q(\RFU.rf[12][15] ), .QN(_09948_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_17 ( .D(_01044_ ), .CK(clock ), .Q(\RFU.rf[12][14] ), .QN(_09947_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_18 ( .D(_01045_ ), .CK(clock ), .Q(\RFU.rf[12][13] ), .QN(_09946_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_19 ( .D(_01046_ ), .CK(clock ), .Q(\RFU.rf[12][12] ), .QN(_09945_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_2 ( .D(_01047_ ), .CK(clock ), .Q(\RFU.rf[12][29] ), .QN(_09944_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_20 ( .D(_01048_ ), .CK(clock ), .Q(\RFU.rf[12][11] ), .QN(_09943_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_21 ( .D(_01049_ ), .CK(clock ), .Q(\RFU.rf[12][10] ), .QN(_09942_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_22 ( .D(_01050_ ), .CK(clock ), .Q(\RFU.rf[12][9] ), .QN(_09941_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_23 ( .D(_01051_ ), .CK(clock ), .Q(\RFU.rf[12][8] ), .QN(_09940_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_24 ( .D(_01052_ ), .CK(clock ), .Q(\RFU.rf[12][7] ), .QN(_09939_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_25 ( .D(_01053_ ), .CK(clock ), .Q(\RFU.rf[12][6] ), .QN(_09938_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_26 ( .D(_01054_ ), .CK(clock ), .Q(\RFU.rf[12][5] ), .QN(_09937_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_27 ( .D(_01055_ ), .CK(clock ), .Q(\RFU.rf[12][4] ), .QN(_09936_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_28 ( .D(_01056_ ), .CK(clock ), .Q(\RFU.rf[12][3] ), .QN(_09935_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_29 ( .D(_01057_ ), .CK(clock ), .Q(\RFU.rf[12][2] ), .QN(_09934_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_3 ( .D(_01058_ ), .CK(clock ), .Q(\RFU.rf[12][28] ), .QN(_09933_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_30 ( .D(_01059_ ), .CK(clock ), .Q(\RFU.rf[12][1] ), .QN(_09932_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_31 ( .D(_01060_ ), .CK(clock ), .Q(\RFU.rf[12][0] ), .QN(_09931_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_4 ( .D(_01061_ ), .CK(clock ), .Q(\RFU.rf[12][27] ), .QN(_09930_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_5 ( .D(_01062_ ), .CK(clock ), .Q(\RFU.rf[12][26] ), .QN(_09929_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_6 ( .D(_01063_ ), .CK(clock ), .Q(\RFU.rf[12][25] ), .QN(_09928_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_7 ( .D(_01064_ ), .CK(clock ), .Q(\RFU.rf[12][24] ), .QN(_09927_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_8 ( .D(_01065_ ), .CK(clock ), .Q(\RFU.rf[12][23] ), .QN(_09926_ ) );
DFF_X1 \RFU.rf[12]_$_DFFE_PP__Q_9 ( .D(_01066_ ), .CK(clock ), .Q(\RFU.rf[12][22] ), .QN(_09925_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q ( .D(_01067_ ), .CK(clock ), .Q(\RFU.rf[13][31] ), .QN(_09924_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_1 ( .D(_01068_ ), .CK(clock ), .Q(\RFU.rf[13][30] ), .QN(_09923_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_10 ( .D(_01069_ ), .CK(clock ), .Q(\RFU.rf[13][21] ), .QN(_09922_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_11 ( .D(_01070_ ), .CK(clock ), .Q(\RFU.rf[13][20] ), .QN(_09921_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_12 ( .D(_01071_ ), .CK(clock ), .Q(\RFU.rf[13][19] ), .QN(_09920_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_13 ( .D(_01072_ ), .CK(clock ), .Q(\RFU.rf[13][18] ), .QN(_09919_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_14 ( .D(_01073_ ), .CK(clock ), .Q(\RFU.rf[13][17] ), .QN(_09918_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_15 ( .D(_01074_ ), .CK(clock ), .Q(\RFU.rf[13][16] ), .QN(_09917_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_16 ( .D(_01075_ ), .CK(clock ), .Q(\RFU.rf[13][15] ), .QN(_09916_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_17 ( .D(_01076_ ), .CK(clock ), .Q(\RFU.rf[13][14] ), .QN(_09915_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_18 ( .D(_01077_ ), .CK(clock ), .Q(\RFU.rf[13][13] ), .QN(_09914_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_19 ( .D(_01078_ ), .CK(clock ), .Q(\RFU.rf[13][12] ), .QN(_09913_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_2 ( .D(_01079_ ), .CK(clock ), .Q(\RFU.rf[13][29] ), .QN(_09912_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_20 ( .D(_01080_ ), .CK(clock ), .Q(\RFU.rf[13][11] ), .QN(_09911_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_21 ( .D(_01081_ ), .CK(clock ), .Q(\RFU.rf[13][10] ), .QN(_09910_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_22 ( .D(_01082_ ), .CK(clock ), .Q(\RFU.rf[13][9] ), .QN(_09909_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_23 ( .D(_01083_ ), .CK(clock ), .Q(\RFU.rf[13][8] ), .QN(_09908_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_24 ( .D(_01084_ ), .CK(clock ), .Q(\RFU.rf[13][7] ), .QN(_09907_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_25 ( .D(_01085_ ), .CK(clock ), .Q(\RFU.rf[13][6] ), .QN(_09906_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_26 ( .D(_01086_ ), .CK(clock ), .Q(\RFU.rf[13][5] ), .QN(_09905_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_27 ( .D(_01087_ ), .CK(clock ), .Q(\RFU.rf[13][4] ), .QN(_09904_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_28 ( .D(_01088_ ), .CK(clock ), .Q(\RFU.rf[13][3] ), .QN(_09903_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_29 ( .D(_01089_ ), .CK(clock ), .Q(\RFU.rf[13][2] ), .QN(_09902_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_3 ( .D(_01090_ ), .CK(clock ), .Q(\RFU.rf[13][28] ), .QN(_09901_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_30 ( .D(_01091_ ), .CK(clock ), .Q(\RFU.rf[13][1] ), .QN(_09900_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_31 ( .D(_01092_ ), .CK(clock ), .Q(\RFU.rf[13][0] ), .QN(_09899_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_4 ( .D(_01093_ ), .CK(clock ), .Q(\RFU.rf[13][27] ), .QN(_09898_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_5 ( .D(_01094_ ), .CK(clock ), .Q(\RFU.rf[13][26] ), .QN(_09897_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_6 ( .D(_01095_ ), .CK(clock ), .Q(\RFU.rf[13][25] ), .QN(_09896_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_7 ( .D(_01096_ ), .CK(clock ), .Q(\RFU.rf[13][24] ), .QN(_09895_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_8 ( .D(_01097_ ), .CK(clock ), .Q(\RFU.rf[13][23] ), .QN(_09894_ ) );
DFF_X1 \RFU.rf[13]_$_DFFE_PP__Q_9 ( .D(_01098_ ), .CK(clock ), .Q(\RFU.rf[13][22] ), .QN(_09893_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q ( .D(_01099_ ), .CK(clock ), .Q(\RFU.rf[14][31] ), .QN(_09892_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_1 ( .D(_01100_ ), .CK(clock ), .Q(\RFU.rf[14][30] ), .QN(_09891_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_10 ( .D(_01101_ ), .CK(clock ), .Q(\RFU.rf[14][21] ), .QN(_09890_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_11 ( .D(_01102_ ), .CK(clock ), .Q(\RFU.rf[14][20] ), .QN(_09889_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_12 ( .D(_01103_ ), .CK(clock ), .Q(\RFU.rf[14][19] ), .QN(_09888_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_13 ( .D(_01104_ ), .CK(clock ), .Q(\RFU.rf[14][18] ), .QN(_09887_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_14 ( .D(_01105_ ), .CK(clock ), .Q(\RFU.rf[14][17] ), .QN(_09886_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_15 ( .D(_01106_ ), .CK(clock ), .Q(\RFU.rf[14][16] ), .QN(_09885_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_16 ( .D(_01107_ ), .CK(clock ), .Q(\RFU.rf[14][15] ), .QN(_09884_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_17 ( .D(_01108_ ), .CK(clock ), .Q(\RFU.rf[14][14] ), .QN(_09883_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_18 ( .D(_01109_ ), .CK(clock ), .Q(\RFU.rf[14][13] ), .QN(_09882_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_19 ( .D(_01110_ ), .CK(clock ), .Q(\RFU.rf[14][12] ), .QN(_09881_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_2 ( .D(_01111_ ), .CK(clock ), .Q(\RFU.rf[14][29] ), .QN(_09880_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_20 ( .D(_01112_ ), .CK(clock ), .Q(\RFU.rf[14][11] ), .QN(_09879_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_21 ( .D(_01113_ ), .CK(clock ), .Q(\RFU.rf[14][10] ), .QN(_09878_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_22 ( .D(_01114_ ), .CK(clock ), .Q(\RFU.rf[14][9] ), .QN(_09877_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_23 ( .D(_01115_ ), .CK(clock ), .Q(\RFU.rf[14][8] ), .QN(_09876_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_24 ( .D(_01116_ ), .CK(clock ), .Q(\RFU.rf[14][7] ), .QN(_09875_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_25 ( .D(_01117_ ), .CK(clock ), .Q(\RFU.rf[14][6] ), .QN(_09874_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_26 ( .D(_01118_ ), .CK(clock ), .Q(\RFU.rf[14][5] ), .QN(_09873_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_27 ( .D(_01119_ ), .CK(clock ), .Q(\RFU.rf[14][4] ), .QN(_09872_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_28 ( .D(_01120_ ), .CK(clock ), .Q(\RFU.rf[14][3] ), .QN(_09871_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_29 ( .D(_01121_ ), .CK(clock ), .Q(\RFU.rf[14][2] ), .QN(_09870_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_3 ( .D(_01122_ ), .CK(clock ), .Q(\RFU.rf[14][28] ), .QN(_09869_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_30 ( .D(_01123_ ), .CK(clock ), .Q(\RFU.rf[14][1] ), .QN(_09868_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_31 ( .D(_01124_ ), .CK(clock ), .Q(\RFU.rf[14][0] ), .QN(_09867_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_4 ( .D(_01125_ ), .CK(clock ), .Q(\RFU.rf[14][27] ), .QN(_09866_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_5 ( .D(_01126_ ), .CK(clock ), .Q(\RFU.rf[14][26] ), .QN(_09865_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_6 ( .D(_01127_ ), .CK(clock ), .Q(\RFU.rf[14][25] ), .QN(_09864_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_7 ( .D(_01128_ ), .CK(clock ), .Q(\RFU.rf[14][24] ), .QN(_09863_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_8 ( .D(_01129_ ), .CK(clock ), .Q(\RFU.rf[14][23] ), .QN(_09862_ ) );
DFF_X1 \RFU.rf[14]_$_DFFE_PP__Q_9 ( .D(_01130_ ), .CK(clock ), .Q(\RFU.rf[14][22] ), .QN(_09861_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q ( .D(_01131_ ), .CK(clock ), .Q(\RFU.rf[15][31] ), .QN(_09860_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_1 ( .D(_01132_ ), .CK(clock ), .Q(\RFU.rf[15][30] ), .QN(_09859_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_10 ( .D(_01133_ ), .CK(clock ), .Q(\RFU.rf[15][21] ), .QN(_09858_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_11 ( .D(_01134_ ), .CK(clock ), .Q(\RFU.rf[15][20] ), .QN(_09857_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_12 ( .D(_01135_ ), .CK(clock ), .Q(\RFU.rf[15][19] ), .QN(_09856_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_13 ( .D(_01136_ ), .CK(clock ), .Q(\RFU.rf[15][18] ), .QN(_09855_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_14 ( .D(_01137_ ), .CK(clock ), .Q(\RFU.rf[15][17] ), .QN(_09854_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_15 ( .D(_01138_ ), .CK(clock ), .Q(\RFU.rf[15][16] ), .QN(_09853_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_16 ( .D(_01139_ ), .CK(clock ), .Q(\RFU.rf[15][15] ), .QN(_09852_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_17 ( .D(_01140_ ), .CK(clock ), .Q(\RFU.rf[15][14] ), .QN(_09851_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_18 ( .D(_01141_ ), .CK(clock ), .Q(\RFU.rf[15][13] ), .QN(_09850_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_19 ( .D(_01142_ ), .CK(clock ), .Q(\RFU.rf[15][12] ), .QN(_09849_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_2 ( .D(_01143_ ), .CK(clock ), .Q(\RFU.rf[15][29] ), .QN(_09848_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_20 ( .D(_01144_ ), .CK(clock ), .Q(\RFU.rf[15][11] ), .QN(_09847_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_21 ( .D(_01145_ ), .CK(clock ), .Q(\RFU.rf[15][10] ), .QN(_09846_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_22 ( .D(_01146_ ), .CK(clock ), .Q(\RFU.rf[15][9] ), .QN(_09845_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_23 ( .D(_01147_ ), .CK(clock ), .Q(\RFU.rf[15][8] ), .QN(_09844_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_24 ( .D(_01148_ ), .CK(clock ), .Q(\RFU.rf[15][7] ), .QN(_09843_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_25 ( .D(_01149_ ), .CK(clock ), .Q(\RFU.rf[15][6] ), .QN(_09842_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_26 ( .D(_01150_ ), .CK(clock ), .Q(\RFU.rf[15][5] ), .QN(_09841_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_27 ( .D(_01151_ ), .CK(clock ), .Q(\RFU.rf[15][4] ), .QN(_09840_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_28 ( .D(_01152_ ), .CK(clock ), .Q(\RFU.rf[15][3] ), .QN(_09839_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_29 ( .D(_01153_ ), .CK(clock ), .Q(\RFU.rf[15][2] ), .QN(_09838_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_3 ( .D(_01154_ ), .CK(clock ), .Q(\RFU.rf[15][28] ), .QN(_09837_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_30 ( .D(_01155_ ), .CK(clock ), .Q(\RFU.rf[15][1] ), .QN(_09836_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_31 ( .D(_01156_ ), .CK(clock ), .Q(\RFU.rf[15][0] ), .QN(_09835_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_4 ( .D(_01157_ ), .CK(clock ), .Q(\RFU.rf[15][27] ), .QN(_09834_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_5 ( .D(_01158_ ), .CK(clock ), .Q(\RFU.rf[15][26] ), .QN(_09833_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_6 ( .D(_01159_ ), .CK(clock ), .Q(\RFU.rf[15][25] ), .QN(_09832_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_7 ( .D(_01160_ ), .CK(clock ), .Q(\RFU.rf[15][24] ), .QN(_09831_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_8 ( .D(_01161_ ), .CK(clock ), .Q(\RFU.rf[15][23] ), .QN(_09830_ ) );
DFF_X1 \RFU.rf[15]_$_DFFE_PP__Q_9 ( .D(_01162_ ), .CK(clock ), .Q(\RFU.rf[15][22] ), .QN(_09829_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q ( .D(_01163_ ), .CK(clock ), .Q(\RFU.rf[1][31] ), .QN(_09828_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_1 ( .D(_01164_ ), .CK(clock ), .Q(\RFU.rf[1][30] ), .QN(_09827_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_10 ( .D(_01165_ ), .CK(clock ), .Q(\RFU.rf[1][21] ), .QN(_09826_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_11 ( .D(_01166_ ), .CK(clock ), .Q(\RFU.rf[1][20] ), .QN(_09825_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_12 ( .D(_01167_ ), .CK(clock ), .Q(\RFU.rf[1][19] ), .QN(_09824_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_13 ( .D(_01168_ ), .CK(clock ), .Q(\RFU.rf[1][18] ), .QN(_09823_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_14 ( .D(_01169_ ), .CK(clock ), .Q(\RFU.rf[1][17] ), .QN(_09822_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_15 ( .D(_01170_ ), .CK(clock ), .Q(\RFU.rf[1][16] ), .QN(_09821_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_16 ( .D(_01171_ ), .CK(clock ), .Q(\RFU.rf[1][15] ), .QN(_09820_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_17 ( .D(_01172_ ), .CK(clock ), .Q(\RFU.rf[1][14] ), .QN(_09819_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_18 ( .D(_01173_ ), .CK(clock ), .Q(\RFU.rf[1][13] ), .QN(_09818_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_19 ( .D(_01174_ ), .CK(clock ), .Q(\RFU.rf[1][12] ), .QN(_09817_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_2 ( .D(_01175_ ), .CK(clock ), .Q(\RFU.rf[1][29] ), .QN(_09816_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_20 ( .D(_01176_ ), .CK(clock ), .Q(\RFU.rf[1][11] ), .QN(_09815_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_21 ( .D(_01177_ ), .CK(clock ), .Q(\RFU.rf[1][10] ), .QN(_09814_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_22 ( .D(_01178_ ), .CK(clock ), .Q(\RFU.rf[1][9] ), .QN(_09813_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_23 ( .D(_01179_ ), .CK(clock ), .Q(\RFU.rf[1][8] ), .QN(_09812_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_24 ( .D(_01180_ ), .CK(clock ), .Q(\RFU.rf[1][7] ), .QN(_09811_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_25 ( .D(_01181_ ), .CK(clock ), .Q(\RFU.rf[1][6] ), .QN(_09810_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_26 ( .D(_01182_ ), .CK(clock ), .Q(\RFU.rf[1][5] ), .QN(_09809_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_27 ( .D(_01183_ ), .CK(clock ), .Q(\RFU.rf[1][4] ), .QN(_09808_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_28 ( .D(_01184_ ), .CK(clock ), .Q(\RFU.rf[1][3] ), .QN(_09807_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_29 ( .D(_01185_ ), .CK(clock ), .Q(\RFU.rf[1][2] ), .QN(_09806_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_3 ( .D(_01186_ ), .CK(clock ), .Q(\RFU.rf[1][28] ), .QN(_09805_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_30 ( .D(_01187_ ), .CK(clock ), .Q(\RFU.rf[1][1] ), .QN(_09804_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_31 ( .D(_01188_ ), .CK(clock ), .Q(\RFU.rf[1][0] ), .QN(_09803_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_4 ( .D(_01189_ ), .CK(clock ), .Q(\RFU.rf[1][27] ), .QN(_09802_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_5 ( .D(_01190_ ), .CK(clock ), .Q(\RFU.rf[1][26] ), .QN(_09801_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_6 ( .D(_01191_ ), .CK(clock ), .Q(\RFU.rf[1][25] ), .QN(_09800_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_7 ( .D(_01192_ ), .CK(clock ), .Q(\RFU.rf[1][24] ), .QN(_09799_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_8 ( .D(_01193_ ), .CK(clock ), .Q(\RFU.rf[1][23] ), .QN(_09798_ ) );
DFF_X1 \RFU.rf[1]_$_DFFE_PP__Q_9 ( .D(_01194_ ), .CK(clock ), .Q(\RFU.rf[1][22] ), .QN(_09797_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q ( .D(_01195_ ), .CK(clock ), .Q(\RFU.rf[2][31] ), .QN(_09796_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_1 ( .D(_01196_ ), .CK(clock ), .Q(\RFU.rf[2][30] ), .QN(_09795_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_10 ( .D(_01197_ ), .CK(clock ), .Q(\RFU.rf[2][21] ), .QN(_09794_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_11 ( .D(_01198_ ), .CK(clock ), .Q(\RFU.rf[2][20] ), .QN(_09793_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_12 ( .D(_01199_ ), .CK(clock ), .Q(\RFU.rf[2][19] ), .QN(_09792_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_13 ( .D(_01200_ ), .CK(clock ), .Q(\RFU.rf[2][18] ), .QN(_09791_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_14 ( .D(_01201_ ), .CK(clock ), .Q(\RFU.rf[2][17] ), .QN(_09790_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_15 ( .D(_01202_ ), .CK(clock ), .Q(\RFU.rf[2][16] ), .QN(_09789_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_16 ( .D(_01203_ ), .CK(clock ), .Q(\RFU.rf[2][15] ), .QN(_09788_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_17 ( .D(_01204_ ), .CK(clock ), .Q(\RFU.rf[2][14] ), .QN(_09787_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_18 ( .D(_01205_ ), .CK(clock ), .Q(\RFU.rf[2][13] ), .QN(_09786_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_19 ( .D(_01206_ ), .CK(clock ), .Q(\RFU.rf[2][12] ), .QN(_09785_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_2 ( .D(_01207_ ), .CK(clock ), .Q(\RFU.rf[2][29] ), .QN(_09784_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_20 ( .D(_01208_ ), .CK(clock ), .Q(\RFU.rf[2][11] ), .QN(_09783_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_21 ( .D(_01209_ ), .CK(clock ), .Q(\RFU.rf[2][10] ), .QN(_09782_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_22 ( .D(_01210_ ), .CK(clock ), .Q(\RFU.rf[2][9] ), .QN(_09781_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_23 ( .D(_01211_ ), .CK(clock ), .Q(\RFU.rf[2][8] ), .QN(_09780_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_24 ( .D(_01212_ ), .CK(clock ), .Q(\RFU.rf[2][7] ), .QN(_09779_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_25 ( .D(_01213_ ), .CK(clock ), .Q(\RFU.rf[2][6] ), .QN(_09778_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_26 ( .D(_01214_ ), .CK(clock ), .Q(\RFU.rf[2][5] ), .QN(_09777_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_27 ( .D(_01215_ ), .CK(clock ), .Q(\RFU.rf[2][4] ), .QN(_09776_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_28 ( .D(_01216_ ), .CK(clock ), .Q(\RFU.rf[2][3] ), .QN(_09775_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_29 ( .D(_01217_ ), .CK(clock ), .Q(\RFU.rf[2][2] ), .QN(_09774_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_3 ( .D(_01218_ ), .CK(clock ), .Q(\RFU.rf[2][28] ), .QN(_09773_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_30 ( .D(_01219_ ), .CK(clock ), .Q(\RFU.rf[2][1] ), .QN(_09772_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_31 ( .D(_01220_ ), .CK(clock ), .Q(\RFU.rf[2][0] ), .QN(_09771_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_4 ( .D(_01221_ ), .CK(clock ), .Q(\RFU.rf[2][27] ), .QN(_09770_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_5 ( .D(_01222_ ), .CK(clock ), .Q(\RFU.rf[2][26] ), .QN(_09769_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_6 ( .D(_01223_ ), .CK(clock ), .Q(\RFU.rf[2][25] ), .QN(_09768_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_7 ( .D(_01224_ ), .CK(clock ), .Q(\RFU.rf[2][24] ), .QN(_09767_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_8 ( .D(_01225_ ), .CK(clock ), .Q(\RFU.rf[2][23] ), .QN(_09766_ ) );
DFF_X1 \RFU.rf[2]_$_DFFE_PP__Q_9 ( .D(_01226_ ), .CK(clock ), .Q(\RFU.rf[2][22] ), .QN(_09765_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q ( .D(_01227_ ), .CK(clock ), .Q(\RFU.rf[3][31] ), .QN(_09764_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_1 ( .D(_01228_ ), .CK(clock ), .Q(\RFU.rf[3][30] ), .QN(_09763_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_10 ( .D(_01229_ ), .CK(clock ), .Q(\RFU.rf[3][21] ), .QN(_09762_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_11 ( .D(_01230_ ), .CK(clock ), .Q(\RFU.rf[3][20] ), .QN(_09761_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_12 ( .D(_01231_ ), .CK(clock ), .Q(\RFU.rf[3][19] ), .QN(_09760_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_13 ( .D(_01232_ ), .CK(clock ), .Q(\RFU.rf[3][18] ), .QN(_09759_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_14 ( .D(_01233_ ), .CK(clock ), .Q(\RFU.rf[3][17] ), .QN(_09758_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_15 ( .D(_01234_ ), .CK(clock ), .Q(\RFU.rf[3][16] ), .QN(_09757_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_16 ( .D(_01235_ ), .CK(clock ), .Q(\RFU.rf[3][15] ), .QN(_09756_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_17 ( .D(_01236_ ), .CK(clock ), .Q(\RFU.rf[3][14] ), .QN(_09755_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_18 ( .D(_01237_ ), .CK(clock ), .Q(\RFU.rf[3][13] ), .QN(_09754_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_19 ( .D(_01238_ ), .CK(clock ), .Q(\RFU.rf[3][12] ), .QN(_09753_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_2 ( .D(_01239_ ), .CK(clock ), .Q(\RFU.rf[3][29] ), .QN(_09752_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_20 ( .D(_01240_ ), .CK(clock ), .Q(\RFU.rf[3][11] ), .QN(_09751_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_21 ( .D(_01241_ ), .CK(clock ), .Q(\RFU.rf[3][10] ), .QN(_09750_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_22 ( .D(_01242_ ), .CK(clock ), .Q(\RFU.rf[3][9] ), .QN(_09749_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_23 ( .D(_01243_ ), .CK(clock ), .Q(\RFU.rf[3][8] ), .QN(_09748_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_24 ( .D(_01244_ ), .CK(clock ), .Q(\RFU.rf[3][7] ), .QN(_09747_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_25 ( .D(_01245_ ), .CK(clock ), .Q(\RFU.rf[3][6] ), .QN(_09746_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_26 ( .D(_01246_ ), .CK(clock ), .Q(\RFU.rf[3][5] ), .QN(_09745_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_27 ( .D(_01247_ ), .CK(clock ), .Q(\RFU.rf[3][4] ), .QN(_09744_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_28 ( .D(_01248_ ), .CK(clock ), .Q(\RFU.rf[3][3] ), .QN(_09743_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_29 ( .D(_01249_ ), .CK(clock ), .Q(\RFU.rf[3][2] ), .QN(_09742_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_3 ( .D(_01250_ ), .CK(clock ), .Q(\RFU.rf[3][28] ), .QN(_09741_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_30 ( .D(_01251_ ), .CK(clock ), .Q(\RFU.rf[3][1] ), .QN(_09740_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_31 ( .D(_01252_ ), .CK(clock ), .Q(\RFU.rf[3][0] ), .QN(_09739_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_4 ( .D(_01253_ ), .CK(clock ), .Q(\RFU.rf[3][27] ), .QN(_09738_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_5 ( .D(_01254_ ), .CK(clock ), .Q(\RFU.rf[3][26] ), .QN(_09737_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_6 ( .D(_01255_ ), .CK(clock ), .Q(\RFU.rf[3][25] ), .QN(_09736_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_7 ( .D(_01256_ ), .CK(clock ), .Q(\RFU.rf[3][24] ), .QN(_09735_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_8 ( .D(_01257_ ), .CK(clock ), .Q(\RFU.rf[3][23] ), .QN(_09734_ ) );
DFF_X1 \RFU.rf[3]_$_DFFE_PP__Q_9 ( .D(_01258_ ), .CK(clock ), .Q(\RFU.rf[3][22] ), .QN(_09733_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q ( .D(_01259_ ), .CK(clock ), .Q(\RFU.rf[4][31] ), .QN(_09732_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_1 ( .D(_01260_ ), .CK(clock ), .Q(\RFU.rf[4][30] ), .QN(_09731_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_10 ( .D(_01261_ ), .CK(clock ), .Q(\RFU.rf[4][21] ), .QN(_09730_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_11 ( .D(_01262_ ), .CK(clock ), .Q(\RFU.rf[4][20] ), .QN(_09729_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_12 ( .D(_01263_ ), .CK(clock ), .Q(\RFU.rf[4][19] ), .QN(_09728_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_13 ( .D(_01264_ ), .CK(clock ), .Q(\RFU.rf[4][18] ), .QN(_09727_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_14 ( .D(_01265_ ), .CK(clock ), .Q(\RFU.rf[4][17] ), .QN(_09726_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_15 ( .D(_01266_ ), .CK(clock ), .Q(\RFU.rf[4][16] ), .QN(_09725_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_16 ( .D(_01267_ ), .CK(clock ), .Q(\RFU.rf[4][15] ), .QN(_09724_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_17 ( .D(_01268_ ), .CK(clock ), .Q(\RFU.rf[4][14] ), .QN(_09723_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_18 ( .D(_01269_ ), .CK(clock ), .Q(\RFU.rf[4][13] ), .QN(_09722_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_19 ( .D(_01270_ ), .CK(clock ), .Q(\RFU.rf[4][12] ), .QN(_09721_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_2 ( .D(_01271_ ), .CK(clock ), .Q(\RFU.rf[4][29] ), .QN(_09720_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_20 ( .D(_01272_ ), .CK(clock ), .Q(\RFU.rf[4][11] ), .QN(_09719_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_21 ( .D(_01273_ ), .CK(clock ), .Q(\RFU.rf[4][10] ), .QN(_09718_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_22 ( .D(_01274_ ), .CK(clock ), .Q(\RFU.rf[4][9] ), .QN(_09717_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_23 ( .D(_01275_ ), .CK(clock ), .Q(\RFU.rf[4][8] ), .QN(_09716_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_24 ( .D(_01276_ ), .CK(clock ), .Q(\RFU.rf[4][7] ), .QN(_09715_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_25 ( .D(_01277_ ), .CK(clock ), .Q(\RFU.rf[4][6] ), .QN(_09714_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_26 ( .D(_01278_ ), .CK(clock ), .Q(\RFU.rf[4][5] ), .QN(_09713_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_27 ( .D(_01279_ ), .CK(clock ), .Q(\RFU.rf[4][4] ), .QN(_09712_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_28 ( .D(_01280_ ), .CK(clock ), .Q(\RFU.rf[4][3] ), .QN(_09711_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_29 ( .D(_01281_ ), .CK(clock ), .Q(\RFU.rf[4][2] ), .QN(_09710_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_3 ( .D(_01282_ ), .CK(clock ), .Q(\RFU.rf[4][28] ), .QN(_09709_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_30 ( .D(_01283_ ), .CK(clock ), .Q(\RFU.rf[4][1] ), .QN(_09708_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_31 ( .D(_01284_ ), .CK(clock ), .Q(\RFU.rf[4][0] ), .QN(_09707_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_4 ( .D(_01285_ ), .CK(clock ), .Q(\RFU.rf[4][27] ), .QN(_09706_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_5 ( .D(_01286_ ), .CK(clock ), .Q(\RFU.rf[4][26] ), .QN(_09705_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_6 ( .D(_01287_ ), .CK(clock ), .Q(\RFU.rf[4][25] ), .QN(_09704_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_7 ( .D(_01288_ ), .CK(clock ), .Q(\RFU.rf[4][24] ), .QN(_09703_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_8 ( .D(_01289_ ), .CK(clock ), .Q(\RFU.rf[4][23] ), .QN(_09702_ ) );
DFF_X1 \RFU.rf[4]_$_DFFE_PP__Q_9 ( .D(_01290_ ), .CK(clock ), .Q(\RFU.rf[4][22] ), .QN(_09701_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q ( .D(_01291_ ), .CK(clock ), .Q(\RFU.rf[5][31] ), .QN(_09700_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_1 ( .D(_01292_ ), .CK(clock ), .Q(\RFU.rf[5][30] ), .QN(_09699_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_10 ( .D(_01293_ ), .CK(clock ), .Q(\RFU.rf[5][21] ), .QN(_09698_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_11 ( .D(_01294_ ), .CK(clock ), .Q(\RFU.rf[5][20] ), .QN(_09697_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_12 ( .D(_01295_ ), .CK(clock ), .Q(\RFU.rf[5][19] ), .QN(_09696_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_13 ( .D(_01296_ ), .CK(clock ), .Q(\RFU.rf[5][18] ), .QN(_09695_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_14 ( .D(_01297_ ), .CK(clock ), .Q(\RFU.rf[5][17] ), .QN(_09694_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_15 ( .D(_01298_ ), .CK(clock ), .Q(\RFU.rf[5][16] ), .QN(_09693_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_16 ( .D(_01299_ ), .CK(clock ), .Q(\RFU.rf[5][15] ), .QN(_09692_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_17 ( .D(_01300_ ), .CK(clock ), .Q(\RFU.rf[5][14] ), .QN(_09691_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_18 ( .D(_01301_ ), .CK(clock ), .Q(\RFU.rf[5][13] ), .QN(_09690_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_19 ( .D(_01302_ ), .CK(clock ), .Q(\RFU.rf[5][12] ), .QN(_09689_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_2 ( .D(_01303_ ), .CK(clock ), .Q(\RFU.rf[5][29] ), .QN(_09688_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_20 ( .D(_01304_ ), .CK(clock ), .Q(\RFU.rf[5][11] ), .QN(_09687_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_21 ( .D(_01305_ ), .CK(clock ), .Q(\RFU.rf[5][10] ), .QN(_09686_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_22 ( .D(_01306_ ), .CK(clock ), .Q(\RFU.rf[5][9] ), .QN(_09685_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_23 ( .D(_01307_ ), .CK(clock ), .Q(\RFU.rf[5][8] ), .QN(_09684_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_24 ( .D(_01308_ ), .CK(clock ), .Q(\RFU.rf[5][7] ), .QN(_09683_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_25 ( .D(_01309_ ), .CK(clock ), .Q(\RFU.rf[5][6] ), .QN(_09682_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_26 ( .D(_01310_ ), .CK(clock ), .Q(\RFU.rf[5][5] ), .QN(_09681_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_27 ( .D(_01311_ ), .CK(clock ), .Q(\RFU.rf[5][4] ), .QN(_09680_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_28 ( .D(_01312_ ), .CK(clock ), .Q(\RFU.rf[5][3] ), .QN(_09679_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_29 ( .D(_01313_ ), .CK(clock ), .Q(\RFU.rf[5][2] ), .QN(_09678_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_3 ( .D(_01314_ ), .CK(clock ), .Q(\RFU.rf[5][28] ), .QN(_09677_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_30 ( .D(_01315_ ), .CK(clock ), .Q(\RFU.rf[5][1] ), .QN(_09676_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_31 ( .D(_01316_ ), .CK(clock ), .Q(\RFU.rf[5][0] ), .QN(_09675_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_4 ( .D(_01317_ ), .CK(clock ), .Q(\RFU.rf[5][27] ), .QN(_09674_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_5 ( .D(_01318_ ), .CK(clock ), .Q(\RFU.rf[5][26] ), .QN(_09673_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_6 ( .D(_01319_ ), .CK(clock ), .Q(\RFU.rf[5][25] ), .QN(_09672_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_7 ( .D(_01320_ ), .CK(clock ), .Q(\RFU.rf[5][24] ), .QN(_09671_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_8 ( .D(_01321_ ), .CK(clock ), .Q(\RFU.rf[5][23] ), .QN(_09670_ ) );
DFF_X1 \RFU.rf[5]_$_DFFE_PP__Q_9 ( .D(_01322_ ), .CK(clock ), .Q(\RFU.rf[5][22] ), .QN(_09669_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q ( .D(_01323_ ), .CK(clock ), .Q(\RFU.rf[6][31] ), .QN(_09668_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_1 ( .D(_01324_ ), .CK(clock ), .Q(\RFU.rf[6][30] ), .QN(_09667_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_10 ( .D(_01325_ ), .CK(clock ), .Q(\RFU.rf[6][21] ), .QN(_09666_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_11 ( .D(_01326_ ), .CK(clock ), .Q(\RFU.rf[6][20] ), .QN(_09665_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_12 ( .D(_01327_ ), .CK(clock ), .Q(\RFU.rf[6][19] ), .QN(_09664_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_13 ( .D(_01328_ ), .CK(clock ), .Q(\RFU.rf[6][18] ), .QN(_09663_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_14 ( .D(_01329_ ), .CK(clock ), .Q(\RFU.rf[6][17] ), .QN(_09662_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_15 ( .D(_01330_ ), .CK(clock ), .Q(\RFU.rf[6][16] ), .QN(_09661_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_16 ( .D(_01331_ ), .CK(clock ), .Q(\RFU.rf[6][15] ), .QN(_09660_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_17 ( .D(_01332_ ), .CK(clock ), .Q(\RFU.rf[6][14] ), .QN(_09659_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_18 ( .D(_01333_ ), .CK(clock ), .Q(\RFU.rf[6][13] ), .QN(_09658_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_19 ( .D(_01334_ ), .CK(clock ), .Q(\RFU.rf[6][12] ), .QN(_09657_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_2 ( .D(_01335_ ), .CK(clock ), .Q(\RFU.rf[6][29] ), .QN(_09656_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_20 ( .D(_01336_ ), .CK(clock ), .Q(\RFU.rf[6][11] ), .QN(_09655_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_21 ( .D(_01337_ ), .CK(clock ), .Q(\RFU.rf[6][10] ), .QN(_09654_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_22 ( .D(_01338_ ), .CK(clock ), .Q(\RFU.rf[6][9] ), .QN(_09653_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_23 ( .D(_01339_ ), .CK(clock ), .Q(\RFU.rf[6][8] ), .QN(_09652_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_24 ( .D(_01340_ ), .CK(clock ), .Q(\RFU.rf[6][7] ), .QN(_09651_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_25 ( .D(_01341_ ), .CK(clock ), .Q(\RFU.rf[6][6] ), .QN(_09650_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_26 ( .D(_01342_ ), .CK(clock ), .Q(\RFU.rf[6][5] ), .QN(_09649_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_27 ( .D(_01343_ ), .CK(clock ), .Q(\RFU.rf[6][4] ), .QN(_09648_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_28 ( .D(_01344_ ), .CK(clock ), .Q(\RFU.rf[6][3] ), .QN(_09647_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_29 ( .D(_01345_ ), .CK(clock ), .Q(\RFU.rf[6][2] ), .QN(_09646_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_3 ( .D(_01346_ ), .CK(clock ), .Q(\RFU.rf[6][28] ), .QN(_09645_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_30 ( .D(_01347_ ), .CK(clock ), .Q(\RFU.rf[6][1] ), .QN(_09644_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_31 ( .D(_01348_ ), .CK(clock ), .Q(\RFU.rf[6][0] ), .QN(_09643_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_4 ( .D(_01349_ ), .CK(clock ), .Q(\RFU.rf[6][27] ), .QN(_09642_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_5 ( .D(_01350_ ), .CK(clock ), .Q(\RFU.rf[6][26] ), .QN(_09641_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_6 ( .D(_01351_ ), .CK(clock ), .Q(\RFU.rf[6][25] ), .QN(_09640_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_7 ( .D(_01352_ ), .CK(clock ), .Q(\RFU.rf[6][24] ), .QN(_09639_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_8 ( .D(_01353_ ), .CK(clock ), .Q(\RFU.rf[6][23] ), .QN(_09638_ ) );
DFF_X1 \RFU.rf[6]_$_DFFE_PP__Q_9 ( .D(_01354_ ), .CK(clock ), .Q(\RFU.rf[6][22] ), .QN(_09637_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q ( .D(_01355_ ), .CK(clock ), .Q(\RFU.rf[7][31] ), .QN(_09636_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_1 ( .D(_01356_ ), .CK(clock ), .Q(\RFU.rf[7][30] ), .QN(_09635_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_10 ( .D(_01357_ ), .CK(clock ), .Q(\RFU.rf[7][21] ), .QN(_09634_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_11 ( .D(_01358_ ), .CK(clock ), .Q(\RFU.rf[7][20] ), .QN(_09633_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_12 ( .D(_01359_ ), .CK(clock ), .Q(\RFU.rf[7][19] ), .QN(_09632_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_13 ( .D(_01360_ ), .CK(clock ), .Q(\RFU.rf[7][18] ), .QN(_09631_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_14 ( .D(_01361_ ), .CK(clock ), .Q(\RFU.rf[7][17] ), .QN(_09630_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_15 ( .D(_01362_ ), .CK(clock ), .Q(\RFU.rf[7][16] ), .QN(_09629_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_16 ( .D(_01363_ ), .CK(clock ), .Q(\RFU.rf[7][15] ), .QN(_09628_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_17 ( .D(_01364_ ), .CK(clock ), .Q(\RFU.rf[7][14] ), .QN(_09627_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_18 ( .D(_01365_ ), .CK(clock ), .Q(\RFU.rf[7][13] ), .QN(_09626_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_19 ( .D(_01366_ ), .CK(clock ), .Q(\RFU.rf[7][12] ), .QN(_09625_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_2 ( .D(_01367_ ), .CK(clock ), .Q(\RFU.rf[7][29] ), .QN(_09624_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_20 ( .D(_01368_ ), .CK(clock ), .Q(\RFU.rf[7][11] ), .QN(_09623_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_21 ( .D(_01369_ ), .CK(clock ), .Q(\RFU.rf[7][10] ), .QN(_09622_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_22 ( .D(_01370_ ), .CK(clock ), .Q(\RFU.rf[7][9] ), .QN(_09621_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_23 ( .D(_01371_ ), .CK(clock ), .Q(\RFU.rf[7][8] ), .QN(_09620_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_24 ( .D(_01372_ ), .CK(clock ), .Q(\RFU.rf[7][7] ), .QN(_09619_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_25 ( .D(_01373_ ), .CK(clock ), .Q(\RFU.rf[7][6] ), .QN(_09618_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_26 ( .D(_01374_ ), .CK(clock ), .Q(\RFU.rf[7][5] ), .QN(_09617_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_27 ( .D(_01375_ ), .CK(clock ), .Q(\RFU.rf[7][4] ), .QN(_09616_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_28 ( .D(_01376_ ), .CK(clock ), .Q(\RFU.rf[7][3] ), .QN(_09615_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_29 ( .D(_01377_ ), .CK(clock ), .Q(\RFU.rf[7][2] ), .QN(_09614_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_3 ( .D(_01378_ ), .CK(clock ), .Q(\RFU.rf[7][28] ), .QN(_09613_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_30 ( .D(_01379_ ), .CK(clock ), .Q(\RFU.rf[7][1] ), .QN(_09612_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_31 ( .D(_01380_ ), .CK(clock ), .Q(\RFU.rf[7][0] ), .QN(_09611_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_4 ( .D(_01381_ ), .CK(clock ), .Q(\RFU.rf[7][27] ), .QN(_09610_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_5 ( .D(_01382_ ), .CK(clock ), .Q(\RFU.rf[7][26] ), .QN(_09609_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_6 ( .D(_01383_ ), .CK(clock ), .Q(\RFU.rf[7][25] ), .QN(_09608_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_7 ( .D(_01384_ ), .CK(clock ), .Q(\RFU.rf[7][24] ), .QN(_09607_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_8 ( .D(_01385_ ), .CK(clock ), .Q(\RFU.rf[7][23] ), .QN(_09606_ ) );
DFF_X1 \RFU.rf[7]_$_DFFE_PP__Q_9 ( .D(_01386_ ), .CK(clock ), .Q(\RFU.rf[7][22] ), .QN(_09605_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q ( .D(_01387_ ), .CK(clock ), .Q(\RFU.rf[8][31] ), .QN(_09604_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_1 ( .D(_01388_ ), .CK(clock ), .Q(\RFU.rf[8][30] ), .QN(_09603_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_10 ( .D(_01389_ ), .CK(clock ), .Q(\RFU.rf[8][21] ), .QN(_09602_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_11 ( .D(_01390_ ), .CK(clock ), .Q(\RFU.rf[8][20] ), .QN(_09601_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_12 ( .D(_01391_ ), .CK(clock ), .Q(\RFU.rf[8][19] ), .QN(_09600_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_13 ( .D(_01392_ ), .CK(clock ), .Q(\RFU.rf[8][18] ), .QN(_09599_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_14 ( .D(_01393_ ), .CK(clock ), .Q(\RFU.rf[8][17] ), .QN(_09598_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_15 ( .D(_01394_ ), .CK(clock ), .Q(\RFU.rf[8][16] ), .QN(_09597_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_16 ( .D(_01395_ ), .CK(clock ), .Q(\RFU.rf[8][15] ), .QN(_09596_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_17 ( .D(_01396_ ), .CK(clock ), .Q(\RFU.rf[8][14] ), .QN(_09595_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_18 ( .D(_01397_ ), .CK(clock ), .Q(\RFU.rf[8][13] ), .QN(_09594_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_19 ( .D(_01398_ ), .CK(clock ), .Q(\RFU.rf[8][12] ), .QN(_09593_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_2 ( .D(_01399_ ), .CK(clock ), .Q(\RFU.rf[8][29] ), .QN(_09592_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_20 ( .D(_01400_ ), .CK(clock ), .Q(\RFU.rf[8][11] ), .QN(_09591_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_21 ( .D(_01401_ ), .CK(clock ), .Q(\RFU.rf[8][10] ), .QN(_09590_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_22 ( .D(_01402_ ), .CK(clock ), .Q(\RFU.rf[8][9] ), .QN(_09589_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_23 ( .D(_01403_ ), .CK(clock ), .Q(\RFU.rf[8][8] ), .QN(_09588_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_24 ( .D(_01404_ ), .CK(clock ), .Q(\RFU.rf[8][7] ), .QN(_09587_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_25 ( .D(_01405_ ), .CK(clock ), .Q(\RFU.rf[8][6] ), .QN(_09586_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_26 ( .D(_01406_ ), .CK(clock ), .Q(\RFU.rf[8][5] ), .QN(_09585_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_27 ( .D(_01407_ ), .CK(clock ), .Q(\RFU.rf[8][4] ), .QN(_09584_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_28 ( .D(_01408_ ), .CK(clock ), .Q(\RFU.rf[8][3] ), .QN(_09583_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_29 ( .D(_01409_ ), .CK(clock ), .Q(\RFU.rf[8][2] ), .QN(_09582_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_3 ( .D(_01410_ ), .CK(clock ), .Q(\RFU.rf[8][28] ), .QN(_09581_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_30 ( .D(_01411_ ), .CK(clock ), .Q(\RFU.rf[8][1] ), .QN(_09580_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_31 ( .D(_01412_ ), .CK(clock ), .Q(\RFU.rf[8][0] ), .QN(_09579_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_4 ( .D(_01413_ ), .CK(clock ), .Q(\RFU.rf[8][27] ), .QN(_09578_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_5 ( .D(_01414_ ), .CK(clock ), .Q(\RFU.rf[8][26] ), .QN(_09577_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_6 ( .D(_01415_ ), .CK(clock ), .Q(\RFU.rf[8][25] ), .QN(_09576_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_7 ( .D(_01416_ ), .CK(clock ), .Q(\RFU.rf[8][24] ), .QN(_09575_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_8 ( .D(_01417_ ), .CK(clock ), .Q(\RFU.rf[8][23] ), .QN(_09574_ ) );
DFF_X1 \RFU.rf[8]_$_DFFE_PP__Q_9 ( .D(_01418_ ), .CK(clock ), .Q(\RFU.rf[8][22] ), .QN(_09573_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q ( .D(_01419_ ), .CK(clock ), .Q(\RFU.rf[9][31] ), .QN(_09572_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_1 ( .D(_01420_ ), .CK(clock ), .Q(\RFU.rf[9][30] ), .QN(_09571_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_10 ( .D(_01421_ ), .CK(clock ), .Q(\RFU.rf[9][21] ), .QN(_09570_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_11 ( .D(_01422_ ), .CK(clock ), .Q(\RFU.rf[9][20] ), .QN(_09569_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_12 ( .D(_01423_ ), .CK(clock ), .Q(\RFU.rf[9][19] ), .QN(_09568_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_13 ( .D(_01424_ ), .CK(clock ), .Q(\RFU.rf[9][18] ), .QN(_09567_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_14 ( .D(_01425_ ), .CK(clock ), .Q(\RFU.rf[9][17] ), .QN(_09566_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_15 ( .D(_01426_ ), .CK(clock ), .Q(\RFU.rf[9][16] ), .QN(_09565_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_16 ( .D(_01427_ ), .CK(clock ), .Q(\RFU.rf[9][15] ), .QN(_09564_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_17 ( .D(_01428_ ), .CK(clock ), .Q(\RFU.rf[9][14] ), .QN(_09563_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_18 ( .D(_01429_ ), .CK(clock ), .Q(\RFU.rf[9][13] ), .QN(_09562_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_19 ( .D(_01430_ ), .CK(clock ), .Q(\RFU.rf[9][12] ), .QN(_09561_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_2 ( .D(_01431_ ), .CK(clock ), .Q(\RFU.rf[9][29] ), .QN(_09560_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_20 ( .D(_01432_ ), .CK(clock ), .Q(\RFU.rf[9][11] ), .QN(_09559_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_21 ( .D(_01433_ ), .CK(clock ), .Q(\RFU.rf[9][10] ), .QN(_09558_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_22 ( .D(_01434_ ), .CK(clock ), .Q(\RFU.rf[9][9] ), .QN(_09557_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_23 ( .D(_01435_ ), .CK(clock ), .Q(\RFU.rf[9][8] ), .QN(_09556_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_24 ( .D(_01436_ ), .CK(clock ), .Q(\RFU.rf[9][7] ), .QN(_09555_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_25 ( .D(_01437_ ), .CK(clock ), .Q(\RFU.rf[9][6] ), .QN(_09554_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_26 ( .D(_01438_ ), .CK(clock ), .Q(\RFU.rf[9][5] ), .QN(_09553_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_27 ( .D(_01439_ ), .CK(clock ), .Q(\RFU.rf[9][4] ), .QN(_09552_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_28 ( .D(_01440_ ), .CK(clock ), .Q(\RFU.rf[9][3] ), .QN(_09551_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_29 ( .D(_01441_ ), .CK(clock ), .Q(\RFU.rf[9][2] ), .QN(_09550_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_3 ( .D(_01442_ ), .CK(clock ), .Q(\RFU.rf[9][28] ), .QN(_09549_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_30 ( .D(_01443_ ), .CK(clock ), .Q(\RFU.rf[9][1] ), .QN(_09548_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_31 ( .D(_01444_ ), .CK(clock ), .Q(\RFU.rf[9][0] ), .QN(_09547_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_4 ( .D(_01445_ ), .CK(clock ), .Q(\RFU.rf[9][27] ), .QN(_09546_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_5 ( .D(_01446_ ), .CK(clock ), .Q(\RFU.rf[9][26] ), .QN(_09545_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_6 ( .D(_01447_ ), .CK(clock ), .Q(\RFU.rf[9][25] ), .QN(_09544_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_7 ( .D(_01448_ ), .CK(clock ), .Q(\RFU.rf[9][24] ), .QN(_09543_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_8 ( .D(_01449_ ), .CK(clock ), .Q(\RFU.rf[9][23] ), .QN(_09542_ ) );
DFF_X1 \RFU.rf[9]_$_DFFE_PP__Q_9 ( .D(_01450_ ), .CK(clock ), .Q(\RFU.rf[9][22] ), .QN(_10797_ ) );
DFF_X1 \Xbar.state_$_DFF_P__Q ( .D(\Xbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\Xbar.state [2] ), .QN(_10798_ ) );
DFF_X1 \Xbar.state_$_DFF_P__Q_1 ( .D(\Xbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\Xbar.state [1] ), .QN(_10799_ ) );
DFF_X1 \Xbar.state_$_DFF_P__Q_2 ( .D(\Xbar.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\Xbar.state [0] ), .QN(_09541_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q ( .D(_01451_ ), .CK(clock ), .Q(\EXU.mcause_i [31] ), .QN(_09540_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_1 ( .D(_01452_ ), .CK(clock ), .Q(\EXU.mcause_i [30] ), .QN(_09539_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_10 ( .D(_01453_ ), .CK(clock ), .Q(\EXU.mcause_i [21] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_10_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_11 ( .D(_01454_ ), .CK(clock ), .Q(\EXU.mcause_i [20] ), .QN(_09538_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_12 ( .D(_01455_ ), .CK(clock ), .Q(\EXU.mcause_i [19] ), .QN(_09537_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_13 ( .D(_01456_ ), .CK(clock ), .Q(\EXU.mcause_i [18] ), .QN(_09536_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_14 ( .D(_01457_ ), .CK(clock ), .Q(\EXU.mcause_i [17] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_14_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_15 ( .D(_01458_ ), .CK(clock ), .Q(\EXU.mcause_i [16] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_15_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_16 ( .D(_01459_ ), .CK(clock ), .Q(\EXU.mcause_i [15] ), .QN(_09535_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_17 ( .D(_01460_ ), .CK(clock ), .Q(\EXU.mcause_i [14] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_17_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_18 ( .D(_01461_ ), .CK(clock ), .Q(\EXU.mcause_i [13] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_18_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_19 ( .D(_01462_ ), .CK(clock ), .Q(\EXU.mcause_i [12] ), .QN(_09534_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_2 ( .D(_01463_ ), .CK(clock ), .Q(\EXU.mcause_i [29] ), .QN(_09533_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_20 ( .D(_01464_ ), .CK(clock ), .Q(\EXU.mcause_i [11] ), .QN(_09532_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_21 ( .D(_01465_ ), .CK(clock ), .Q(\EXU.mcause_i [10] ), .QN(_09531_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_22 ( .D(_01466_ ), .CK(clock ), .Q(\EXU.mcause_i [9] ), .QN(_09530_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_23 ( .D(_01467_ ), .CK(clock ), .Q(\EXU.mcause_i [8] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_23_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_24 ( .D(_01468_ ), .CK(clock ), .Q(\EXU.mcause_i [7] ), .QN(_09529_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_25 ( .D(_01469_ ), .CK(clock ), .Q(\EXU.mcause_i [6] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_25_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_26 ( .D(_01470_ ), .CK(clock ), .Q(\EXU.mcause_i [5] ), .QN(_09528_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_27 ( .D(_01471_ ), .CK(clock ), .Q(\EXU.mcause_i [4] ), .QN(_09527_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_28 ( .D(_01472_ ), .CK(clock ), .Q(\EXU.mcause_i [3] ), .QN(_09526_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_29 ( .D(_01473_ ), .CK(clock ), .Q(\EXU.mcause_i [2] ), .QN(_09525_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_3 ( .D(_01474_ ), .CK(clock ), .Q(\EXU.mcause_i [28] ), .QN(_09524_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_30 ( .D(_01475_ ), .CK(clock ), .Q(\EXU.mcause_i [1] ), .QN(_09523_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_31 ( .D(_01476_ ), .CK(clock ), .Q(\EXU.mcause_i [0] ), .QN(\EXU.dnpc_$_MUX__Y_31_B_$_MUX__B_Y_$_MUX__B_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_4 ( .D(_01477_ ), .CK(clock ), .Q(\EXU.mcause_i [27] ), .QN(_09522_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_5 ( .D(_01478_ ), .CK(clock ), .Q(\EXU.mcause_i [26] ), .QN(_09521_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_6 ( .D(_01479_ ), .CK(clock ), .Q(\EXU.mcause_i [25] ), .QN(_09520_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_7 ( .D(_01480_ ), .CK(clock ), .Q(\EXU.mcause_i [24] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_8 ( .D(_01481_ ), .CK(clock ), .Q(\EXU.mcause_i [23] ), .QN(_09519_ ) );
DFF_X1 \mcause_reg.dout_$_SDFFE_PP0P__Q_9 ( .D(_01482_ ), .CK(clock ), .Q(\EXU.mcause_i [22] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q ( .D(_01483_ ), .CK(clock ), .Q(\EXU.mepc_i [31] ), .QN(_09518_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_1 ( .D(_01484_ ), .CK(clock ), .Q(\EXU.mepc_i [30] ), .QN(_09517_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_10 ( .D(_01485_ ), .CK(clock ), .Q(\EXU.mepc_i [21] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_10_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_11 ( .D(_01486_ ), .CK(clock ), .Q(\EXU.mepc_i [20] ), .QN(_09516_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_12 ( .D(_01487_ ), .CK(clock ), .Q(\EXU.mepc_i [19] ), .QN(_09515_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_13 ( .D(_01488_ ), .CK(clock ), .Q(\EXU.mepc_i [18] ), .QN(_09514_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_14 ( .D(_01489_ ), .CK(clock ), .Q(\EXU.mepc_i [17] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_14_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_15 ( .D(_01490_ ), .CK(clock ), .Q(\EXU.mepc_i [16] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_15_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_16 ( .D(_01491_ ), .CK(clock ), .Q(\EXU.mepc_i [15] ), .QN(_09513_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_17 ( .D(_01492_ ), .CK(clock ), .Q(\EXU.mepc_i [14] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_17_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_18 ( .D(_01493_ ), .CK(clock ), .Q(\EXU.mepc_i [13] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_18_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_19 ( .D(_01494_ ), .CK(clock ), .Q(\EXU.mepc_i [12] ), .QN(_09512_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_2 ( .D(_01495_ ), .CK(clock ), .Q(\EXU.mepc_i [29] ), .QN(_09511_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_20 ( .D(_01496_ ), .CK(clock ), .Q(\EXU.mepc_i [11] ), .QN(_09510_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_21 ( .D(_01497_ ), .CK(clock ), .Q(\EXU.mepc_i [10] ), .QN(_09509_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_22 ( .D(_01498_ ), .CK(clock ), .Q(\EXU.mepc_i [9] ), .QN(_09508_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_23 ( .D(_01499_ ), .CK(clock ), .Q(\EXU.mepc_i [8] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_23_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_24 ( .D(_01500_ ), .CK(clock ), .Q(\EXU.mepc_i [7] ), .QN(_09507_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_25 ( .D(_01501_ ), .CK(clock ), .Q(\EXU.mepc_i [6] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_25_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_26 ( .D(_01502_ ), .CK(clock ), .Q(\EXU.mepc_i [5] ), .QN(_09506_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_27 ( .D(_01503_ ), .CK(clock ), .Q(\EXU.mepc_i [4] ), .QN(_09505_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_28 ( .D(_01504_ ), .CK(clock ), .Q(\EXU.mepc_i [3] ), .QN(_09504_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_29 ( .D(_01505_ ), .CK(clock ), .Q(\EXU.mepc_i [2] ), .QN(_09503_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_3 ( .D(_01506_ ), .CK(clock ), .Q(\EXU.mepc_i [28] ), .QN(_09502_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_30 ( .D(_01507_ ), .CK(clock ), .Q(\EXU.mepc_i [1] ), .QN(_09501_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_31 ( .D(_01508_ ), .CK(clock ), .Q(\EXU.mepc_i [0] ), .QN(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_B_$_MUX__A_B ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_4 ( .D(_01509_ ), .CK(clock ), .Q(\EXU.mepc_i [27] ), .QN(_09500_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_5 ( .D(_01510_ ), .CK(clock ), .Q(\EXU.mepc_i [26] ), .QN(_09499_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_6 ( .D(_01511_ ), .CK(clock ), .Q(\EXU.mepc_i [25] ), .QN(_09498_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_7 ( .D(_01512_ ), .CK(clock ), .Q(\EXU.mepc_i [24] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_8 ( .D(_01513_ ), .CK(clock ), .Q(\EXU.mepc_i [23] ), .QN(_09497_ ) );
DFF_X1 \mepc_reg.dout_$_SDFFE_PP0P__Q_9 ( .D(_01514_ ), .CK(clock ), .Q(\EXU.mepc_i [22] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q ( .D(_01515_ ), .CK(clock ), .Q(\EXU.mstatus_i [31] ), .QN(_09496_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_1 ( .D(_01516_ ), .CK(clock ), .Q(\EXU.mstatus_i [30] ), .QN(_09495_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_10 ( .D(_01517_ ), .CK(clock ), .Q(\EXU.mstatus_i [21] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_10_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_11 ( .D(_01518_ ), .CK(clock ), .Q(\EXU.mstatus_i [20] ), .QN(_09494_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_12 ( .D(_01519_ ), .CK(clock ), .Q(\EXU.mstatus_i [19] ), .QN(_09493_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_13 ( .D(_01520_ ), .CK(clock ), .Q(\EXU.mstatus_i [18] ), .QN(_09492_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_14 ( .D(_01521_ ), .CK(clock ), .Q(\EXU.mstatus_i [17] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_14_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_15 ( .D(_01522_ ), .CK(clock ), .Q(\EXU.mstatus_i [16] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_15_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_16 ( .D(_01523_ ), .CK(clock ), .Q(\EXU.mstatus_i [15] ), .QN(_09491_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_17 ( .D(_01524_ ), .CK(clock ), .Q(\EXU.mstatus_i [14] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_17_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_18 ( .D(_01525_ ), .CK(clock ), .Q(\EXU.mstatus_i [13] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_18_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_19 ( .D(_01526_ ), .CK(clock ), .Q(\EXU.mstatus_i [10] ), .QN(_09490_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_2 ( .D(_01527_ ), .CK(clock ), .Q(\EXU.mstatus_i [29] ), .QN(_09489_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_20 ( .D(_01528_ ), .CK(clock ), .Q(\EXU.mstatus_i [9] ), .QN(_09488_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_21 ( .D(_01529_ ), .CK(clock ), .Q(\EXU.mstatus_i [8] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_23_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_22 ( .D(_01530_ ), .CK(clock ), .Q(\EXU.mstatus_i [7] ), .QN(_09487_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_23 ( .D(_01531_ ), .CK(clock ), .Q(\EXU.mstatus_i [6] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_25_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_24 ( .D(_01532_ ), .CK(clock ), .Q(\EXU.mstatus_i [5] ), .QN(_09486_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_25 ( .D(_01533_ ), .CK(clock ), .Q(\EXU.mstatus_i [4] ), .QN(_09485_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_26 ( .D(_01534_ ), .CK(clock ), .Q(\EXU.mstatus_i [3] ), .QN(_09484_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_27 ( .D(_01535_ ), .CK(clock ), .Q(\EXU.mstatus_i [2] ), .QN(_09483_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_28 ( .D(_01536_ ), .CK(clock ), .Q(\EXU.mstatus_i [1] ), .QN(_09482_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_29 ( .D(_01537_ ), .CK(clock ), .Q(\EXU.mstatus_i [0] ), .QN(\EXU.dnpc_$_MUX__Y_31_B_$_MUX__B_Y_$_MUX__B_A_$_MUX__Y_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_3 ( .D(_01538_ ), .CK(clock ), .Q(\EXU.mstatus_i [28] ), .QN(_09481_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_4 ( .D(_01539_ ), .CK(clock ), .Q(\EXU.mstatus_i [27] ), .QN(_09480_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_5 ( .D(_01540_ ), .CK(clock ), .Q(\EXU.mstatus_i [26] ), .QN(_09479_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_6 ( .D(_01541_ ), .CK(clock ), .Q(\EXU.mstatus_i [25] ), .QN(_09478_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_7 ( .D(_01542_ ), .CK(clock ), .Q(\EXU.mstatus_i [24] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_8 ( .D(_01543_ ), .CK(clock ), .Q(\EXU.mstatus_i [23] ), .QN(_09477_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP0P__Q_9 ( .D(_01544_ ), .CK(clock ), .Q(\EXU.mstatus_i [22] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP1P__Q ( .D(_01545_ ), .CK(clock ), .Q(\EXU.mstatus_i [12] ), .QN(_09476_ ) );
DFF_X1 \mstatus_reg.dout_$_SDFFE_PP1P__Q_1 ( .D(_01546_ ), .CK(clock ), .Q(\EXU.mstatus_i [11] ), .QN(_09475_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q ( .D(_01547_ ), .CK(clock ), .Q(\EXU.mtvec_i [31] ), .QN(_09474_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_1 ( .D(_01548_ ), .CK(clock ), .Q(\EXU.mtvec_i [30] ), .QN(_09473_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_10 ( .D(_01549_ ), .CK(clock ), .Q(\EXU.mtvec_i [21] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_10_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_11 ( .D(_01550_ ), .CK(clock ), .Q(\EXU.mtvec_i [20] ), .QN(_09472_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_12 ( .D(_01551_ ), .CK(clock ), .Q(\EXU.mtvec_i [19] ), .QN(_09471_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_13 ( .D(_01552_ ), .CK(clock ), .Q(\EXU.mtvec_i [18] ), .QN(_09470_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_14 ( .D(_01553_ ), .CK(clock ), .Q(\EXU.mtvec_i [17] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_14_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_15 ( .D(_01554_ ), .CK(clock ), .Q(\EXU.mtvec_i [16] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_15_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_16 ( .D(_01555_ ), .CK(clock ), .Q(\EXU.mtvec_i [15] ), .QN(_09469_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_17 ( .D(_01556_ ), .CK(clock ), .Q(\EXU.mtvec_i [14] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_17_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_18 ( .D(_01557_ ), .CK(clock ), .Q(\EXU.mtvec_i [13] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_18_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_19 ( .D(_01558_ ), .CK(clock ), .Q(\EXU.mtvec_i [12] ), .QN(_09468_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_2 ( .D(_01559_ ), .CK(clock ), .Q(\EXU.mtvec_i [29] ), .QN(_09467_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_20 ( .D(_01560_ ), .CK(clock ), .Q(\EXU.mtvec_i [11] ), .QN(_09466_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_21 ( .D(_01561_ ), .CK(clock ), .Q(\EXU.mtvec_i [10] ), .QN(_09465_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_22 ( .D(_01562_ ), .CK(clock ), .Q(\EXU.mtvec_i [9] ), .QN(_09464_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_23 ( .D(_01563_ ), .CK(clock ), .Q(\EXU.mtvec_i [8] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_23_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_24 ( .D(_01564_ ), .CK(clock ), .Q(\EXU.mtvec_i [7] ), .QN(_09463_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_25 ( .D(_01565_ ), .CK(clock ), .Q(\EXU.mtvec_i [6] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_25_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_26 ( .D(_01566_ ), .CK(clock ), .Q(\EXU.mtvec_i [5] ), .QN(_09462_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_27 ( .D(_01567_ ), .CK(clock ), .Q(\EXU.mtvec_i [4] ), .QN(_09461_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_28 ( .D(_01568_ ), .CK(clock ), .Q(\EXU.mtvec_i [3] ), .QN(_09460_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_29 ( .D(_01569_ ), .CK(clock ), .Q(\EXU.mtvec_i [2] ), .QN(_09459_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_3 ( .D(_01570_ ), .CK(clock ), .Q(\EXU.mtvec_i [28] ), .QN(_09458_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_30 ( .D(_01571_ ), .CK(clock ), .Q(\EXU.mtvec_i [1] ), .QN(_09457_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_31 ( .D(_01572_ ), .CK(clock ), .Q(\EXU.mtvec_i [0] ), .QN(\EXU.ls_addr_o_$_ANDNOT__Y_B_$_XOR__Y_A_$_NOR__Y_B_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_A ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_4 ( .D(_01573_ ), .CK(clock ), .Q(\EXU.mtvec_i [27] ), .QN(_09456_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_5 ( .D(_01574_ ), .CK(clock ), .Q(\EXU.mtvec_i [26] ), .QN(_09455_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_6 ( .D(_01575_ ), .CK(clock ), .Q(\EXU.mtvec_i [25] ), .QN(_09454_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_7 ( .D(_01576_ ), .CK(clock ), .Q(\EXU.mtvec_i [24] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_7_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_8 ( .D(_01577_ ), .CK(clock ), .Q(\EXU.mtvec_i [23] ), .QN(_09453_ ) );
DFF_X1 \mtvec_reg.dout_$_SDFFE_PP0P__Q_9 ( .D(_01578_ ), .CK(clock ), .Q(\EXU.mtvec_i [22] ), .QN(\EXU.xrd_o_$_SDFFCE_PP0P__Q_9_D_$_MUX__Y_B_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
BUF_X8 fanout_buf_1 ( .A(\EXU.csrs_wen_o [0] ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(\EXU.csrs_wen_o [1] ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(\EXU.csrs_wen_o [2] ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(\EXU.csrs_wen_o [3] ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\EXU.funct3_i [0] ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\EXU.funct3_i [1] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\EXU.op_i [4] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\EXU.xrd_o_$_SDFFCE_PP0P__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_XOR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\IFU.pc_$_DFFE_PP__Q_31_E_$_MUX__S_Y_$_DFF_P__D_Q ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(io_master_arsize_$_ANDNOT__Y_1_B_$_OR__Y_A_$_OR__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_AND__Y_B_$_OR__Y_B ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(reset ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(reset ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(reset ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(reset ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(reset ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(reset ), .Z(fanout_net_16 ) );

endmodule
