//Generate the verilog at 2025-09-28T22:05:40 by iSTA.
module ysyx_23060229_netlist (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire _08922_ ;
wire _08923_ ;
wire _08924_ ;
wire _08925_ ;
wire _08926_ ;
wire _08927_ ;
wire _08928_ ;
wire _08929_ ;
wire _08930_ ;
wire _08931_ ;
wire _08932_ ;
wire _08933_ ;
wire _08934_ ;
wire _08935_ ;
wire _08936_ ;
wire _08937_ ;
wire _08938_ ;
wire _08939_ ;
wire _08940_ ;
wire _08941_ ;
wire _08942_ ;
wire _08943_ ;
wire _08944_ ;
wire _08945_ ;
wire _08946_ ;
wire _08947_ ;
wire _08948_ ;
wire _08949_ ;
wire _08950_ ;
wire _08951_ ;
wire _08952_ ;
wire _08953_ ;
wire _08954_ ;
wire _08955_ ;
wire _08956_ ;
wire _08957_ ;
wire _08958_ ;
wire _08959_ ;
wire _08960_ ;
wire _08961_ ;
wire _08962_ ;
wire _08963_ ;
wire _08964_ ;
wire _08965_ ;
wire _08966_ ;
wire _08967_ ;
wire _08968_ ;
wire _08969_ ;
wire _08970_ ;
wire _08971_ ;
wire _08972_ ;
wire _08973_ ;
wire _08974_ ;
wire _08975_ ;
wire _08976_ ;
wire _08977_ ;
wire _08978_ ;
wire _08979_ ;
wire _08980_ ;
wire _08981_ ;
wire _08982_ ;
wire _08983_ ;
wire _08984_ ;
wire _08985_ ;
wire _08986_ ;
wire _08987_ ;
wire _08988_ ;
wire _08989_ ;
wire _08990_ ;
wire _08991_ ;
wire _08992_ ;
wire _08993_ ;
wire _08994_ ;
wire _08995_ ;
wire _08996_ ;
wire _08997_ ;
wire _08998_ ;
wire _08999_ ;
wire _09000_ ;
wire _09001_ ;
wire _09002_ ;
wire _09003_ ;
wire _09004_ ;
wire _09005_ ;
wire _09006_ ;
wire _09007_ ;
wire _09008_ ;
wire _09009_ ;
wire _09010_ ;
wire _09011_ ;
wire _09012_ ;
wire EXU_valid_LSU ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire check_assert ;
wire check_quest ;
wire exception_quest_IDU ;
wire excp_written ;
wire fc_disenable ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire loaduse_clear ;
wire \myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ;
wire \myclint.rvalid ;
wire \myclint.state_r_$_NOT__A_Y ;
wire \mycsreg.CSReg[0][0] ;
wire \mycsreg.CSReg[0][10] ;
wire \mycsreg.CSReg[0][11] ;
wire \mycsreg.CSReg[0][12] ;
wire \mycsreg.CSReg[0][13] ;
wire \mycsreg.CSReg[0][14] ;
wire \mycsreg.CSReg[0][15] ;
wire \mycsreg.CSReg[0][16] ;
wire \mycsreg.CSReg[0][17] ;
wire \mycsreg.CSReg[0][18] ;
wire \mycsreg.CSReg[0][19] ;
wire \mycsreg.CSReg[0][1] ;
wire \mycsreg.CSReg[0][20] ;
wire \mycsreg.CSReg[0][21] ;
wire \mycsreg.CSReg[0][22] ;
wire \mycsreg.CSReg[0][23] ;
wire \mycsreg.CSReg[0][24] ;
wire \mycsreg.CSReg[0][25] ;
wire \mycsreg.CSReg[0][26] ;
wire \mycsreg.CSReg[0][27] ;
wire \mycsreg.CSReg[0][28] ;
wire \mycsreg.CSReg[0][29] ;
wire \mycsreg.CSReg[0][2] ;
wire \mycsreg.CSReg[0][30] ;
wire \mycsreg.CSReg[0][31] ;
wire \mycsreg.CSReg[0][3] ;
wire \mycsreg.CSReg[0][4] ;
wire \mycsreg.CSReg[0][5] ;
wire \mycsreg.CSReg[0][6] ;
wire \mycsreg.CSReg[0][7] ;
wire \mycsreg.CSReg[0][8] ;
wire \mycsreg.CSReg[0][9] ;
wire \mycsreg.CSReg[3][0] ;
wire \mycsreg.CSReg[3][10] ;
wire \mycsreg.CSReg[3][11] ;
wire \mycsreg.CSReg[3][12] ;
wire \mycsreg.CSReg[3][13] ;
wire \mycsreg.CSReg[3][14] ;
wire \mycsreg.CSReg[3][15] ;
wire \mycsreg.CSReg[3][16] ;
wire \mycsreg.CSReg[3][17] ;
wire \mycsreg.CSReg[3][18] ;
wire \mycsreg.CSReg[3][19] ;
wire \mycsreg.CSReg[3][1] ;
wire \mycsreg.CSReg[3][20] ;
wire \mycsreg.CSReg[3][21] ;
wire \mycsreg.CSReg[3][22] ;
wire \mycsreg.CSReg[3][23] ;
wire \mycsreg.CSReg[3][24] ;
wire \mycsreg.CSReg[3][25] ;
wire \mycsreg.CSReg[3][26] ;
wire \mycsreg.CSReg[3][27] ;
wire \mycsreg.CSReg[3][28] ;
wire \mycsreg.CSReg[3][29] ;
wire \mycsreg.CSReg[3][2] ;
wire \mycsreg.CSReg[3][30] ;
wire \mycsreg.CSReg[3][31] ;
wire \mycsreg.CSReg[3][3] ;
wire \mycsreg.CSReg[3][4] ;
wire \mycsreg.CSReg[3][5] ;
wire \mycsreg.CSReg[3][6] ;
wire \mycsreg.CSReg[3][7] ;
wire \mycsreg.CSReg[3][8] ;
wire \mycsreg.CSReg[3][9] ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_D ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__B_Y_$_ORNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_10_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_11_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_12_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_13_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_14_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_15_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_16_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_17_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_18_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_19_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_1_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_20_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_21_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_22_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_23_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_24_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_25_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_26_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_27_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_28_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_29_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_2_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_30_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_31_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_3_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_4_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_5_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_6_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_7_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_8_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_9_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_D ;
wire \myec.state_$_SDFFE_PP0P__Q_E ;
wire \myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_10_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_12_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_14_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_15_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_16_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_18_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_19_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_20_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_22_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_23_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_24_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_26_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_27_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_28_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_2_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_30_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_4_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_6_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_7_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_8_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_D ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.state_$_ANDNOT__B_Y ;
wire \myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ;
wire \myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_fencei ;
wire \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ;
wire \myidu.stall_quest_loaduse ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ;
wire \myidu.state_$_DFF_P__Q_1_D ;
wire \myidu.state_$_DFF_P__Q_2_D ;
wire \myidu.state_$_DFF_P__Q_D ;
wire \myidu.typ_$_SDFFE_PP0P__Q_E ;
wire \myifu.check_assert_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[0][0] ;
wire \myifu.myicache.data[0][10] ;
wire \myifu.myicache.data[0][11] ;
wire \myifu.myicache.data[0][12] ;
wire \myifu.myicache.data[0][13] ;
wire \myifu.myicache.data[0][14] ;
wire \myifu.myicache.data[0][15] ;
wire \myifu.myicache.data[0][16] ;
wire \myifu.myicache.data[0][17] ;
wire \myifu.myicache.data[0][18] ;
wire \myifu.myicache.data[0][19] ;
wire \myifu.myicache.data[0][1] ;
wire \myifu.myicache.data[0][20] ;
wire \myifu.myicache.data[0][21] ;
wire \myifu.myicache.data[0][22] ;
wire \myifu.myicache.data[0][23] ;
wire \myifu.myicache.data[0][24] ;
wire \myifu.myicache.data[0][25] ;
wire \myifu.myicache.data[0][26] ;
wire \myifu.myicache.data[0][27] ;
wire \myifu.myicache.data[0][28] ;
wire \myifu.myicache.data[0][29] ;
wire \myifu.myicache.data[0][2] ;
wire \myifu.myicache.data[0][30] ;
wire \myifu.myicache.data[0][31] ;
wire \myifu.myicache.data[0][3] ;
wire \myifu.myicache.data[0][4] ;
wire \myifu.myicache.data[0][5] ;
wire \myifu.myicache.data[0][6] ;
wire \myifu.myicache.data[0][7] ;
wire \myifu.myicache.data[0][8] ;
wire \myifu.myicache.data[0][9] ;
wire \myifu.myicache.data[0]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[1][0] ;
wire \myifu.myicache.data[1][10] ;
wire \myifu.myicache.data[1][11] ;
wire \myifu.myicache.data[1][12] ;
wire \myifu.myicache.data[1][13] ;
wire \myifu.myicache.data[1][14] ;
wire \myifu.myicache.data[1][15] ;
wire \myifu.myicache.data[1][16] ;
wire \myifu.myicache.data[1][17] ;
wire \myifu.myicache.data[1][18] ;
wire \myifu.myicache.data[1][19] ;
wire \myifu.myicache.data[1][1] ;
wire \myifu.myicache.data[1][20] ;
wire \myifu.myicache.data[1][21] ;
wire \myifu.myicache.data[1][22] ;
wire \myifu.myicache.data[1][23] ;
wire \myifu.myicache.data[1][24] ;
wire \myifu.myicache.data[1][25] ;
wire \myifu.myicache.data[1][26] ;
wire \myifu.myicache.data[1][27] ;
wire \myifu.myicache.data[1][28] ;
wire \myifu.myicache.data[1][29] ;
wire \myifu.myicache.data[1][2] ;
wire \myifu.myicache.data[1][30] ;
wire \myifu.myicache.data[1][31] ;
wire \myifu.myicache.data[1][3] ;
wire \myifu.myicache.data[1][4] ;
wire \myifu.myicache.data[1][5] ;
wire \myifu.myicache.data[1][6] ;
wire \myifu.myicache.data[1][7] ;
wire \myifu.myicache.data[1][8] ;
wire \myifu.myicache.data[1][9] ;
wire \myifu.myicache.data[1]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[2][0] ;
wire \myifu.myicache.data[2][10] ;
wire \myifu.myicache.data[2][11] ;
wire \myifu.myicache.data[2][12] ;
wire \myifu.myicache.data[2][13] ;
wire \myifu.myicache.data[2][14] ;
wire \myifu.myicache.data[2][15] ;
wire \myifu.myicache.data[2][16] ;
wire \myifu.myicache.data[2][17] ;
wire \myifu.myicache.data[2][18] ;
wire \myifu.myicache.data[2][19] ;
wire \myifu.myicache.data[2][1] ;
wire \myifu.myicache.data[2][20] ;
wire \myifu.myicache.data[2][21] ;
wire \myifu.myicache.data[2][22] ;
wire \myifu.myicache.data[2][23] ;
wire \myifu.myicache.data[2][24] ;
wire \myifu.myicache.data[2][25] ;
wire \myifu.myicache.data[2][26] ;
wire \myifu.myicache.data[2][27] ;
wire \myifu.myicache.data[2][28] ;
wire \myifu.myicache.data[2][29] ;
wire \myifu.myicache.data[2][2] ;
wire \myifu.myicache.data[2][30] ;
wire \myifu.myicache.data[2][31] ;
wire \myifu.myicache.data[2][3] ;
wire \myifu.myicache.data[2][4] ;
wire \myifu.myicache.data[2][5] ;
wire \myifu.myicache.data[2][6] ;
wire \myifu.myicache.data[2][7] ;
wire \myifu.myicache.data[2][8] ;
wire \myifu.myicache.data[2][9] ;
wire \myifu.myicache.data[2]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[3][0] ;
wire \myifu.myicache.data[3][10] ;
wire \myifu.myicache.data[3][11] ;
wire \myifu.myicache.data[3][12] ;
wire \myifu.myicache.data[3][13] ;
wire \myifu.myicache.data[3][14] ;
wire \myifu.myicache.data[3][15] ;
wire \myifu.myicache.data[3][16] ;
wire \myifu.myicache.data[3][17] ;
wire \myifu.myicache.data[3][18] ;
wire \myifu.myicache.data[3][19] ;
wire \myifu.myicache.data[3][1] ;
wire \myifu.myicache.data[3][20] ;
wire \myifu.myicache.data[3][21] ;
wire \myifu.myicache.data[3][22] ;
wire \myifu.myicache.data[3][23] ;
wire \myifu.myicache.data[3][24] ;
wire \myifu.myicache.data[3][25] ;
wire \myifu.myicache.data[3][26] ;
wire \myifu.myicache.data[3][27] ;
wire \myifu.myicache.data[3][28] ;
wire \myifu.myicache.data[3][29] ;
wire \myifu.myicache.data[3][2] ;
wire \myifu.myicache.data[3][30] ;
wire \myifu.myicache.data[3][31] ;
wire \myifu.myicache.data[3][3] ;
wire \myifu.myicache.data[3][4] ;
wire \myifu.myicache.data[3][5] ;
wire \myifu.myicache.data[3][6] ;
wire \myifu.myicache.data[3][7] ;
wire \myifu.myicache.data[3][8] ;
wire \myifu.myicache.data[3][9] ;
wire \myifu.myicache.data[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[4][0] ;
wire \myifu.myicache.data[4][10] ;
wire \myifu.myicache.data[4][11] ;
wire \myifu.myicache.data[4][12] ;
wire \myifu.myicache.data[4][13] ;
wire \myifu.myicache.data[4][14] ;
wire \myifu.myicache.data[4][15] ;
wire \myifu.myicache.data[4][16] ;
wire \myifu.myicache.data[4][17] ;
wire \myifu.myicache.data[4][18] ;
wire \myifu.myicache.data[4][19] ;
wire \myifu.myicache.data[4][1] ;
wire \myifu.myicache.data[4][20] ;
wire \myifu.myicache.data[4][21] ;
wire \myifu.myicache.data[4][22] ;
wire \myifu.myicache.data[4][23] ;
wire \myifu.myicache.data[4][24] ;
wire \myifu.myicache.data[4][25] ;
wire \myifu.myicache.data[4][26] ;
wire \myifu.myicache.data[4][27] ;
wire \myifu.myicache.data[4][28] ;
wire \myifu.myicache.data[4][29] ;
wire \myifu.myicache.data[4][2] ;
wire \myifu.myicache.data[4][30] ;
wire \myifu.myicache.data[4][31] ;
wire \myifu.myicache.data[4][3] ;
wire \myifu.myicache.data[4][4] ;
wire \myifu.myicache.data[4][5] ;
wire \myifu.myicache.data[4][6] ;
wire \myifu.myicache.data[4][7] ;
wire \myifu.myicache.data[4][8] ;
wire \myifu.myicache.data[4][9] ;
wire \myifu.myicache.data[4]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[5][0] ;
wire \myifu.myicache.data[5][10] ;
wire \myifu.myicache.data[5][11] ;
wire \myifu.myicache.data[5][12] ;
wire \myifu.myicache.data[5][13] ;
wire \myifu.myicache.data[5][14] ;
wire \myifu.myicache.data[5][15] ;
wire \myifu.myicache.data[5][16] ;
wire \myifu.myicache.data[5][17] ;
wire \myifu.myicache.data[5][18] ;
wire \myifu.myicache.data[5][19] ;
wire \myifu.myicache.data[5][1] ;
wire \myifu.myicache.data[5][20] ;
wire \myifu.myicache.data[5][21] ;
wire \myifu.myicache.data[5][22] ;
wire \myifu.myicache.data[5][23] ;
wire \myifu.myicache.data[5][24] ;
wire \myifu.myicache.data[5][25] ;
wire \myifu.myicache.data[5][26] ;
wire \myifu.myicache.data[5][27] ;
wire \myifu.myicache.data[5][28] ;
wire \myifu.myicache.data[5][29] ;
wire \myifu.myicache.data[5][2] ;
wire \myifu.myicache.data[5][30] ;
wire \myifu.myicache.data[5][31] ;
wire \myifu.myicache.data[5][3] ;
wire \myifu.myicache.data[5][4] ;
wire \myifu.myicache.data[5][5] ;
wire \myifu.myicache.data[5][6] ;
wire \myifu.myicache.data[5][7] ;
wire \myifu.myicache.data[5][8] ;
wire \myifu.myicache.data[5][9] ;
wire \myifu.myicache.data[5]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[6][0] ;
wire \myifu.myicache.data[6][10] ;
wire \myifu.myicache.data[6][11] ;
wire \myifu.myicache.data[6][12] ;
wire \myifu.myicache.data[6][13] ;
wire \myifu.myicache.data[6][14] ;
wire \myifu.myicache.data[6][15] ;
wire \myifu.myicache.data[6][16] ;
wire \myifu.myicache.data[6][17] ;
wire \myifu.myicache.data[6][18] ;
wire \myifu.myicache.data[6][19] ;
wire \myifu.myicache.data[6][1] ;
wire \myifu.myicache.data[6][20] ;
wire \myifu.myicache.data[6][21] ;
wire \myifu.myicache.data[6][22] ;
wire \myifu.myicache.data[6][23] ;
wire \myifu.myicache.data[6][24] ;
wire \myifu.myicache.data[6][25] ;
wire \myifu.myicache.data[6][26] ;
wire \myifu.myicache.data[6][27] ;
wire \myifu.myicache.data[6][28] ;
wire \myifu.myicache.data[6][29] ;
wire \myifu.myicache.data[6][2] ;
wire \myifu.myicache.data[6][30] ;
wire \myifu.myicache.data[6][31] ;
wire \myifu.myicache.data[6][3] ;
wire \myifu.myicache.data[6][4] ;
wire \myifu.myicache.data[6][5] ;
wire \myifu.myicache.data[6][6] ;
wire \myifu.myicache.data[6][7] ;
wire \myifu.myicache.data[6][8] ;
wire \myifu.myicache.data[6][9] ;
wire \myifu.myicache.data[6]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[7][0] ;
wire \myifu.myicache.data[7][10] ;
wire \myifu.myicache.data[7][11] ;
wire \myifu.myicache.data[7][12] ;
wire \myifu.myicache.data[7][13] ;
wire \myifu.myicache.data[7][14] ;
wire \myifu.myicache.data[7][15] ;
wire \myifu.myicache.data[7][16] ;
wire \myifu.myicache.data[7][17] ;
wire \myifu.myicache.data[7][18] ;
wire \myifu.myicache.data[7][19] ;
wire \myifu.myicache.data[7][1] ;
wire \myifu.myicache.data[7][20] ;
wire \myifu.myicache.data[7][21] ;
wire \myifu.myicache.data[7][22] ;
wire \myifu.myicache.data[7][23] ;
wire \myifu.myicache.data[7][24] ;
wire \myifu.myicache.data[7][25] ;
wire \myifu.myicache.data[7][26] ;
wire \myifu.myicache.data[7][27] ;
wire \myifu.myicache.data[7][28] ;
wire \myifu.myicache.data[7][29] ;
wire \myifu.myicache.data[7][2] ;
wire \myifu.myicache.data[7][30] ;
wire \myifu.myicache.data[7][31] ;
wire \myifu.myicache.data[7][3] ;
wire \myifu.myicache.data[7][4] ;
wire \myifu.myicache.data[7][5] ;
wire \myifu.myicache.data[7][6] ;
wire \myifu.myicache.data[7][7] ;
wire \myifu.myicache.data[7][8] ;
wire \myifu.myicache.data[7][9] ;
wire \myifu.myicache.data[7]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.tag[0][0] ;
wire \myifu.myicache.tag[0][10] ;
wire \myifu.myicache.tag[0][11] ;
wire \myifu.myicache.tag[0][12] ;
wire \myifu.myicache.tag[0][13] ;
wire \myifu.myicache.tag[0][14] ;
wire \myifu.myicache.tag[0][15] ;
wire \myifu.myicache.tag[0][16] ;
wire \myifu.myicache.tag[0][17] ;
wire \myifu.myicache.tag[0][18] ;
wire \myifu.myicache.tag[0][19] ;
wire \myifu.myicache.tag[0][1] ;
wire \myifu.myicache.tag[0][20] ;
wire \myifu.myicache.tag[0][21] ;
wire \myifu.myicache.tag[0][22] ;
wire \myifu.myicache.tag[0][23] ;
wire \myifu.myicache.tag[0][24] ;
wire \myifu.myicache.tag[0][25] ;
wire \myifu.myicache.tag[0][26] ;
wire \myifu.myicache.tag[0][2] ;
wire \myifu.myicache.tag[0][3] ;
wire \myifu.myicache.tag[0][4] ;
wire \myifu.myicache.tag[0][5] ;
wire \myifu.myicache.tag[0][6] ;
wire \myifu.myicache.tag[0][7] ;
wire \myifu.myicache.tag[0][8] ;
wire \myifu.myicache.tag[0][9] ;
wire \myifu.myicache.tag[0]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.tag[1][0] ;
wire \myifu.myicache.tag[1][10] ;
wire \myifu.myicache.tag[1][11] ;
wire \myifu.myicache.tag[1][12] ;
wire \myifu.myicache.tag[1][13] ;
wire \myifu.myicache.tag[1][14] ;
wire \myifu.myicache.tag[1][15] ;
wire \myifu.myicache.tag[1][16] ;
wire \myifu.myicache.tag[1][17] ;
wire \myifu.myicache.tag[1][18] ;
wire \myifu.myicache.tag[1][19] ;
wire \myifu.myicache.tag[1][1] ;
wire \myifu.myicache.tag[1][20] ;
wire \myifu.myicache.tag[1][21] ;
wire \myifu.myicache.tag[1][22] ;
wire \myifu.myicache.tag[1][23] ;
wire \myifu.myicache.tag[1][24] ;
wire \myifu.myicache.tag[1][25] ;
wire \myifu.myicache.tag[1][26] ;
wire \myifu.myicache.tag[1][2] ;
wire \myifu.myicache.tag[1][3] ;
wire \myifu.myicache.tag[1][4] ;
wire \myifu.myicache.tag[1][5] ;
wire \myifu.myicache.tag[1][6] ;
wire \myifu.myicache.tag[1][7] ;
wire \myifu.myicache.tag[1][8] ;
wire \myifu.myicache.tag[1][9] ;
wire \myifu.myicache.tag[1]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.tag[2][0] ;
wire \myifu.myicache.tag[2][10] ;
wire \myifu.myicache.tag[2][11] ;
wire \myifu.myicache.tag[2][12] ;
wire \myifu.myicache.tag[2][13] ;
wire \myifu.myicache.tag[2][14] ;
wire \myifu.myicache.tag[2][15] ;
wire \myifu.myicache.tag[2][16] ;
wire \myifu.myicache.tag[2][17] ;
wire \myifu.myicache.tag[2][18] ;
wire \myifu.myicache.tag[2][19] ;
wire \myifu.myicache.tag[2][1] ;
wire \myifu.myicache.tag[2][20] ;
wire \myifu.myicache.tag[2][21] ;
wire \myifu.myicache.tag[2][22] ;
wire \myifu.myicache.tag[2][23] ;
wire \myifu.myicache.tag[2][24] ;
wire \myifu.myicache.tag[2][25] ;
wire \myifu.myicache.tag[2][26] ;
wire \myifu.myicache.tag[2][2] ;
wire \myifu.myicache.tag[2][3] ;
wire \myifu.myicache.tag[2][4] ;
wire \myifu.myicache.tag[2][5] ;
wire \myifu.myicache.tag[2][6] ;
wire \myifu.myicache.tag[2][7] ;
wire \myifu.myicache.tag[2][8] ;
wire \myifu.myicache.tag[2][9] ;
wire \myifu.myicache.tag[2]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.tag[3][0] ;
wire \myifu.myicache.tag[3][10] ;
wire \myifu.myicache.tag[3][11] ;
wire \myifu.myicache.tag[3][12] ;
wire \myifu.myicache.tag[3][13] ;
wire \myifu.myicache.tag[3][14] ;
wire \myifu.myicache.tag[3][15] ;
wire \myifu.myicache.tag[3][16] ;
wire \myifu.myicache.tag[3][17] ;
wire \myifu.myicache.tag[3][18] ;
wire \myifu.myicache.tag[3][19] ;
wire \myifu.myicache.tag[3][1] ;
wire \myifu.myicache.tag[3][20] ;
wire \myifu.myicache.tag[3][21] ;
wire \myifu.myicache.tag[3][22] ;
wire \myifu.myicache.tag[3][23] ;
wire \myifu.myicache.tag[3][24] ;
wire \myifu.myicache.tag[3][25] ;
wire \myifu.myicache.tag[3][26] ;
wire \myifu.myicache.tag[3][2] ;
wire \myifu.myicache.tag[3][3] ;
wire \myifu.myicache.tag[3][4] ;
wire \myifu.myicache.tag[3][5] ;
wire \myifu.myicache.tag[3][6] ;
wire \myifu.myicache.tag[3][7] ;
wire \myifu.myicache.tag[3][8] ;
wire \myifu.myicache.tag[3][9] ;
wire \myifu.myicache.tag[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid_data_in ;
wire \myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_E ;
wire \myifu.pc_$_SDFFE_PP1P__Q_E ;
wire \myifu.state_$_DFF_P__Q_1_D ;
wire \myifu.state_$_DFF_P__Q_2_D ;
wire \myifu.state_$_DFF_P__Q_D ;
wire \myifu.tmp_offset_$_SDFFE_PP0P__Q_E ;
wire \myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ;
wire \myifu.to_reset ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ;
wire \myifu.wen_$_ANDNOT__A_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.pc_out_$_SDFFE_PN0P__Q_E ;
wire \mylsu.previous_load_done ;
wire \mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ;
wire \mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_1_D ;
wire \mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ;
wire \mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_2_D ;
wire \mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ;
wire \mylsu.state_$_DFF_P__Q_3_D ;
wire \mylsu.state_$_DFF_P__Q_4_D ;
wire \mylsu.state_$_DFF_P__Q_D ;
wire \mylsu.typ_tmp_$_NOT__A_Y ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_D ;
wire \mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ;
wire \myminixbar.state_$_DFF_P__Q_1_D ;
wire \myminixbar.state_$_DFF_P__Q_D ;
wire \myreg.Reg[0][0] ;
wire \myreg.Reg[0][10] ;
wire \myreg.Reg[0][11] ;
wire \myreg.Reg[0][12] ;
wire \myreg.Reg[0][13] ;
wire \myreg.Reg[0][14] ;
wire \myreg.Reg[0][15] ;
wire \myreg.Reg[0][16] ;
wire \myreg.Reg[0][17] ;
wire \myreg.Reg[0][18] ;
wire \myreg.Reg[0][19] ;
wire \myreg.Reg[0][1] ;
wire \myreg.Reg[0][20] ;
wire \myreg.Reg[0][21] ;
wire \myreg.Reg[0][22] ;
wire \myreg.Reg[0][23] ;
wire \myreg.Reg[0][24] ;
wire \myreg.Reg[0][25] ;
wire \myreg.Reg[0][26] ;
wire \myreg.Reg[0][27] ;
wire \myreg.Reg[0][28] ;
wire \myreg.Reg[0][29] ;
wire \myreg.Reg[0][2] ;
wire \myreg.Reg[0][30] ;
wire \myreg.Reg[0][31] ;
wire \myreg.Reg[0][3] ;
wire \myreg.Reg[0][4] ;
wire \myreg.Reg[0][5] ;
wire \myreg.Reg[0][6] ;
wire \myreg.Reg[0][7] ;
wire \myreg.Reg[0][8] ;
wire \myreg.Reg[0][9] ;
wire \myreg.Reg[10][0] ;
wire \myreg.Reg[10][10] ;
wire \myreg.Reg[10][11] ;
wire \myreg.Reg[10][12] ;
wire \myreg.Reg[10][13] ;
wire \myreg.Reg[10][14] ;
wire \myreg.Reg[10][15] ;
wire \myreg.Reg[10][16] ;
wire \myreg.Reg[10][17] ;
wire \myreg.Reg[10][18] ;
wire \myreg.Reg[10][19] ;
wire \myreg.Reg[10][1] ;
wire \myreg.Reg[10][20] ;
wire \myreg.Reg[10][21] ;
wire \myreg.Reg[10][22] ;
wire \myreg.Reg[10][23] ;
wire \myreg.Reg[10][24] ;
wire \myreg.Reg[10][25] ;
wire \myreg.Reg[10][26] ;
wire \myreg.Reg[10][27] ;
wire \myreg.Reg[10][28] ;
wire \myreg.Reg[10][29] ;
wire \myreg.Reg[10][2] ;
wire \myreg.Reg[10][30] ;
wire \myreg.Reg[10][31] ;
wire \myreg.Reg[10][3] ;
wire \myreg.Reg[10][4] ;
wire \myreg.Reg[10][5] ;
wire \myreg.Reg[10][6] ;
wire \myreg.Reg[10][7] ;
wire \myreg.Reg[10][8] ;
wire \myreg.Reg[10][9] ;
wire \myreg.Reg[11][0] ;
wire \myreg.Reg[11][10] ;
wire \myreg.Reg[11][11] ;
wire \myreg.Reg[11][12] ;
wire \myreg.Reg[11][13] ;
wire \myreg.Reg[11][14] ;
wire \myreg.Reg[11][15] ;
wire \myreg.Reg[11][16] ;
wire \myreg.Reg[11][17] ;
wire \myreg.Reg[11][18] ;
wire \myreg.Reg[11][19] ;
wire \myreg.Reg[11][1] ;
wire \myreg.Reg[11][20] ;
wire \myreg.Reg[11][21] ;
wire \myreg.Reg[11][22] ;
wire \myreg.Reg[11][23] ;
wire \myreg.Reg[11][24] ;
wire \myreg.Reg[11][25] ;
wire \myreg.Reg[11][26] ;
wire \myreg.Reg[11][27] ;
wire \myreg.Reg[11][28] ;
wire \myreg.Reg[11][29] ;
wire \myreg.Reg[11][2] ;
wire \myreg.Reg[11][30] ;
wire \myreg.Reg[11][31] ;
wire \myreg.Reg[11][3] ;
wire \myreg.Reg[11][4] ;
wire \myreg.Reg[11][5] ;
wire \myreg.Reg[11][6] ;
wire \myreg.Reg[11][7] ;
wire \myreg.Reg[11][8] ;
wire \myreg.Reg[11][9] ;
wire \myreg.Reg[12][0] ;
wire \myreg.Reg[12][10] ;
wire \myreg.Reg[12][11] ;
wire \myreg.Reg[12][12] ;
wire \myreg.Reg[12][13] ;
wire \myreg.Reg[12][14] ;
wire \myreg.Reg[12][15] ;
wire \myreg.Reg[12][16] ;
wire \myreg.Reg[12][17] ;
wire \myreg.Reg[12][18] ;
wire \myreg.Reg[12][19] ;
wire \myreg.Reg[12][1] ;
wire \myreg.Reg[12][20] ;
wire \myreg.Reg[12][21] ;
wire \myreg.Reg[12][22] ;
wire \myreg.Reg[12][23] ;
wire \myreg.Reg[12][24] ;
wire \myreg.Reg[12][25] ;
wire \myreg.Reg[12][26] ;
wire \myreg.Reg[12][27] ;
wire \myreg.Reg[12][28] ;
wire \myreg.Reg[12][29] ;
wire \myreg.Reg[12][2] ;
wire \myreg.Reg[12][30] ;
wire \myreg.Reg[12][31] ;
wire \myreg.Reg[12][3] ;
wire \myreg.Reg[12][4] ;
wire \myreg.Reg[12][5] ;
wire \myreg.Reg[12][6] ;
wire \myreg.Reg[12][7] ;
wire \myreg.Reg[12][8] ;
wire \myreg.Reg[12][9] ;
wire \myreg.Reg[13][0] ;
wire \myreg.Reg[13][10] ;
wire \myreg.Reg[13][11] ;
wire \myreg.Reg[13][12] ;
wire \myreg.Reg[13][13] ;
wire \myreg.Reg[13][14] ;
wire \myreg.Reg[13][15] ;
wire \myreg.Reg[13][16] ;
wire \myreg.Reg[13][17] ;
wire \myreg.Reg[13][18] ;
wire \myreg.Reg[13][19] ;
wire \myreg.Reg[13][1] ;
wire \myreg.Reg[13][20] ;
wire \myreg.Reg[13][21] ;
wire \myreg.Reg[13][22] ;
wire \myreg.Reg[13][23] ;
wire \myreg.Reg[13][24] ;
wire \myreg.Reg[13][25] ;
wire \myreg.Reg[13][26] ;
wire \myreg.Reg[13][27] ;
wire \myreg.Reg[13][28] ;
wire \myreg.Reg[13][29] ;
wire \myreg.Reg[13][2] ;
wire \myreg.Reg[13][30] ;
wire \myreg.Reg[13][31] ;
wire \myreg.Reg[13][3] ;
wire \myreg.Reg[13][4] ;
wire \myreg.Reg[13][5] ;
wire \myreg.Reg[13][6] ;
wire \myreg.Reg[13][7] ;
wire \myreg.Reg[13][8] ;
wire \myreg.Reg[13][9] ;
wire \myreg.Reg[14][0] ;
wire \myreg.Reg[14][10] ;
wire \myreg.Reg[14][11] ;
wire \myreg.Reg[14][12] ;
wire \myreg.Reg[14][13] ;
wire \myreg.Reg[14][14] ;
wire \myreg.Reg[14][15] ;
wire \myreg.Reg[14][16] ;
wire \myreg.Reg[14][17] ;
wire \myreg.Reg[14][18] ;
wire \myreg.Reg[14][19] ;
wire \myreg.Reg[14][1] ;
wire \myreg.Reg[14][20] ;
wire \myreg.Reg[14][21] ;
wire \myreg.Reg[14][22] ;
wire \myreg.Reg[14][23] ;
wire \myreg.Reg[14][24] ;
wire \myreg.Reg[14][25] ;
wire \myreg.Reg[14][26] ;
wire \myreg.Reg[14][27] ;
wire \myreg.Reg[14][28] ;
wire \myreg.Reg[14][29] ;
wire \myreg.Reg[14][2] ;
wire \myreg.Reg[14][30] ;
wire \myreg.Reg[14][31] ;
wire \myreg.Reg[14][3] ;
wire \myreg.Reg[14][4] ;
wire \myreg.Reg[14][5] ;
wire \myreg.Reg[14][6] ;
wire \myreg.Reg[14][7] ;
wire \myreg.Reg[14][8] ;
wire \myreg.Reg[14][9] ;
wire \myreg.Reg[15][0] ;
wire \myreg.Reg[15][10] ;
wire \myreg.Reg[15][11] ;
wire \myreg.Reg[15][12] ;
wire \myreg.Reg[15][13] ;
wire \myreg.Reg[15][14] ;
wire \myreg.Reg[15][15] ;
wire \myreg.Reg[15][16] ;
wire \myreg.Reg[15][17] ;
wire \myreg.Reg[15][18] ;
wire \myreg.Reg[15][19] ;
wire \myreg.Reg[15][1] ;
wire \myreg.Reg[15][20] ;
wire \myreg.Reg[15][21] ;
wire \myreg.Reg[15][22] ;
wire \myreg.Reg[15][23] ;
wire \myreg.Reg[15][24] ;
wire \myreg.Reg[15][25] ;
wire \myreg.Reg[15][26] ;
wire \myreg.Reg[15][27] ;
wire \myreg.Reg[15][28] ;
wire \myreg.Reg[15][29] ;
wire \myreg.Reg[15][2] ;
wire \myreg.Reg[15][30] ;
wire \myreg.Reg[15][31] ;
wire \myreg.Reg[15][3] ;
wire \myreg.Reg[15][4] ;
wire \myreg.Reg[15][5] ;
wire \myreg.Reg[15][6] ;
wire \myreg.Reg[15][7] ;
wire \myreg.Reg[15][8] ;
wire \myreg.Reg[15][9] ;
wire \myreg.Reg[1][0] ;
wire \myreg.Reg[1][10] ;
wire \myreg.Reg[1][11] ;
wire \myreg.Reg[1][12] ;
wire \myreg.Reg[1][13] ;
wire \myreg.Reg[1][14] ;
wire \myreg.Reg[1][15] ;
wire \myreg.Reg[1][16] ;
wire \myreg.Reg[1][17] ;
wire \myreg.Reg[1][18] ;
wire \myreg.Reg[1][19] ;
wire \myreg.Reg[1][1] ;
wire \myreg.Reg[1][20] ;
wire \myreg.Reg[1][21] ;
wire \myreg.Reg[1][22] ;
wire \myreg.Reg[1][23] ;
wire \myreg.Reg[1][24] ;
wire \myreg.Reg[1][25] ;
wire \myreg.Reg[1][26] ;
wire \myreg.Reg[1][27] ;
wire \myreg.Reg[1][28] ;
wire \myreg.Reg[1][29] ;
wire \myreg.Reg[1][2] ;
wire \myreg.Reg[1][30] ;
wire \myreg.Reg[1][31] ;
wire \myreg.Reg[1][3] ;
wire \myreg.Reg[1][4] ;
wire \myreg.Reg[1][5] ;
wire \myreg.Reg[1][6] ;
wire \myreg.Reg[1][7] ;
wire \myreg.Reg[1][8] ;
wire \myreg.Reg[1][9] ;
wire \myreg.Reg[2][0] ;
wire \myreg.Reg[2][10] ;
wire \myreg.Reg[2][11] ;
wire \myreg.Reg[2][12] ;
wire \myreg.Reg[2][13] ;
wire \myreg.Reg[2][14] ;
wire \myreg.Reg[2][15] ;
wire \myreg.Reg[2][16] ;
wire \myreg.Reg[2][17] ;
wire \myreg.Reg[2][18] ;
wire \myreg.Reg[2][19] ;
wire \myreg.Reg[2][1] ;
wire \myreg.Reg[2][20] ;
wire \myreg.Reg[2][21] ;
wire \myreg.Reg[2][22] ;
wire \myreg.Reg[2][23] ;
wire \myreg.Reg[2][24] ;
wire \myreg.Reg[2][25] ;
wire \myreg.Reg[2][26] ;
wire \myreg.Reg[2][27] ;
wire \myreg.Reg[2][28] ;
wire \myreg.Reg[2][29] ;
wire \myreg.Reg[2][2] ;
wire \myreg.Reg[2][30] ;
wire \myreg.Reg[2][31] ;
wire \myreg.Reg[2][3] ;
wire \myreg.Reg[2][4] ;
wire \myreg.Reg[2][5] ;
wire \myreg.Reg[2][6] ;
wire \myreg.Reg[2][7] ;
wire \myreg.Reg[2][8] ;
wire \myreg.Reg[2][9] ;
wire \myreg.Reg[3][0] ;
wire \myreg.Reg[3][10] ;
wire \myreg.Reg[3][11] ;
wire \myreg.Reg[3][12] ;
wire \myreg.Reg[3][13] ;
wire \myreg.Reg[3][14] ;
wire \myreg.Reg[3][15] ;
wire \myreg.Reg[3][16] ;
wire \myreg.Reg[3][17] ;
wire \myreg.Reg[3][18] ;
wire \myreg.Reg[3][19] ;
wire \myreg.Reg[3][1] ;
wire \myreg.Reg[3][20] ;
wire \myreg.Reg[3][21] ;
wire \myreg.Reg[3][22] ;
wire \myreg.Reg[3][23] ;
wire \myreg.Reg[3][24] ;
wire \myreg.Reg[3][25] ;
wire \myreg.Reg[3][26] ;
wire \myreg.Reg[3][27] ;
wire \myreg.Reg[3][28] ;
wire \myreg.Reg[3][29] ;
wire \myreg.Reg[3][2] ;
wire \myreg.Reg[3][30] ;
wire \myreg.Reg[3][31] ;
wire \myreg.Reg[3][3] ;
wire \myreg.Reg[3][4] ;
wire \myreg.Reg[3][5] ;
wire \myreg.Reg[3][6] ;
wire \myreg.Reg[3][7] ;
wire \myreg.Reg[3][8] ;
wire \myreg.Reg[3][9] ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_10_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_11_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_12_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_13_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_14_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_15_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_16_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_17_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_18_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_19_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_1_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_20_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_21_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_22_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_23_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_24_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_25_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_26_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_27_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_28_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_29_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_2_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_30_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_31_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_3_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_4_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_5_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_6_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_7_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_8_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_9_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_D ;
wire \myreg.Reg[4][0] ;
wire \myreg.Reg[4][10] ;
wire \myreg.Reg[4][11] ;
wire \myreg.Reg[4][12] ;
wire \myreg.Reg[4][13] ;
wire \myreg.Reg[4][14] ;
wire \myreg.Reg[4][15] ;
wire \myreg.Reg[4][16] ;
wire \myreg.Reg[4][17] ;
wire \myreg.Reg[4][18] ;
wire \myreg.Reg[4][19] ;
wire \myreg.Reg[4][1] ;
wire \myreg.Reg[4][20] ;
wire \myreg.Reg[4][21] ;
wire \myreg.Reg[4][22] ;
wire \myreg.Reg[4][23] ;
wire \myreg.Reg[4][24] ;
wire \myreg.Reg[4][25] ;
wire \myreg.Reg[4][26] ;
wire \myreg.Reg[4][27] ;
wire \myreg.Reg[4][28] ;
wire \myreg.Reg[4][29] ;
wire \myreg.Reg[4][2] ;
wire \myreg.Reg[4][30] ;
wire \myreg.Reg[4][31] ;
wire \myreg.Reg[4][3] ;
wire \myreg.Reg[4][4] ;
wire \myreg.Reg[4][5] ;
wire \myreg.Reg[4][6] ;
wire \myreg.Reg[4][7] ;
wire \myreg.Reg[4][8] ;
wire \myreg.Reg[4][9] ;
wire \myreg.Reg[5][0] ;
wire \myreg.Reg[5][10] ;
wire \myreg.Reg[5][11] ;
wire \myreg.Reg[5][12] ;
wire \myreg.Reg[5][13] ;
wire \myreg.Reg[5][14] ;
wire \myreg.Reg[5][15] ;
wire \myreg.Reg[5][16] ;
wire \myreg.Reg[5][17] ;
wire \myreg.Reg[5][18] ;
wire \myreg.Reg[5][19] ;
wire \myreg.Reg[5][1] ;
wire \myreg.Reg[5][20] ;
wire \myreg.Reg[5][21] ;
wire \myreg.Reg[5][22] ;
wire \myreg.Reg[5][23] ;
wire \myreg.Reg[5][24] ;
wire \myreg.Reg[5][25] ;
wire \myreg.Reg[5][26] ;
wire \myreg.Reg[5][27] ;
wire \myreg.Reg[5][28] ;
wire \myreg.Reg[5][29] ;
wire \myreg.Reg[5][2] ;
wire \myreg.Reg[5][30] ;
wire \myreg.Reg[5][31] ;
wire \myreg.Reg[5][3] ;
wire \myreg.Reg[5][4] ;
wire \myreg.Reg[5][5] ;
wire \myreg.Reg[5][6] ;
wire \myreg.Reg[5][7] ;
wire \myreg.Reg[5][8] ;
wire \myreg.Reg[5][9] ;
wire \myreg.Reg[6][0] ;
wire \myreg.Reg[6][10] ;
wire \myreg.Reg[6][11] ;
wire \myreg.Reg[6][12] ;
wire \myreg.Reg[6][13] ;
wire \myreg.Reg[6][14] ;
wire \myreg.Reg[6][15] ;
wire \myreg.Reg[6][16] ;
wire \myreg.Reg[6][17] ;
wire \myreg.Reg[6][18] ;
wire \myreg.Reg[6][19] ;
wire \myreg.Reg[6][1] ;
wire \myreg.Reg[6][20] ;
wire \myreg.Reg[6][21] ;
wire \myreg.Reg[6][22] ;
wire \myreg.Reg[6][23] ;
wire \myreg.Reg[6][24] ;
wire \myreg.Reg[6][25] ;
wire \myreg.Reg[6][26] ;
wire \myreg.Reg[6][27] ;
wire \myreg.Reg[6][28] ;
wire \myreg.Reg[6][29] ;
wire \myreg.Reg[6][2] ;
wire \myreg.Reg[6][30] ;
wire \myreg.Reg[6][31] ;
wire \myreg.Reg[6][3] ;
wire \myreg.Reg[6][4] ;
wire \myreg.Reg[6][5] ;
wire \myreg.Reg[6][6] ;
wire \myreg.Reg[6][7] ;
wire \myreg.Reg[6][8] ;
wire \myreg.Reg[6][9] ;
wire \myreg.Reg[7][0] ;
wire \myreg.Reg[7][10] ;
wire \myreg.Reg[7][11] ;
wire \myreg.Reg[7][12] ;
wire \myreg.Reg[7][13] ;
wire \myreg.Reg[7][14] ;
wire \myreg.Reg[7][15] ;
wire \myreg.Reg[7][16] ;
wire \myreg.Reg[7][17] ;
wire \myreg.Reg[7][18] ;
wire \myreg.Reg[7][19] ;
wire \myreg.Reg[7][1] ;
wire \myreg.Reg[7][20] ;
wire \myreg.Reg[7][21] ;
wire \myreg.Reg[7][22] ;
wire \myreg.Reg[7][23] ;
wire \myreg.Reg[7][24] ;
wire \myreg.Reg[7][25] ;
wire \myreg.Reg[7][26] ;
wire \myreg.Reg[7][27] ;
wire \myreg.Reg[7][28] ;
wire \myreg.Reg[7][29] ;
wire \myreg.Reg[7][2] ;
wire \myreg.Reg[7][30] ;
wire \myreg.Reg[7][31] ;
wire \myreg.Reg[7][3] ;
wire \myreg.Reg[7][4] ;
wire \myreg.Reg[7][5] ;
wire \myreg.Reg[7][6] ;
wire \myreg.Reg[7][7] ;
wire \myreg.Reg[7][8] ;
wire \myreg.Reg[7][9] ;
wire \myreg.Reg[8][0] ;
wire \myreg.Reg[8][10] ;
wire \myreg.Reg[8][11] ;
wire \myreg.Reg[8][12] ;
wire \myreg.Reg[8][13] ;
wire \myreg.Reg[8][14] ;
wire \myreg.Reg[8][15] ;
wire \myreg.Reg[8][16] ;
wire \myreg.Reg[8][17] ;
wire \myreg.Reg[8][18] ;
wire \myreg.Reg[8][19] ;
wire \myreg.Reg[8][1] ;
wire \myreg.Reg[8][20] ;
wire \myreg.Reg[8][21] ;
wire \myreg.Reg[8][22] ;
wire \myreg.Reg[8][23] ;
wire \myreg.Reg[8][24] ;
wire \myreg.Reg[8][25] ;
wire \myreg.Reg[8][26] ;
wire \myreg.Reg[8][27] ;
wire \myreg.Reg[8][28] ;
wire \myreg.Reg[8][29] ;
wire \myreg.Reg[8][2] ;
wire \myreg.Reg[8][30] ;
wire \myreg.Reg[8][31] ;
wire \myreg.Reg[8][3] ;
wire \myreg.Reg[8][4] ;
wire \myreg.Reg[8][5] ;
wire \myreg.Reg[8][6] ;
wire \myreg.Reg[8][7] ;
wire \myreg.Reg[8][8] ;
wire \myreg.Reg[8][9] ;
wire \myreg.Reg[9][0] ;
wire \myreg.Reg[9][10] ;
wire \myreg.Reg[9][11] ;
wire \myreg.Reg[9][12] ;
wire \myreg.Reg[9][13] ;
wire \myreg.Reg[9][14] ;
wire \myreg.Reg[9][15] ;
wire \myreg.Reg[9][16] ;
wire \myreg.Reg[9][17] ;
wire \myreg.Reg[9][18] ;
wire \myreg.Reg[9][19] ;
wire \myreg.Reg[9][1] ;
wire \myreg.Reg[9][20] ;
wire \myreg.Reg[9][21] ;
wire \myreg.Reg[9][22] ;
wire \myreg.Reg[9][23] ;
wire \myreg.Reg[9][24] ;
wire \myreg.Reg[9][25] ;
wire \myreg.Reg[9][26] ;
wire \myreg.Reg[9][27] ;
wire \myreg.Reg[9][28] ;
wire \myreg.Reg[9][29] ;
wire \myreg.Reg[9][2] ;
wire \myreg.Reg[9][30] ;
wire \myreg.Reg[9][31] ;
wire \myreg.Reg[9][3] ;
wire \myreg.Reg[9][4] ;
wire \myreg.Reg[9][5] ;
wire \myreg.Reg[9][6] ;
wire \myreg.Reg[9][7] ;
wire \myreg.Reg[9][8] ;
wire \myreg.Reg[9][9] ;
wire \mysc.state_$_DFF_P__Q_1_D ;
wire \mysc.state_$_DFF_P__Q_2_D ;
wire \mysc.state_$_DFF_P__Q_D ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire fanout_net_41 ;
wire fanout_net_42 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [4:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [3:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] mepc ;
wire [31:0] mtvec ;
wire [63:0] \myclint.mtime ;
wire [0:0] \myclint.mtime_$_SDFF_PP0__Q_63_D ;
wire [31:0] \myec.mepc_tmp ;
wire [1:0] \myec.state ;
wire [31:0] \myexu.pc_jump ;
wire [3:0] \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [3:0] \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [2:0] \myidu.state ;
wire [31:0] \myifu.data_in ;
wire [3:0] \myifu.myicache.valid ;
wire [1:0] \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y ;
wire [2:0] \myifu.state ;
wire [2:0] \myifu.tmp_offset ;
wire [31:0] \mylsu.araddr_tmp ;
wire [31:0] \mylsu.awaddr_tmp ;
wire [4:0] \mylsu.state ;
wire [2:0] \mylsu.typ_tmp ;
wire [2:0] \myminixbar.state ;
wire [2:0] \mysc.state ;

assign \io_master_awid [1] = \io_master_awid [0] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [0] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awid [0] ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [0] = \io_master_arburst [0] ;
assign \io_master_arlen [1] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;

AND3_X4 _09013_ ( .A1(\myclint.mtime [2] ), .A2(\myclint.mtime [0] ), .A3(\myclint.mtime [1] ), .ZN(_01499_ ) );
AND3_X4 _09014_ ( .A1(_01499_ ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [3] ), .ZN(_01500_ ) );
AND3_X4 _09015_ ( .A1(_01500_ ), .A2(\myclint.mtime [6] ), .A3(\myclint.mtime [5] ), .ZN(_01501_ ) );
AND2_X2 _09016_ ( .A1(_01501_ ), .A2(\myclint.mtime [7] ), .ZN(_01502_ ) );
AND4_X1 _09017_ ( .A1(\myclint.mtime [14] ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .A4(\myclint.mtime [15] ), .ZN(_01503_ ) );
AND2_X1 _09018_ ( .A1(\myclint.mtime [8] ), .A2(\myclint.mtime [9] ), .ZN(_01504_ ) );
AND4_X1 _09019_ ( .A1(\myclint.mtime [10] ), .A2(_01503_ ), .A3(\myclint.mtime [11] ), .A4(_01504_ ), .ZN(_01505_ ) );
NAND2_X1 _09020_ ( .A1(_01502_ ), .A2(_01505_ ), .ZN(_01506_ ) );
AND2_X1 _09021_ ( .A1(\myclint.mtime [16] ), .A2(\myclint.mtime [17] ), .ZN(_01507_ ) );
AND3_X1 _09022_ ( .A1(_01507_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [19] ), .ZN(_01508_ ) );
AND4_X1 _09023_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_01509_ ) );
AND2_X1 _09024_ ( .A1(_01508_ ), .A2(_01509_ ), .ZN(_01510_ ) );
AND2_X1 _09025_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [31] ), .ZN(_01511_ ) );
AND2_X1 _09026_ ( .A1(\myclint.mtime [28] ), .A2(\myclint.mtime [29] ), .ZN(_01512_ ) );
AND2_X1 _09027_ ( .A1(\myclint.mtime [26] ), .A2(\myclint.mtime [27] ), .ZN(_01513_ ) );
AND3_X1 _09028_ ( .A1(_01513_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [25] ), .ZN(_01514_ ) );
NAND4_X1 _09029_ ( .A1(_01510_ ), .A2(_01511_ ), .A3(_01512_ ), .A4(_01514_ ), .ZN(_01515_ ) );
NOR2_X1 _09030_ ( .A1(_01506_ ), .A2(_01515_ ), .ZN(_01516_ ) );
AND2_X1 _09031_ ( .A1(\myclint.mtime [33] ), .A2(\myclint.mtime [32] ), .ZN(_01517_ ) );
AND3_X1 _09032_ ( .A1(_01517_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01518_ ) );
AND2_X1 _09033_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [39] ), .ZN(_01519_ ) );
AND2_X1 _09034_ ( .A1(\myclint.mtime [36] ), .A2(\myclint.mtime [37] ), .ZN(_01520_ ) );
AND3_X1 _09035_ ( .A1(_01518_ ), .A2(_01519_ ), .A3(_01520_ ), .ZN(_01521_ ) );
AND2_X1 _09036_ ( .A1(\myclint.mtime [44] ), .A2(\myclint.mtime [45] ), .ZN(_01522_ ) );
AND3_X1 _09037_ ( .A1(_01522_ ), .A2(\myclint.mtime [46] ), .A3(\myclint.mtime [47] ), .ZN(_01523_ ) );
AND2_X1 _09038_ ( .A1(\myclint.mtime [40] ), .A2(\myclint.mtime [41] ), .ZN(_01524_ ) );
AND3_X1 _09039_ ( .A1(_01524_ ), .A2(\myclint.mtime [42] ), .A3(\myclint.mtime [43] ), .ZN(_01525_ ) );
AND3_X1 _09040_ ( .A1(_01521_ ), .A2(_01523_ ), .A3(_01525_ ), .ZN(_01526_ ) );
AND2_X1 _09041_ ( .A1(_01516_ ), .A2(_01526_ ), .ZN(_01527_ ) );
AND2_X1 _09042_ ( .A1(\myclint.mtime [54] ), .A2(\myclint.mtime [55] ), .ZN(_01528_ ) );
AND2_X1 _09043_ ( .A1(\myclint.mtime [52] ), .A2(\myclint.mtime [53] ), .ZN(_01529_ ) );
AND2_X1 _09044_ ( .A1(\myclint.mtime [50] ), .A2(\myclint.mtime [51] ), .ZN(_01530_ ) );
AND2_X1 _09045_ ( .A1(\myclint.mtime [48] ), .A2(\myclint.mtime [49] ), .ZN(_01531_ ) );
AND4_X1 _09046_ ( .A1(_01528_ ), .A2(_01529_ ), .A3(_01530_ ), .A4(_01531_ ), .ZN(_01532_ ) );
AND2_X1 _09047_ ( .A1(_01527_ ), .A2(_01532_ ), .ZN(_01533_ ) );
AND4_X1 _09048_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .A4(\myclint.mtime [59] ), .ZN(_01534_ ) );
AND2_X1 _09049_ ( .A1(_01533_ ), .A2(_01534_ ), .ZN(_01535_ ) );
AND3_X1 _09050_ ( .A1(_01535_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01536_ ) );
INV_X1 _09051_ ( .A(_01536_ ), .ZN(_01537_ ) );
OR3_X1 _09052_ ( .A1(_01537_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [63] ), .ZN(_01538_ ) );
OAI21_X1 _09053_ ( .A(\myclint.mtime [63] ), .B1(_01537_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01539_ ) );
AOI21_X1 _09054_ ( .A(fanout_net_1 ), .B1(_01538_ ), .B2(_01539_ ), .ZN(_00000_ ) );
XNOR2_X1 _09055_ ( .A(_01536_ ), .B(\myclint.mtime [62] ), .ZN(_01540_ ) );
NOR2_X1 _09056_ ( .A1(_01540_ ), .A2(fanout_net_1 ), .ZN(_00001_ ) );
AND2_X1 _09057_ ( .A1(_01530_ ), .A2(_01531_ ), .ZN(_01541_ ) );
AND2_X1 _09058_ ( .A1(_01527_ ), .A2(_01541_ ), .ZN(_01542_ ) );
INV_X1 _09059_ ( .A(_01542_ ), .ZN(_01543_ ) );
OR3_X1 _09060_ ( .A1(_01543_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [53] ), .ZN(_01544_ ) );
OAI21_X1 _09061_ ( .A(\myclint.mtime [53] ), .B1(_01543_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01545_ ) );
AOI21_X1 _09062_ ( .A(fanout_net_1 ), .B1(_01544_ ), .B2(_01545_ ), .ZN(_00002_ ) );
XNOR2_X1 _09063_ ( .A(_01542_ ), .B(\myclint.mtime [52] ), .ZN(_01546_ ) );
NOR2_X1 _09064_ ( .A1(_01546_ ), .A2(fanout_net_1 ), .ZN(_00003_ ) );
INV_X1 _09065_ ( .A(fanout_net_1 ), .ZN(_01547_ ) );
BUF_X4 _09066_ ( .A(_01547_ ), .Z(_01548_ ) );
AND3_X4 _09067_ ( .A1(_01501_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [7] ), .ZN(_01549_ ) );
AND3_X4 _09068_ ( .A1(_01549_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [9] ), .ZN(_01550_ ) );
AND3_X4 _09069_ ( .A1(_01550_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [11] ), .ZN(_01551_ ) );
AND3_X4 _09070_ ( .A1(_01551_ ), .A2(\myclint.mtime [14] ), .A3(\myclint.mtime [13] ), .ZN(_01552_ ) );
AND3_X4 _09071_ ( .A1(_01552_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [15] ), .ZN(_01553_ ) );
AND3_X4 _09072_ ( .A1(_01553_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [17] ), .ZN(_01554_ ) );
AND3_X4 _09073_ ( .A1(_01554_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [19] ), .ZN(_01555_ ) );
AND3_X4 _09074_ ( .A1(_01555_ ), .A2(\myclint.mtime [22] ), .A3(\myclint.mtime [21] ), .ZN(_01556_ ) );
AND3_X4 _09075_ ( .A1(_01556_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [23] ), .ZN(_01557_ ) );
AND3_X2 _09076_ ( .A1(_01557_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [25] ), .ZN(_01558_ ) );
AND2_X4 _09077_ ( .A1(_01558_ ), .A2(\myclint.mtime [27] ), .ZN(_01559_ ) );
AND4_X1 _09078_ ( .A1(\myclint.mtime [33] ), .A2(_01559_ ), .A3(_01511_ ), .A4(_01512_ ), .ZN(_01560_ ) );
AND3_X2 _09079_ ( .A1(_01560_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01561_ ) );
AND2_X1 _09080_ ( .A1(_01561_ ), .A2(\myclint.mtime [35] ), .ZN(_01562_ ) );
AND3_X1 _09081_ ( .A1(_01562_ ), .A2(_01519_ ), .A3(_01520_ ), .ZN(_01563_ ) );
NAND2_X2 _09082_ ( .A1(_01563_ ), .A2(\myclint.mtime [40] ), .ZN(_01564_ ) );
INV_X1 _09083_ ( .A(\myclint.mtime [42] ), .ZN(_01565_ ) );
INV_X1 _09084_ ( .A(\myclint.mtime [41] ), .ZN(_01566_ ) );
NOR3_X4 _09085_ ( .A1(_01564_ ), .A2(_01565_ ), .A3(_01566_ ), .ZN(_01567_ ) );
AND2_X4 _09086_ ( .A1(_01567_ ), .A2(\myclint.mtime [43] ), .ZN(_01568_ ) );
NAND2_X1 _09087_ ( .A1(_01568_ ), .A2(_01523_ ), .ZN(_01569_ ) );
INV_X1 _09088_ ( .A(_01531_ ), .ZN(_01570_ ) );
NOR3_X1 _09089_ ( .A1(_01569_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01570_ ), .ZN(_01571_ ) );
OAI21_X1 _09090_ ( .A(_01548_ ), .B1(_01571_ ), .B2(\myclint.mtime [51] ), .ZN(_01572_ ) );
AND2_X1 _09091_ ( .A1(_01559_ ), .A2(_01512_ ), .ZN(_01573_ ) );
AND3_X1 _09092_ ( .A1(_01573_ ), .A2(_01517_ ), .A3(_01511_ ), .ZN(_01574_ ) );
AND2_X1 _09093_ ( .A1(_01574_ ), .A2(\myclint.mtime [34] ), .ZN(_01575_ ) );
AND2_X1 _09094_ ( .A1(_01575_ ), .A2(\myclint.mtime [35] ), .ZN(_01576_ ) );
AND3_X1 _09095_ ( .A1(_01576_ ), .A2(_01519_ ), .A3(_01520_ ), .ZN(_01577_ ) );
NAND2_X1 _09096_ ( .A1(_01577_ ), .A2(\myclint.mtime [40] ), .ZN(_01578_ ) );
NOR3_X1 _09097_ ( .A1(_01578_ ), .A2(_01565_ ), .A3(_01566_ ), .ZN(_01579_ ) );
AND2_X1 _09098_ ( .A1(_01579_ ), .A2(\myclint.mtime [43] ), .ZN(_01580_ ) );
AND2_X1 _09099_ ( .A1(_01580_ ), .A2(_01523_ ), .ZN(_01581_ ) );
INV_X1 _09100_ ( .A(_01581_ ), .ZN(_01582_ ) );
NOR3_X1 _09101_ ( .A1(_01582_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01570_ ), .ZN(_01583_ ) );
AOI21_X1 _09102_ ( .A(_01572_ ), .B1(_01583_ ), .B2(\myclint.mtime [51] ), .ZN(_00004_ ) );
INV_X1 _09103_ ( .A(_01516_ ), .ZN(_01584_ ) );
INV_X1 _09104_ ( .A(_01526_ ), .ZN(_01585_ ) );
OR4_X1 _09105_ ( .A1(\myclint.mtime [50] ), .A2(_01584_ ), .A3(_01570_ ), .A4(_01585_ ), .ZN(_01586_ ) );
AND3_X1 _09106_ ( .A1(_01516_ ), .A2(_01531_ ), .A3(_01526_ ), .ZN(_01587_ ) );
INV_X1 _09107_ ( .A(_01587_ ), .ZN(_01588_ ) );
NAND2_X1 _09108_ ( .A1(_01588_ ), .A2(\myclint.mtime [50] ), .ZN(_01589_ ) );
AOI21_X1 _09109_ ( .A(fanout_net_1 ), .B1(_01586_ ), .B2(_01589_ ), .ZN(_00005_ ) );
INV_X1 _09110_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01590_ ) );
AND4_X1 _09111_ ( .A1(\myclint.mtime [49] ), .A2(_01580_ ), .A3(_01590_ ), .A4(_01523_ ), .ZN(_01591_ ) );
BUF_X2 _09112_ ( .A(_01547_ ), .Z(_01592_ ) );
AND3_X1 _09113_ ( .A1(_01568_ ), .A2(_01590_ ), .A3(_01523_ ), .ZN(_01593_ ) );
OAI21_X1 _09114_ ( .A(_01592_ ), .B1(_01593_ ), .B2(\myclint.mtime [49] ), .ZN(_01594_ ) );
NOR2_X1 _09115_ ( .A1(_01591_ ), .A2(_01594_ ), .ZN(_00006_ ) );
OAI21_X1 _09116_ ( .A(\myclint.mtime [48] ), .B1(_01584_ ), .B2(_01585_ ), .ZN(_01595_ ) );
OR4_X1 _09117_ ( .A1(\myclint.mtime [48] ), .A2(_01506_ ), .A3(_01585_ ), .A4(_01515_ ), .ZN(_01596_ ) );
AOI21_X1 _09118_ ( .A(fanout_net_1 ), .B1(_01595_ ), .B2(_01596_ ), .ZN(_00007_ ) );
NAND3_X1 _09119_ ( .A1(_01567_ ), .A2(\myclint.mtime [43] ), .A3(_01522_ ), .ZN(_01597_ ) );
NOR2_X1 _09120_ ( .A1(_01597_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01598_ ) );
OAI21_X1 _09121_ ( .A(_01548_ ), .B1(_01598_ ), .B2(\myclint.mtime [47] ), .ZN(_01599_ ) );
NAND3_X1 _09122_ ( .A1(_01579_ ), .A2(\myclint.mtime [44] ), .A3(\myclint.mtime [43] ), .ZN(_01600_ ) );
INV_X1 _09123_ ( .A(\myclint.mtime [45] ), .ZN(_01601_ ) );
NOR3_X1 _09124_ ( .A1(_01600_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01601_ ), .ZN(_01602_ ) );
AOI21_X1 _09125_ ( .A(_01599_ ), .B1(_01602_ ), .B2(\myclint.mtime [47] ), .ZN(_00008_ ) );
AND2_X1 _09126_ ( .A1(_01516_ ), .A2(_01521_ ), .ZN(_01603_ ) );
AND3_X1 _09127_ ( .A1(_01603_ ), .A2(_01522_ ), .A3(_01525_ ), .ZN(_01604_ ) );
XNOR2_X1 _09128_ ( .A(_01604_ ), .B(\myclint.mtime [46] ), .ZN(_01605_ ) );
NOR2_X1 _09129_ ( .A1(_01605_ ), .A2(fanout_net_1 ), .ZN(_00009_ ) );
INV_X1 _09130_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01606_ ) );
NAND3_X1 _09131_ ( .A1(_01567_ ), .A2(_01606_ ), .A3(\myclint.mtime [43] ), .ZN(_01607_ ) );
AOI21_X1 _09132_ ( .A(fanout_net_1 ), .B1(_01607_ ), .B2(_01601_ ), .ZN(_01608_ ) );
NAND4_X1 _09133_ ( .A1(_01579_ ), .A2(\myclint.mtime [45] ), .A3(_01606_ ), .A4(\myclint.mtime [43] ), .ZN(_01609_ ) );
AND2_X1 _09134_ ( .A1(_01608_ ), .A2(_01609_ ), .ZN(_00010_ ) );
AND2_X1 _09135_ ( .A1(_01603_ ), .A2(_01525_ ), .ZN(_01610_ ) );
XNOR2_X1 _09136_ ( .A(_01610_ ), .B(\myclint.mtime [44] ), .ZN(_01611_ ) );
NOR2_X1 _09137_ ( .A1(_01611_ ), .A2(fanout_net_1 ), .ZN(_00011_ ) );
INV_X1 _09138_ ( .A(_01535_ ), .ZN(_01612_ ) );
OR3_X1 _09139_ ( .A1(_01612_ ), .A2(\myclint.mtime [61] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01613_ ) );
OAI21_X1 _09140_ ( .A(\myclint.mtime [61] ), .B1(_01612_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01614_ ) );
AOI21_X1 _09141_ ( .A(fanout_net_1 ), .B1(_01613_ ), .B2(_01614_ ), .ZN(_00012_ ) );
NOR3_X1 _09142_ ( .A1(_01564_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01566_ ), .ZN(_01615_ ) );
OAI21_X1 _09143_ ( .A(_01548_ ), .B1(_01615_ ), .B2(\myclint.mtime [43] ), .ZN(_01616_ ) );
NOR3_X1 _09144_ ( .A1(_01578_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01566_ ), .ZN(_01617_ ) );
AOI21_X1 _09145_ ( .A(_01616_ ), .B1(_01617_ ), .B2(\myclint.mtime [43] ), .ZN(_00013_ ) );
BUF_X2 _09146_ ( .A(_01548_ ), .Z(_01618_ ) );
AND3_X1 _09147_ ( .A1(_01563_ ), .A2(\myclint.mtime [40] ), .A3(\myclint.mtime [41] ), .ZN(_01619_ ) );
OAI21_X1 _09148_ ( .A(_01618_ ), .B1(_01619_ ), .B2(\myclint.mtime [42] ), .ZN(_01620_ ) );
NOR2_X1 _09149_ ( .A1(_01620_ ), .A2(_01567_ ), .ZN(_00014_ ) );
INV_X1 _09150_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01621_ ) );
NAND2_X1 _09151_ ( .A1(_01563_ ), .A2(_01621_ ), .ZN(_01622_ ) );
AOI21_X1 _09152_ ( .A(fanout_net_1 ), .B1(_01622_ ), .B2(_01566_ ), .ZN(_01623_ ) );
AND2_X1 _09153_ ( .A1(_01576_ ), .A2(_01520_ ), .ZN(_01624_ ) );
NAND4_X1 _09154_ ( .A1(_01624_ ), .A2(\myclint.mtime [41] ), .A3(_01621_ ), .A4(_01519_ ), .ZN(_01625_ ) );
AND2_X1 _09155_ ( .A1(_01623_ ), .A2(_01625_ ), .ZN(_00015_ ) );
XNOR2_X1 _09156_ ( .A(_01603_ ), .B(\myclint.mtime [40] ), .ZN(_01626_ ) );
NOR2_X1 _09157_ ( .A1(_01626_ ), .A2(fanout_net_1 ), .ZN(_00016_ ) );
NAND3_X1 _09158_ ( .A1(_01516_ ), .A2(_01520_ ), .A3(_01518_ ), .ZN(_01627_ ) );
OR3_X1 _09159_ ( .A1(_01627_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [39] ), .ZN(_01628_ ) );
OAI21_X1 _09160_ ( .A(\myclint.mtime [39] ), .B1(_01627_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01629_ ) );
AOI21_X1 _09161_ ( .A(fanout_net_1 ), .B1(_01628_ ), .B2(_01629_ ), .ZN(_00017_ ) );
OR2_X1 _09162_ ( .A1(_01627_ ), .A2(\myclint.mtime [38] ), .ZN(_01630_ ) );
NAND2_X1 _09163_ ( .A1(_01627_ ), .A2(\myclint.mtime [38] ), .ZN(_01631_ ) );
AOI21_X1 _09164_ ( .A(fanout_net_1 ), .B1(_01630_ ), .B2(_01631_ ), .ZN(_00018_ ) );
INV_X1 _09165_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01632_ ) );
AND4_X1 _09166_ ( .A1(\myclint.mtime [37] ), .A2(_01575_ ), .A3(_01632_ ), .A4(\myclint.mtime [35] ), .ZN(_01633_ ) );
AND3_X1 _09167_ ( .A1(_01561_ ), .A2(_01632_ ), .A3(\myclint.mtime [35] ), .ZN(_01634_ ) );
OAI21_X1 _09168_ ( .A(_01592_ ), .B1(_01634_ ), .B2(\myclint.mtime [37] ), .ZN(_01635_ ) );
NOR2_X1 _09169_ ( .A1(_01633_ ), .A2(_01635_ ), .ZN(_00019_ ) );
AND2_X1 _09170_ ( .A1(_01516_ ), .A2(_01518_ ), .ZN(_01636_ ) );
XNOR2_X1 _09171_ ( .A(_01636_ ), .B(\myclint.mtime [36] ), .ZN(_01637_ ) );
NOR2_X1 _09172_ ( .A1(_01637_ ), .A2(fanout_net_1 ), .ZN(_00020_ ) );
AND2_X1 _09173_ ( .A1(_01502_ ), .A2(_01505_ ), .ZN(_01638_ ) );
AND4_X1 _09174_ ( .A1(_01511_ ), .A2(_01510_ ), .A3(_01512_ ), .A4(_01514_ ), .ZN(_01639_ ) );
NAND3_X1 _09175_ ( .A1(_01638_ ), .A2(_01517_ ), .A3(_01639_ ), .ZN(_01640_ ) );
OR3_X1 _09176_ ( .A1(_01640_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [35] ), .ZN(_01641_ ) );
OAI21_X1 _09177_ ( .A(\myclint.mtime [35] ), .B1(_01640_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01642_ ) );
AOI21_X1 _09178_ ( .A(fanout_net_1 ), .B1(_01641_ ), .B2(_01642_ ), .ZN(_00021_ ) );
NAND4_X1 _09179_ ( .A1(_01559_ ), .A2(\myclint.mtime [33] ), .A3(_01511_ ), .A4(_01512_ ), .ZN(_01643_ ) );
INV_X1 _09180_ ( .A(\myclint.mtime [32] ), .ZN(_01644_ ) );
NOR2_X1 _09181_ ( .A1(_01643_ ), .A2(_01644_ ), .ZN(_01645_ ) );
OAI21_X1 _09182_ ( .A(_01618_ ), .B1(_01645_ ), .B2(\myclint.mtime [34] ), .ZN(_01646_ ) );
NOR2_X1 _09183_ ( .A1(_01646_ ), .A2(_01561_ ), .ZN(_00022_ ) );
XNOR2_X1 _09184_ ( .A(_01535_ ), .B(\myclint.mtime [60] ), .ZN(_01647_ ) );
NOR2_X1 _09185_ ( .A1(_01647_ ), .A2(fanout_net_1 ), .ZN(_00023_ ) );
OR3_X1 _09186_ ( .A1(_01506_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_01515_ ), .ZN(_01648_ ) );
NAND2_X1 _09187_ ( .A1(_01648_ ), .A2(\myclint.mtime [33] ), .ZN(_01649_ ) );
OR4_X1 _09188_ ( .A1(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A2(_01506_ ), .A3(\myclint.mtime [33] ), .A4(_01515_ ), .ZN(_01650_ ) );
AOI21_X1 _09189_ ( .A(fanout_net_1 ), .B1(_01649_ ), .B2(_01650_ ), .ZN(_00024_ ) );
OAI21_X1 _09190_ ( .A(\myclint.mtime [32] ), .B1(_01506_ ), .B2(_01515_ ), .ZN(_01651_ ) );
NAND4_X1 _09191_ ( .A1(_01639_ ), .A2(_01502_ ), .A3(_01644_ ), .A4(_01505_ ), .ZN(_01652_ ) );
AOI21_X1 _09192_ ( .A(fanout_net_1 ), .B1(_01651_ ), .B2(_01652_ ), .ZN(_00025_ ) );
AND2_X1 _09193_ ( .A1(_01638_ ), .A2(_01510_ ), .ZN(_01653_ ) );
NAND3_X1 _09194_ ( .A1(_01653_ ), .A2(_01512_ ), .A3(_01514_ ), .ZN(_01654_ ) );
OR3_X1 _09195_ ( .A1(_01654_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [31] ), .ZN(_01655_ ) );
OAI21_X1 _09196_ ( .A(\myclint.mtime [31] ), .B1(_01654_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01656_ ) );
AOI21_X1 _09197_ ( .A(fanout_net_1 ), .B1(_01655_ ), .B2(_01656_ ), .ZN(_00026_ ) );
OR2_X1 _09198_ ( .A1(_01654_ ), .A2(\myclint.mtime [30] ), .ZN(_01657_ ) );
NAND2_X1 _09199_ ( .A1(_01654_ ), .A2(\myclint.mtime [30] ), .ZN(_01658_ ) );
AOI21_X1 _09200_ ( .A(fanout_net_1 ), .B1(_01657_ ), .B2(_01658_ ), .ZN(_00027_ ) );
INV_X1 _09201_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01659_ ) );
AND3_X1 _09202_ ( .A1(_01558_ ), .A2(_01659_ ), .A3(\myclint.mtime [27] ), .ZN(_01660_ ) );
AND2_X1 _09203_ ( .A1(_01660_ ), .A2(\myclint.mtime [29] ), .ZN(_01661_ ) );
OAI21_X1 _09204_ ( .A(_01592_ ), .B1(_01660_ ), .B2(\myclint.mtime [29] ), .ZN(_01662_ ) );
NOR2_X1 _09205_ ( .A1(_01661_ ), .A2(_01662_ ), .ZN(_00028_ ) );
NAND2_X1 _09206_ ( .A1(_01653_ ), .A2(_01514_ ), .ZN(_01663_ ) );
OR2_X1 _09207_ ( .A1(_01663_ ), .A2(\myclint.mtime [28] ), .ZN(_01664_ ) );
NAND2_X1 _09208_ ( .A1(_01663_ ), .A2(\myclint.mtime [28] ), .ZN(_01665_ ) );
AOI21_X1 _09209_ ( .A(fanout_net_1 ), .B1(_01664_ ), .B2(_01665_ ), .ZN(_00029_ ) );
NAND3_X1 _09210_ ( .A1(_01653_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [25] ), .ZN(_01666_ ) );
OR3_X1 _09211_ ( .A1(_01666_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [27] ), .ZN(_01667_ ) );
OAI21_X1 _09212_ ( .A(\myclint.mtime [27] ), .B1(_01666_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01668_ ) );
AOI21_X1 _09213_ ( .A(fanout_net_1 ), .B1(_01667_ ), .B2(_01668_ ), .ZN(_00030_ ) );
BUF_X4 _09214_ ( .A(_01548_ ), .Z(_01669_ ) );
AND2_X1 _09215_ ( .A1(_01557_ ), .A2(\myclint.mtime [25] ), .ZN(_01670_ ) );
OAI21_X1 _09216_ ( .A(_01669_ ), .B1(_01670_ ), .B2(\myclint.mtime [26] ), .ZN(_01671_ ) );
NOR2_X1 _09217_ ( .A1(_01671_ ), .A2(_01558_ ), .ZN(_00031_ ) );
INV_X1 _09218_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01672_ ) );
AND3_X1 _09219_ ( .A1(_01556_ ), .A2(_01672_ ), .A3(\myclint.mtime [23] ), .ZN(_01673_ ) );
AND2_X1 _09220_ ( .A1(_01673_ ), .A2(\myclint.mtime [25] ), .ZN(_01674_ ) );
OAI21_X1 _09221_ ( .A(_01592_ ), .B1(_01673_ ), .B2(\myclint.mtime [25] ), .ZN(_01675_ ) );
NOR2_X1 _09222_ ( .A1(_01674_ ), .A2(_01675_ ), .ZN(_00032_ ) );
AND2_X1 _09223_ ( .A1(_01556_ ), .A2(\myclint.mtime [23] ), .ZN(_01676_ ) );
OAI21_X1 _09224_ ( .A(_01669_ ), .B1(_01676_ ), .B2(\myclint.mtime [24] ), .ZN(_01677_ ) );
NOR2_X1 _09225_ ( .A1(_01677_ ), .A2(_01557_ ), .ZN(_00033_ ) );
AND2_X1 _09226_ ( .A1(\myclint.mtime [56] ), .A2(\myclint.mtime [57] ), .ZN(_01678_ ) );
NAND3_X1 _09227_ ( .A1(_01527_ ), .A2(_01678_ ), .A3(_01532_ ), .ZN(_01679_ ) );
OR3_X1 _09228_ ( .A1(_01679_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [59] ), .ZN(_01680_ ) );
OAI21_X1 _09229_ ( .A(\myclint.mtime [59] ), .B1(_01679_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01681_ ) );
AOI21_X1 _09230_ ( .A(fanout_net_1 ), .B1(_01680_ ), .B2(_01681_ ), .ZN(_00034_ ) );
AND2_X1 _09231_ ( .A1(_01638_ ), .A2(_01508_ ), .ZN(_01682_ ) );
NAND3_X1 _09232_ ( .A1(_01682_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .ZN(_01683_ ) );
OR3_X1 _09233_ ( .A1(_01683_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [23] ), .ZN(_01684_ ) );
OAI21_X1 _09234_ ( .A(\myclint.mtime [23] ), .B1(_01683_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01685_ ) );
AOI21_X1 _09235_ ( .A(fanout_net_1 ), .B1(_01684_ ), .B2(_01685_ ), .ZN(_00035_ ) );
AND2_X1 _09236_ ( .A1(_01555_ ), .A2(\myclint.mtime [21] ), .ZN(_01686_ ) );
OAI21_X1 _09237_ ( .A(_01669_ ), .B1(_01686_ ), .B2(\myclint.mtime [22] ), .ZN(_01687_ ) );
NOR2_X1 _09238_ ( .A1(_01687_ ), .A2(_01556_ ), .ZN(_00036_ ) );
INV_X1 _09239_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01688_ ) );
AND3_X1 _09240_ ( .A1(_01554_ ), .A2(_01688_ ), .A3(\myclint.mtime [19] ), .ZN(_01689_ ) );
AND2_X1 _09241_ ( .A1(_01689_ ), .A2(\myclint.mtime [21] ), .ZN(_01690_ ) );
OAI21_X1 _09242_ ( .A(_01592_ ), .B1(_01689_ ), .B2(\myclint.mtime [21] ), .ZN(_01691_ ) );
NOR2_X1 _09243_ ( .A1(_01690_ ), .A2(_01691_ ), .ZN(_00037_ ) );
AND2_X1 _09244_ ( .A1(_01554_ ), .A2(\myclint.mtime [19] ), .ZN(_01692_ ) );
OAI21_X1 _09245_ ( .A(_01669_ ), .B1(_01692_ ), .B2(\myclint.mtime [20] ), .ZN(_01693_ ) );
NOR2_X1 _09246_ ( .A1(_01693_ ), .A2(_01555_ ), .ZN(_00038_ ) );
NAND3_X1 _09247_ ( .A1(_01502_ ), .A2(_01505_ ), .A3(_01507_ ), .ZN(_01694_ ) );
OR3_X1 _09248_ ( .A1(_01694_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [19] ), .ZN(_01695_ ) );
OAI21_X1 _09249_ ( .A(\myclint.mtime [19] ), .B1(_01694_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01696_ ) );
AOI21_X1 _09250_ ( .A(fanout_net_1 ), .B1(_01695_ ), .B2(_01696_ ), .ZN(_00039_ ) );
AND2_X1 _09251_ ( .A1(_01553_ ), .A2(\myclint.mtime [17] ), .ZN(_01697_ ) );
OAI21_X1 _09252_ ( .A(_01669_ ), .B1(_01697_ ), .B2(\myclint.mtime [18] ), .ZN(_01698_ ) );
NOR2_X1 _09253_ ( .A1(_01698_ ), .A2(_01554_ ), .ZN(_00040_ ) );
INV_X1 _09254_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01699_ ) );
AND3_X1 _09255_ ( .A1(_01552_ ), .A2(_01699_ ), .A3(\myclint.mtime [15] ), .ZN(_01700_ ) );
AND2_X1 _09256_ ( .A1(_01700_ ), .A2(\myclint.mtime [17] ), .ZN(_01701_ ) );
OAI21_X1 _09257_ ( .A(_01592_ ), .B1(_01700_ ), .B2(\myclint.mtime [17] ), .ZN(_01702_ ) );
NOR2_X1 _09258_ ( .A1(_01701_ ), .A2(_01702_ ), .ZN(_00041_ ) );
AND2_X1 _09259_ ( .A1(_01552_ ), .A2(\myclint.mtime [15] ), .ZN(_01703_ ) );
OAI21_X1 _09260_ ( .A(_01669_ ), .B1(_01703_ ), .B2(\myclint.mtime [16] ), .ZN(_01704_ ) );
NOR2_X1 _09261_ ( .A1(_01704_ ), .A2(_01553_ ), .ZN(_00042_ ) );
AND3_X1 _09262_ ( .A1(_01504_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [11] ), .ZN(_01705_ ) );
AND2_X1 _09263_ ( .A1(_01502_ ), .A2(_01705_ ), .ZN(_01706_ ) );
NAND3_X1 _09264_ ( .A1(_01706_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .ZN(_01707_ ) );
OR3_X1 _09265_ ( .A1(_01707_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [15] ), .ZN(_01708_ ) );
OAI21_X1 _09266_ ( .A(\myclint.mtime [15] ), .B1(_01707_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01709_ ) );
AOI21_X1 _09267_ ( .A(fanout_net_1 ), .B1(_01708_ ), .B2(_01709_ ), .ZN(_00043_ ) );
AND2_X1 _09268_ ( .A1(_01551_ ), .A2(\myclint.mtime [13] ), .ZN(_01710_ ) );
OAI21_X1 _09269_ ( .A(_01669_ ), .B1(_01710_ ), .B2(\myclint.mtime [14] ), .ZN(_01711_ ) );
NOR2_X1 _09270_ ( .A1(_01711_ ), .A2(_01552_ ), .ZN(_00044_ ) );
OR2_X1 _09271_ ( .A1(_01679_ ), .A2(\myclint.mtime [58] ), .ZN(_01712_ ) );
NAND2_X1 _09272_ ( .A1(_01679_ ), .A2(\myclint.mtime [58] ), .ZN(_01713_ ) );
AOI21_X1 _09273_ ( .A(fanout_net_1 ), .B1(_01712_ ), .B2(_01713_ ), .ZN(_00045_ ) );
INV_X1 _09274_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01714_ ) );
AND3_X1 _09275_ ( .A1(_01550_ ), .A2(_01714_ ), .A3(\myclint.mtime [11] ), .ZN(_01715_ ) );
AND2_X1 _09276_ ( .A1(_01715_ ), .A2(\myclint.mtime [13] ), .ZN(_01716_ ) );
OAI21_X1 _09277_ ( .A(_01548_ ), .B1(_01715_ ), .B2(\myclint.mtime [13] ), .ZN(_01717_ ) );
NOR2_X1 _09278_ ( .A1(_01716_ ), .A2(_01717_ ), .ZN(_00046_ ) );
AND2_X1 _09279_ ( .A1(_01550_ ), .A2(\myclint.mtime [11] ), .ZN(_01718_ ) );
OAI21_X1 _09280_ ( .A(_01669_ ), .B1(_01718_ ), .B2(\myclint.mtime [12] ), .ZN(_01719_ ) );
NOR2_X1 _09281_ ( .A1(_01719_ ), .A2(_01551_ ), .ZN(_00047_ ) );
INV_X1 _09282_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01720_ ) );
AND3_X1 _09283_ ( .A1(_01549_ ), .A2(_01720_ ), .A3(\myclint.mtime [9] ), .ZN(_01721_ ) );
AND2_X1 _09284_ ( .A1(_01721_ ), .A2(\myclint.mtime [11] ), .ZN(_01722_ ) );
OAI21_X1 _09285_ ( .A(_01548_ ), .B1(_01721_ ), .B2(\myclint.mtime [11] ), .ZN(_01723_ ) );
NOR2_X1 _09286_ ( .A1(_01722_ ), .A2(_01723_ ), .ZN(_00048_ ) );
AOI21_X1 _09287_ ( .A(\myclint.mtime [10] ), .B1(_01549_ ), .B2(\myclint.mtime [9] ), .ZN(_01724_ ) );
NOR3_X1 _09288_ ( .A1(_01550_ ), .A2(_01724_ ), .A3(fanout_net_1 ), .ZN(_00049_ ) );
INV_X1 _09289_ ( .A(_01502_ ), .ZN(_01725_ ) );
OR3_X1 _09290_ ( .A1(_01725_ ), .A2(\myclint.mtime [9] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01726_ ) );
OAI21_X1 _09291_ ( .A(\myclint.mtime [9] ), .B1(_01725_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01727_ ) );
AOI21_X1 _09292_ ( .A(fanout_net_2 ), .B1(_01726_ ), .B2(_01727_ ), .ZN(_00050_ ) );
OAI21_X1 _09293_ ( .A(_01669_ ), .B1(_01502_ ), .B2(\myclint.mtime [8] ), .ZN(_01728_ ) );
NOR2_X1 _09294_ ( .A1(_01728_ ), .A2(_01549_ ), .ZN(_00051_ ) );
AND2_X1 _09295_ ( .A1(_01500_ ), .A2(\myclint.mtime [5] ), .ZN(_01729_ ) );
INV_X1 _09296_ ( .A(_01729_ ), .ZN(_01730_ ) );
OR3_X1 _09297_ ( .A1(_01730_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [7] ), .ZN(_01731_ ) );
OAI21_X1 _09298_ ( .A(\myclint.mtime [7] ), .B1(_01730_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01732_ ) );
AOI21_X1 _09299_ ( .A(fanout_net_2 ), .B1(_01731_ ), .B2(_01732_ ), .ZN(_00052_ ) );
OAI21_X1 _09300_ ( .A(_01669_ ), .B1(_01729_ ), .B2(\myclint.mtime [6] ), .ZN(_01733_ ) );
NOR2_X1 _09301_ ( .A1(_01733_ ), .A2(_01501_ ), .ZN(_00053_ ) );
AND2_X1 _09302_ ( .A1(_01499_ ), .A2(\myclint.mtime [3] ), .ZN(_01734_ ) );
INV_X1 _09303_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01735_ ) );
AND3_X1 _09304_ ( .A1(_01734_ ), .A2(\myclint.mtime [5] ), .A3(_01735_ ), .ZN(_01736_ ) );
AOI21_X1 _09305_ ( .A(\myclint.mtime [5] ), .B1(_01734_ ), .B2(_01735_ ), .ZN(_01737_ ) );
NOR3_X1 _09306_ ( .A1(_01736_ ), .A2(_01737_ ), .A3(fanout_net_2 ), .ZN(_00054_ ) );
OAI21_X1 _09307_ ( .A(_01592_ ), .B1(_01734_ ), .B2(\myclint.mtime [4] ), .ZN(_01738_ ) );
NOR2_X1 _09308_ ( .A1(_01738_ ), .A2(_01500_ ), .ZN(_00055_ ) );
NOR2_X1 _09309_ ( .A1(_01569_ ), .A2(_01570_ ), .ZN(_01739_ ) );
AND2_X1 _09310_ ( .A1(_01739_ ), .A2(_01530_ ), .ZN(_01740_ ) );
AND2_X1 _09311_ ( .A1(_01740_ ), .A2(_01529_ ), .ZN(_01741_ ) );
INV_X1 _09312_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01742_ ) );
AND3_X1 _09313_ ( .A1(_01741_ ), .A2(_01742_ ), .A3(_01528_ ), .ZN(_01743_ ) );
OAI21_X1 _09314_ ( .A(_01548_ ), .B1(_01743_ ), .B2(\myclint.mtime [57] ), .ZN(_01744_ ) );
AND2_X1 _09315_ ( .A1(_01581_ ), .A2(_01531_ ), .ZN(_01745_ ) );
AND2_X1 _09316_ ( .A1(_01745_ ), .A2(_01530_ ), .ZN(_01746_ ) );
AND2_X1 _09317_ ( .A1(_01746_ ), .A2(_01529_ ), .ZN(_01747_ ) );
AND3_X1 _09318_ ( .A1(_01747_ ), .A2(_01742_ ), .A3(_01528_ ), .ZN(_01748_ ) );
AOI21_X1 _09319_ ( .A(_01744_ ), .B1(_01748_ ), .B2(\myclint.mtime [57] ), .ZN(_00056_ ) );
AND2_X1 _09320_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01749_ ) );
INV_X1 _09321_ ( .A(_01749_ ), .ZN(_01750_ ) );
OR3_X1 _09322_ ( .A1(_01750_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [3] ), .ZN(_01751_ ) );
OAI21_X1 _09323_ ( .A(\myclint.mtime [3] ), .B1(_01750_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01752_ ) );
AOI21_X1 _09324_ ( .A(fanout_net_2 ), .B1(_01751_ ), .B2(_01752_ ), .ZN(_00057_ ) );
AOI21_X1 _09325_ ( .A(\myclint.mtime [2] ), .B1(\myclint.mtime [0] ), .B2(\myclint.mtime [1] ), .ZN(_01753_ ) );
NOR3_X1 _09326_ ( .A1(_01499_ ), .A2(_01753_ ), .A3(fanout_net_2 ), .ZN(_00058_ ) );
NOR2_X1 _09327_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01754_ ) );
NOR3_X1 _09328_ ( .A1(_01749_ ), .A2(_01754_ ), .A3(fanout_net_2 ), .ZN(_00059_ ) );
AND2_X1 _09329_ ( .A1(_01618_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_00060_ ) );
XNOR2_X1 _09330_ ( .A(_01533_ ), .B(\myclint.mtime [56] ), .ZN(_01755_ ) );
NOR2_X1 _09331_ ( .A1(_01755_ ), .A2(fanout_net_2 ), .ZN(_00061_ ) );
NAND3_X1 _09332_ ( .A1(_01527_ ), .A2(_01529_ ), .A3(_01541_ ), .ZN(_01756_ ) );
OR3_X1 _09333_ ( .A1(_01756_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [55] ), .ZN(_01757_ ) );
OAI21_X1 _09334_ ( .A(\myclint.mtime [55] ), .B1(_01756_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01758_ ) );
AOI21_X1 _09335_ ( .A(fanout_net_2 ), .B1(_01757_ ), .B2(_01758_ ), .ZN(_00062_ ) );
OR2_X1 _09336_ ( .A1(_01756_ ), .A2(\myclint.mtime [54] ), .ZN(_01759_ ) );
NAND2_X1 _09337_ ( .A1(_01756_ ), .A2(\myclint.mtime [54] ), .ZN(_01760_ ) );
AOI21_X1 _09338_ ( .A(fanout_net_2 ), .B1(_01759_ ), .B2(_01760_ ), .ZN(_00063_ ) );
INV_X32 _09339_ ( .A(fanout_net_40 ), .ZN(_01761_ ) );
BUF_X32 _09340_ ( .A(_01761_ ), .Z(_01762_ ) );
OR2_X1 _09341_ ( .A1(_01762_ ), .A2(\myifu.myicache.tag[1][25] ), .ZN(_01763_ ) );
INV_X32 _09342_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01764_ ) );
BUF_X32 _09343_ ( .A(_01764_ ), .Z(_01765_ ) );
OAI211_X1 _09344_ ( .A(_01763_ ), .B(_01765_ ), .C1(fanout_net_40 ), .C2(\myifu.myicache.tag[0][25] ), .ZN(_01766_ ) );
OR2_X1 _09345_ ( .A1(_01762_ ), .A2(\myifu.myicache.tag[3][25] ), .ZN(_01767_ ) );
OAI211_X1 _09346_ ( .A(_01767_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_40 ), .C2(\myifu.myicache.tag[2][25] ), .ZN(_01768_ ) );
NAND2_X1 _09347_ ( .A1(_01766_ ), .A2(_01768_ ), .ZN(_01769_ ) );
INV_X1 _09348_ ( .A(\IF_ID_pc [30] ), .ZN(_01770_ ) );
XNOR2_X1 _09349_ ( .A(_01769_ ), .B(_01770_ ), .ZN(_01771_ ) );
OR2_X4 _09350_ ( .A1(_01762_ ), .A2(\myifu.myicache.tag[1][23] ), .ZN(_01772_ ) );
OAI211_X2 _09351_ ( .A(_01772_ ), .B(_01765_ ), .C1(fanout_net_40 ), .C2(\myifu.myicache.tag[0][23] ), .ZN(_01773_ ) );
OR2_X1 _09352_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[2][23] ), .ZN(_01774_ ) );
BUF_X16 _09353_ ( .A(_01761_ ), .Z(_01775_ ) );
OAI211_X1 _09354_ ( .A(_01774_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01775_ ), .C2(\myifu.myicache.tag[3][23] ), .ZN(_01776_ ) );
INV_X1 _09355_ ( .A(\IF_ID_pc [28] ), .ZN(_01777_ ) );
AND3_X2 _09356_ ( .A1(_01773_ ), .A2(_01776_ ), .A3(_01777_ ), .ZN(_01778_ ) );
AOI21_X1 _09357_ ( .A(_01777_ ), .B1(_01773_ ), .B2(_01776_ ), .ZN(_01779_ ) );
OR2_X4 _09358_ ( .A1(_01761_ ), .A2(\myifu.myicache.tag[1][6] ), .ZN(_01780_ ) );
OAI211_X1 _09359_ ( .A(_01780_ ), .B(_01765_ ), .C1(fanout_net_40 ), .C2(\myifu.myicache.tag[0][6] ), .ZN(_01781_ ) );
OR2_X4 _09360_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[2][6] ), .ZN(_01782_ ) );
OAI211_X1 _09361_ ( .A(_01782_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01762_ ), .C2(\myifu.myicache.tag[3][6] ), .ZN(_01783_ ) );
INV_X1 _09362_ ( .A(\IF_ID_pc [11] ), .ZN(_01784_ ) );
AND3_X1 _09363_ ( .A1(_01781_ ), .A2(_01783_ ), .A3(_01784_ ), .ZN(_01785_ ) );
AOI21_X1 _09364_ ( .A(_01784_ ), .B1(_01781_ ), .B2(_01783_ ), .ZN(_01786_ ) );
OAI22_X1 _09365_ ( .A1(_01778_ ), .A2(_01779_ ), .B1(_01785_ ), .B2(_01786_ ), .ZN(_01787_ ) );
OR2_X1 _09366_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[0][14] ), .ZN(_01788_ ) );
BUF_X4 _09367_ ( .A(_01762_ ), .Z(_01789_ ) );
OAI211_X1 _09368_ ( .A(_01788_ ), .B(_01765_ ), .C1(_01789_ ), .C2(\myifu.myicache.tag[1][14] ), .ZN(_01790_ ) );
OR2_X1 _09369_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[2][14] ), .ZN(_01791_ ) );
OAI211_X1 _09370_ ( .A(_01791_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01789_ ), .C2(\myifu.myicache.tag[3][14] ), .ZN(_01792_ ) );
AND3_X1 _09371_ ( .A1(_01790_ ), .A2(_01792_ ), .A3(\IF_ID_pc [19] ), .ZN(_01793_ ) );
AOI21_X1 _09372_ ( .A(\IF_ID_pc [19] ), .B1(_01790_ ), .B2(_01792_ ), .ZN(_01794_ ) );
OR4_X2 _09373_ ( .A1(_01771_ ), .A2(_01787_ ), .A3(_01793_ ), .A4(_01794_ ), .ZN(_01795_ ) );
MUX2_X1 _09374_ ( .A(\myifu.myicache.valid [2] ), .B(\myifu.myicache.valid [3] ), .S(fanout_net_40 ), .Z(_01796_ ) );
AND2_X1 _09375_ ( .A1(_01796_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01797_ ) );
BUF_X2 _09376_ ( .A(_01764_ ), .Z(_01798_ ) );
MUX2_X1 _09377_ ( .A(\myifu.myicache.valid [0] ), .B(\myifu.myicache.valid [1] ), .S(fanout_net_40 ), .Z(_01799_ ) );
AOI21_X1 _09378_ ( .A(_01797_ ), .B1(_01798_ ), .B2(_01799_ ), .ZN(_01800_ ) );
OR2_X4 _09379_ ( .A1(_01762_ ), .A2(\myifu.myicache.tag[3][17] ), .ZN(_01801_ ) );
OAI211_X4 _09380_ ( .A(_01801_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_40 ), .C2(\myifu.myicache.tag[2][17] ), .ZN(_01802_ ) );
OR2_X1 _09381_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[0][17] ), .ZN(_01803_ ) );
OAI211_X1 _09382_ ( .A(_01803_ ), .B(_01765_ ), .C1(_01775_ ), .C2(\myifu.myicache.tag[1][17] ), .ZN(_01804_ ) );
AND3_X2 _09383_ ( .A1(_01802_ ), .A2(\IF_ID_pc [22] ), .A3(_01804_ ), .ZN(_01805_ ) );
OR2_X4 _09384_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[0][21] ), .ZN(_01806_ ) );
OAI211_X1 _09385_ ( .A(_01806_ ), .B(_01765_ ), .C1(_01775_ ), .C2(\myifu.myicache.tag[1][21] ), .ZN(_01807_ ) );
OR2_X4 _09386_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[2][21] ), .ZN(_01808_ ) );
OAI211_X1 _09387_ ( .A(_01808_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01775_ ), .C2(\myifu.myicache.tag[3][21] ), .ZN(_01809_ ) );
AND3_X1 _09388_ ( .A1(_01807_ ), .A2(_01809_ ), .A3(\IF_ID_pc [26] ), .ZN(_01810_ ) );
AOI21_X1 _09389_ ( .A(\IF_ID_pc [26] ), .B1(_01807_ ), .B2(_01809_ ), .ZN(_01811_ ) );
NOR4_X1 _09390_ ( .A1(_01800_ ), .A2(_01805_ ), .A3(_01810_ ), .A4(_01811_ ), .ZN(_01812_ ) );
OR2_X1 _09391_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[0][19] ), .ZN(_01813_ ) );
OAI211_X1 _09392_ ( .A(_01813_ ), .B(_01798_ ), .C1(_01789_ ), .C2(\myifu.myicache.tag[1][19] ), .ZN(_01814_ ) );
OR2_X1 _09393_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[2][19] ), .ZN(_01815_ ) );
OAI211_X1 _09394_ ( .A(_01815_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01789_ ), .C2(\myifu.myicache.tag[3][19] ), .ZN(_01816_ ) );
INV_X1 _09395_ ( .A(\IF_ID_pc [24] ), .ZN(_01817_ ) );
AND3_X1 _09396_ ( .A1(_01814_ ), .A2(_01816_ ), .A3(_01817_ ), .ZN(_01818_ ) );
AOI21_X1 _09397_ ( .A(_01817_ ), .B1(_01814_ ), .B2(_01816_ ), .ZN(_01819_ ) );
OR2_X1 _09398_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[0][1] ), .ZN(_01820_ ) );
OAI211_X1 _09399_ ( .A(_01820_ ), .B(_01798_ ), .C1(_01789_ ), .C2(\myifu.myicache.tag[1][1] ), .ZN(_01821_ ) );
OR2_X1 _09400_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[2][1] ), .ZN(_01822_ ) );
OAI211_X1 _09401_ ( .A(_01822_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01789_ ), .C2(\myifu.myicache.tag[3][1] ), .ZN(_01823_ ) );
INV_X1 _09402_ ( .A(\IF_ID_pc [6] ), .ZN(_01824_ ) );
AND3_X1 _09403_ ( .A1(_01821_ ), .A2(_01823_ ), .A3(_01824_ ), .ZN(_01825_ ) );
AOI21_X1 _09404_ ( .A(_01824_ ), .B1(_01821_ ), .B2(_01823_ ), .ZN(_01826_ ) );
OAI221_X1 _09405_ ( .A(_01812_ ), .B1(_01818_ ), .B2(_01819_ ), .C1(_01825_ ), .C2(_01826_ ), .ZN(_01827_ ) );
OR2_X1 _09406_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[0][22] ), .ZN(_01828_ ) );
OAI211_X1 _09407_ ( .A(_01828_ ), .B(_01798_ ), .C1(_01789_ ), .C2(\myifu.myicache.tag[1][22] ), .ZN(_01829_ ) );
OR2_X1 _09408_ ( .A1(fanout_net_40 ), .A2(\myifu.myicache.tag[2][22] ), .ZN(_01830_ ) );
OAI211_X1 _09409_ ( .A(_01830_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01789_ ), .C2(\myifu.myicache.tag[3][22] ), .ZN(_01831_ ) );
AOI21_X1 _09410_ ( .A(\IF_ID_pc [27] ), .B1(_01829_ ), .B2(_01831_ ), .ZN(_01832_ ) );
MUX2_X1 _09411_ ( .A(\myifu.myicache.tag[0][20] ), .B(\myifu.myicache.tag[1][20] ), .S(fanout_net_40 ), .Z(_01833_ ) );
MUX2_X1 _09412_ ( .A(\myifu.myicache.tag[2][20] ), .B(\myifu.myicache.tag[3][20] ), .S(fanout_net_40 ), .Z(_01834_ ) );
MUX2_X1 _09413_ ( .A(_01833_ ), .B(_01834_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01835_ ) );
INV_X1 _09414_ ( .A(\IF_ID_pc [25] ), .ZN(_01836_ ) );
AOI21_X1 _09415_ ( .A(_01832_ ), .B1(_01835_ ), .B2(_01836_ ), .ZN(_01837_ ) );
MUX2_X1 _09416_ ( .A(\myifu.myicache.tag[0][24] ), .B(\myifu.myicache.tag[1][24] ), .S(fanout_net_40 ), .Z(_01838_ ) );
MUX2_X1 _09417_ ( .A(\myifu.myicache.tag[2][24] ), .B(\myifu.myicache.tag[3][24] ), .S(fanout_net_40 ), .Z(_01839_ ) );
MUX2_X1 _09418_ ( .A(_01838_ ), .B(_01839_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01840_ ) );
INV_X1 _09419_ ( .A(\IF_ID_pc [29] ), .ZN(_01841_ ) );
NAND2_X1 _09420_ ( .A1(_01840_ ), .A2(_01841_ ), .ZN(_01842_ ) );
INV_X1 _09421_ ( .A(\IF_ID_pc [21] ), .ZN(_01843_ ) );
MUX2_X1 _09422_ ( .A(\myifu.myicache.tag[0][16] ), .B(\myifu.myicache.tag[1][16] ), .S(fanout_net_40 ), .Z(_01844_ ) );
MUX2_X1 _09423_ ( .A(\myifu.myicache.tag[2][16] ), .B(\myifu.myicache.tag[3][16] ), .S(fanout_net_40 ), .Z(_01845_ ) );
MUX2_X1 _09424_ ( .A(_01844_ ), .B(_01845_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01846_ ) );
OAI211_X1 _09425_ ( .A(_01837_ ), .B(_01842_ ), .C1(_01843_ ), .C2(_01846_ ), .ZN(_01847_ ) );
AOI21_X1 _09426_ ( .A(\IF_ID_pc [22] ), .B1(_01802_ ), .B2(_01804_ ), .ZN(_01848_ ) );
AND3_X1 _09427_ ( .A1(_01829_ ), .A2(_01831_ ), .A3(\IF_ID_pc [27] ), .ZN(_01849_ ) );
NOR2_X1 _09428_ ( .A1(_01848_ ), .A2(_01849_ ), .ZN(_01850_ ) );
INV_X1 _09429_ ( .A(\IF_ID_pc [16] ), .ZN(_01851_ ) );
MUX2_X1 _09430_ ( .A(\myifu.myicache.tag[0][11] ), .B(\myifu.myicache.tag[1][11] ), .S(fanout_net_40 ), .Z(_01852_ ) );
MUX2_X1 _09431_ ( .A(\myifu.myicache.tag[2][11] ), .B(\myifu.myicache.tag[3][11] ), .S(fanout_net_40 ), .Z(_01853_ ) );
MUX2_X2 _09432_ ( .A(_01852_ ), .B(_01853_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01854_ ) );
MUX2_X1 _09433_ ( .A(\myifu.myicache.tag[0][13] ), .B(\myifu.myicache.tag[1][13] ), .S(fanout_net_40 ), .Z(_01855_ ) );
OR2_X1 _09434_ ( .A1(_01855_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01856_ ) );
MUX2_X1 _09435_ ( .A(\myifu.myicache.tag[2][13] ), .B(\myifu.myicache.tag[3][13] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01857_ ) );
OAI21_X1 _09436_ ( .A(_01856_ ), .B1(_01798_ ), .B2(_01857_ ), .ZN(_01858_ ) );
OAI221_X1 _09437_ ( .A(_01850_ ), .B1(_01851_ ), .B2(_01854_ ), .C1(\IF_ID_pc [18] ), .C2(_01858_ ), .ZN(_01859_ ) );
NOR4_X2 _09438_ ( .A1(_01795_ ), .A2(_01827_ ), .A3(_01847_ ), .A4(_01859_ ), .ZN(_01860_ ) );
MUX2_X1 _09439_ ( .A(\myifu.myicache.tag[0][8] ), .B(\myifu.myicache.tag[1][8] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01861_ ) );
MUX2_X1 _09440_ ( .A(\myifu.myicache.tag[2][8] ), .B(\myifu.myicache.tag[3][8] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01862_ ) );
MUX2_X1 _09441_ ( .A(_01861_ ), .B(_01862_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01863_ ) );
INV_X1 _09442_ ( .A(_01863_ ), .ZN(_01864_ ) );
AOI22_X1 _09443_ ( .A1(\IF_ID_pc [13] ), .A2(_01864_ ), .B1(_01858_ ), .B2(\IF_ID_pc [18] ), .ZN(_01865_ ) );
MUX2_X1 _09444_ ( .A(\myifu.myicache.tag[2][9] ), .B(\myifu.myicache.tag[3][9] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01866_ ) );
OR2_X1 _09445_ ( .A1(_01866_ ), .A2(_01798_ ), .ZN(_01867_ ) );
MUX2_X1 _09446_ ( .A(\myifu.myicache.tag[0][9] ), .B(\myifu.myicache.tag[1][9] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01868_ ) );
OAI21_X1 _09447_ ( .A(_01867_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01868_ ), .ZN(_01869_ ) );
MUX2_X1 _09448_ ( .A(\myifu.myicache.tag[2][15] ), .B(\myifu.myicache.tag[3][15] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01870_ ) );
AND2_X1 _09449_ ( .A1(_01870_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01871_ ) );
MUX2_X1 _09450_ ( .A(\myifu.myicache.tag[0][15] ), .B(\myifu.myicache.tag[1][15] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01872_ ) );
AOI21_X1 _09451_ ( .A(_01871_ ), .B1(_01798_ ), .B2(_01872_ ), .ZN(_01873_ ) );
OAI221_X1 _09452_ ( .A(_01865_ ), .B1(\IF_ID_pc [14] ), .B2(_01869_ ), .C1(\IF_ID_pc [20] ), .C2(_01873_ ), .ZN(_01874_ ) );
OR2_X1 _09453_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][0] ), .ZN(_01875_ ) );
OAI211_X1 _09454_ ( .A(_01875_ ), .B(_01765_ ), .C1(_01789_ ), .C2(\myifu.myicache.tag[1][0] ), .ZN(_01876_ ) );
OR2_X1 _09455_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][0] ), .ZN(_01877_ ) );
OAI211_X1 _09456_ ( .A(_01877_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01775_ ), .C2(\myifu.myicache.tag[3][0] ), .ZN(_01878_ ) );
NAND2_X1 _09457_ ( .A1(_01876_ ), .A2(_01878_ ), .ZN(_01879_ ) );
NOR2_X1 _09458_ ( .A1(_01879_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_01880_ ) );
MUX2_X1 _09459_ ( .A(\myifu.myicache.tag[2][26] ), .B(\myifu.myicache.tag[3][26] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01881_ ) );
OR2_X1 _09460_ ( .A1(_01881_ ), .A2(_01798_ ), .ZN(_01882_ ) );
MUX2_X1 _09461_ ( .A(\myifu.myicache.tag[0][26] ), .B(\myifu.myicache.tag[1][26] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01883_ ) );
OAI21_X1 _09462_ ( .A(_01882_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01883_ ), .ZN(_01884_ ) );
AOI21_X1 _09463_ ( .A(_01880_ ), .B1(_01884_ ), .B2(\IF_ID_pc [31] ), .ZN(_01885_ ) );
INV_X1 _09464_ ( .A(\IF_ID_pc [8] ), .ZN(_01886_ ) );
OR2_X1 _09465_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][3] ), .ZN(_01887_ ) );
OAI211_X1 _09466_ ( .A(_01887_ ), .B(_01798_ ), .C1(_01789_ ), .C2(\myifu.myicache.tag[1][3] ), .ZN(_01888_ ) );
AND2_X1 _09467_ ( .A1(_01775_ ), .A2(\myifu.myicache.tag[2][3] ), .ZN(_01889_ ) );
AOI21_X1 _09468_ ( .A(_01889_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myifu.myicache.tag[3][3] ), .ZN(_01890_ ) );
OAI21_X1 _09469_ ( .A(_01888_ ), .B1(_01890_ ), .B2(_01798_ ), .ZN(_01891_ ) );
OAI221_X1 _09470_ ( .A(_01885_ ), .B1(\IF_ID_pc [31] ), .B2(_01884_ ), .C1(_01886_ ), .C2(_01891_ ), .ZN(_01892_ ) );
INV_X1 _09471_ ( .A(\IF_ID_pc [12] ), .ZN(_01893_ ) );
MUX2_X1 _09472_ ( .A(\myifu.myicache.tag[0][7] ), .B(\myifu.myicache.tag[1][7] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01894_ ) );
MUX2_X1 _09473_ ( .A(\myifu.myicache.tag[2][7] ), .B(\myifu.myicache.tag[3][7] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01895_ ) );
MUX2_X2 _09474_ ( .A(_01894_ ), .B(_01895_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01896_ ) );
MUX2_X1 _09475_ ( .A(\myifu.myicache.tag[0][5] ), .B(\myifu.myicache.tag[1][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01897_ ) );
MUX2_X1 _09476_ ( .A(\myifu.myicache.tag[2][5] ), .B(\myifu.myicache.tag[3][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01898_ ) );
MUX2_X2 _09477_ ( .A(_01897_ ), .B(_01898_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01899_ ) );
INV_X1 _09478_ ( .A(\IF_ID_pc [10] ), .ZN(_01900_ ) );
AOI22_X1 _09479_ ( .A1(_01893_ ), .A2(_01896_ ), .B1(_01899_ ), .B2(_01900_ ), .ZN(_01901_ ) );
NAND2_X1 _09480_ ( .A1(_01891_ ), .A2(_01886_ ), .ZN(_01902_ ) );
OAI211_X1 _09481_ ( .A(_01901_ ), .B(_01902_ ), .C1(_01900_ ), .C2(_01899_ ), .ZN(_01903_ ) );
NAND2_X1 _09482_ ( .A1(_01854_ ), .A2(_01851_ ), .ZN(_01904_ ) );
OAI221_X1 _09483_ ( .A(_01904_ ), .B1(_01841_ ), .B2(_01840_ ), .C1(_01864_ ), .C2(\IF_ID_pc [13] ), .ZN(_01905_ ) );
NOR4_X2 _09484_ ( .A1(_01874_ ), .A2(_01892_ ), .A3(_01903_ ), .A4(_01905_ ), .ZN(_01906_ ) );
AOI22_X1 _09485_ ( .A1(_01873_ ), .A2(\IF_ID_pc [20] ), .B1(_01843_ ), .B2(_01846_ ), .ZN(_01907_ ) );
OR2_X1 _09486_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][4] ), .ZN(_01908_ ) );
OAI211_X1 _09487_ ( .A(_01908_ ), .B(_01765_ ), .C1(_01775_ ), .C2(\myifu.myicache.tag[1][4] ), .ZN(_01909_ ) );
OR2_X1 _09488_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][4] ), .ZN(_01910_ ) );
OAI211_X1 _09489_ ( .A(_01910_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01762_ ), .C2(\myifu.myicache.tag[3][4] ), .ZN(_01911_ ) );
NAND2_X1 _09490_ ( .A1(_01909_ ), .A2(_01911_ ), .ZN(_01912_ ) );
INV_X1 _09491_ ( .A(\IF_ID_pc [9] ), .ZN(_01913_ ) );
NAND2_X1 _09492_ ( .A1(_01912_ ), .A2(_01913_ ), .ZN(_01914_ ) );
INV_X1 _09493_ ( .A(\IF_ID_pc [23] ), .ZN(_01915_ ) );
MUX2_X1 _09494_ ( .A(\myifu.myicache.tag[0][18] ), .B(\myifu.myicache.tag[1][18] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01916_ ) );
MUX2_X1 _09495_ ( .A(\myifu.myicache.tag[2][18] ), .B(\myifu.myicache.tag[3][18] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01917_ ) );
MUX2_X2 _09496_ ( .A(_01916_ ), .B(_01917_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01918_ ) );
OAI211_X1 _09497_ ( .A(_01907_ ), .B(_01914_ ), .C1(_01915_ ), .C2(_01918_ ), .ZN(_01919_ ) );
AOI22_X1 _09498_ ( .A1(_01869_ ), .A2(\IF_ID_pc [14] ), .B1(_01915_ ), .B2(_01918_ ), .ZN(_01920_ ) );
NAND2_X1 _09499_ ( .A1(_01879_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_01921_ ) );
OAI211_X1 _09500_ ( .A(_01920_ ), .B(_01921_ ), .C1(_01893_ ), .C2(_01896_ ), .ZN(_01922_ ) );
NOR2_X1 _09501_ ( .A1(_01835_ ), .A2(_01836_ ), .ZN(_01923_ ) );
OR2_X4 _09502_ ( .A1(_01762_ ), .A2(\myifu.myicache.tag[1][12] ), .ZN(_01924_ ) );
OAI211_X2 _09503_ ( .A(_01924_ ), .B(_01765_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][12] ), .ZN(_01925_ ) );
OR2_X1 _09504_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][12] ), .ZN(_01926_ ) );
OAI211_X1 _09505_ ( .A(_01926_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01775_ ), .C2(\myifu.myicache.tag[3][12] ), .ZN(_01927_ ) );
AND3_X1 _09506_ ( .A1(_01925_ ), .A2(_01927_ ), .A3(\IF_ID_pc [17] ), .ZN(_01928_ ) );
OR2_X4 _09507_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][10] ), .ZN(_01929_ ) );
OAI211_X1 _09508_ ( .A(_01929_ ), .B(_01764_ ), .C1(_01762_ ), .C2(\myifu.myicache.tag[1][10] ), .ZN(_01930_ ) );
OR2_X4 _09509_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][10] ), .ZN(_01931_ ) );
OAI211_X1 _09510_ ( .A(_01931_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01762_ ), .C2(\myifu.myicache.tag[3][10] ), .ZN(_01932_ ) );
AND3_X1 _09511_ ( .A1(_01930_ ), .A2(_01932_ ), .A3(\IF_ID_pc [15] ), .ZN(_01933_ ) );
AOI21_X2 _09512_ ( .A(\IF_ID_pc [17] ), .B1(_01925_ ), .B2(_01927_ ), .ZN(_01934_ ) );
OR4_X4 _09513_ ( .A1(_01923_ ), .A2(_01928_ ), .A3(_01933_ ), .A4(_01934_ ), .ZN(_01935_ ) );
OR2_X4 _09514_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][2] ), .ZN(_01936_ ) );
OAI211_X2 _09515_ ( .A(_01936_ ), .B(_01765_ ), .C1(_01775_ ), .C2(\myifu.myicache.tag[1][2] ), .ZN(_01937_ ) );
OR2_X4 _09516_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][2] ), .ZN(_01938_ ) );
OAI211_X2 _09517_ ( .A(_01938_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01775_ ), .C2(\myifu.myicache.tag[3][2] ), .ZN(_01939_ ) );
AND3_X1 _09518_ ( .A1(_01937_ ), .A2(_01939_ ), .A3(\IF_ID_pc [7] ), .ZN(_01940_ ) );
AND3_X1 _09519_ ( .A1(_01909_ ), .A2(_01911_ ), .A3(\IF_ID_pc [9] ), .ZN(_01941_ ) );
AOI21_X1 _09520_ ( .A(\IF_ID_pc [15] ), .B1(_01930_ ), .B2(_01932_ ), .ZN(_01942_ ) );
AOI21_X1 _09521_ ( .A(\IF_ID_pc [7] ), .B1(_01937_ ), .B2(_01939_ ), .ZN(_01943_ ) );
OR4_X2 _09522_ ( .A1(_01940_ ), .A2(_01941_ ), .A3(_01942_ ), .A4(_01943_ ), .ZN(_01944_ ) );
NOR4_X4 _09523_ ( .A1(_01919_ ), .A2(_01922_ ), .A3(_01935_ ), .A4(_01944_ ), .ZN(_01945_ ) );
NAND3_X2 _09524_ ( .A1(_01860_ ), .A2(_01906_ ), .A3(_01945_ ), .ZN(_01946_ ) );
AND2_X4 _09525_ ( .A1(_01946_ ), .A2(\myifu.state [0] ), .ZN(_01947_ ) );
INV_X2 _09526_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01948_ ) );
NOR2_X4 _09527_ ( .A1(_01947_ ), .A2(_01948_ ), .ZN(_01949_ ) );
NOR2_X1 _09528_ ( .A1(\myminixbar.state [2] ), .A2(\myminixbar.state [0] ), .ZN(_01950_ ) );
NOR2_X4 _09529_ ( .A1(_01949_ ), .A2(_01950_ ), .ZN(_01951_ ) );
INV_X32 _09530_ ( .A(\EX_LS_flag [2] ), .ZN(_01952_ ) );
NAND4_X1 _09531_ ( .A1(_01952_ ), .A2(\EX_LS_flag [1] ), .A3(\EX_LS_flag [0] ), .A4(EXU_valid_LSU ), .ZN(_01953_ ) );
NOR2_X1 _09532_ ( .A1(_01953_ ), .A2(fanout_net_42 ), .ZN(_01954_ ) );
INV_X1 _09533_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ), .ZN(_01955_ ) );
NOR2_X1 _09534_ ( .A1(_01954_ ), .A2(_01955_ ), .ZN(_01956_ ) );
NOR2_X4 _09535_ ( .A1(_01951_ ), .A2(_01956_ ), .ZN(_01957_ ) );
BUF_X8 _09536_ ( .A(_01957_ ), .Z(_01958_ ) );
CLKBUF_X2 _09537_ ( .A(_01953_ ), .Z(_01959_ ) );
OR3_X1 _09538_ ( .A1(_01959_ ), .A2(\EX_LS_dest_csreg_mem [21] ), .A3(fanout_net_42 ), .ZN(_01960_ ) );
BUF_X4 _09539_ ( .A(_01954_ ), .Z(_01961_ ) );
OAI211_X1 _09540_ ( .A(_01958_ ), .B(_01960_ ), .C1(\mylsu.araddr_tmp [21] ), .C2(_01961_ ), .ZN(_01962_ ) );
INV_X4 _09541_ ( .A(_01951_ ), .ZN(_01963_ ) );
OAI21_X1 _09542_ ( .A(_01962_ ), .B1(_01843_ ), .B2(_01963_ ), .ZN(\io_master_araddr [21] ) );
OR3_X1 _09543_ ( .A1(_01953_ ), .A2(\EX_LS_dest_csreg_mem [29] ), .A3(fanout_net_42 ), .ZN(_01964_ ) );
OAI211_X1 _09544_ ( .A(_01957_ ), .B(_01964_ ), .C1(\mylsu.araddr_tmp [29] ), .C2(_01954_ ), .ZN(_01965_ ) );
OAI21_X1 _09545_ ( .A(_01965_ ), .B1(_01841_ ), .B2(_01963_ ), .ZN(\io_master_araddr [29] ) );
CLKBUF_X2 _09546_ ( .A(_01957_ ), .Z(_01966_ ) );
CLKBUF_X2 _09547_ ( .A(_01959_ ), .Z(_01967_ ) );
OR3_X1 _09548_ ( .A1(_01967_ ), .A2(\EX_LS_dest_csreg_mem [20] ), .A3(fanout_net_42 ), .ZN(_01968_ ) );
BUF_X4 _09549_ ( .A(_01961_ ), .Z(_01969_ ) );
OAI211_X1 _09550_ ( .A(_01966_ ), .B(_01968_ ), .C1(\mylsu.araddr_tmp [20] ), .C2(_01969_ ), .ZN(_01970_ ) );
INV_X1 _09551_ ( .A(\IF_ID_pc [20] ), .ZN(_01971_ ) );
BUF_X4 _09552_ ( .A(_01963_ ), .Z(_01972_ ) );
OAI21_X1 _09553_ ( .A(_01970_ ), .B1(_01971_ ), .B2(_01972_ ), .ZN(\io_master_araddr [20] ) );
OR3_X1 _09554_ ( .A1(_01959_ ), .A2(\EX_LS_dest_csreg_mem [18] ), .A3(fanout_net_42 ), .ZN(_01973_ ) );
OAI211_X1 _09555_ ( .A(_01958_ ), .B(_01973_ ), .C1(\mylsu.araddr_tmp [18] ), .C2(_01969_ ), .ZN(_01974_ ) );
INV_X1 _09556_ ( .A(\IF_ID_pc [18] ), .ZN(_01975_ ) );
OAI21_X1 _09557_ ( .A(_01974_ ), .B1(_01975_ ), .B2(_01972_ ), .ZN(\io_master_araddr [18] ) );
OR4_X1 _09558_ ( .A1(\io_master_araddr [21] ), .A2(\io_master_araddr [29] ), .A3(\io_master_araddr [20] ), .A4(\io_master_araddr [18] ), .ZN(_01976_ ) );
OR3_X1 _09559_ ( .A1(_01959_ ), .A2(\EX_LS_dest_csreg_mem [23] ), .A3(fanout_net_42 ), .ZN(_01977_ ) );
OAI211_X1 _09560_ ( .A(_01958_ ), .B(_01977_ ), .C1(\mylsu.araddr_tmp [23] ), .C2(_01961_ ), .ZN(_01978_ ) );
OAI21_X1 _09561_ ( .A(_01978_ ), .B1(_01915_ ), .B2(_01963_ ), .ZN(\io_master_araddr [23] ) );
OR3_X1 _09562_ ( .A1(_01959_ ), .A2(\EX_LS_dest_csreg_mem [17] ), .A3(fanout_net_42 ), .ZN(_01979_ ) );
OAI211_X1 _09563_ ( .A(_01958_ ), .B(_01979_ ), .C1(\mylsu.araddr_tmp [17] ), .C2(_01961_ ), .ZN(_01980_ ) );
INV_X1 _09564_ ( .A(\IF_ID_pc [17] ), .ZN(_01981_ ) );
OAI21_X1 _09565_ ( .A(_01980_ ), .B1(_01981_ ), .B2(_01963_ ), .ZN(\io_master_araddr [17] ) );
OR3_X1 _09566_ ( .A1(_01959_ ), .A2(\EX_LS_dest_csreg_mem [19] ), .A3(fanout_net_42 ), .ZN(_01982_ ) );
OAI211_X1 _09567_ ( .A(_01958_ ), .B(_01982_ ), .C1(\mylsu.araddr_tmp [19] ), .C2(_01961_ ), .ZN(_01983_ ) );
OAI221_X1 _09568_ ( .A(\IF_ID_pc [19] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01947_ ), .C2(_01948_ ), .ZN(_01984_ ) );
AND2_X1 _09569_ ( .A1(_01983_ ), .A2(_01984_ ), .ZN(_01985_ ) );
INV_X1 _09570_ ( .A(EXU_valid_LSU ), .ZN(_01986_ ) );
NOR2_X1 _09571_ ( .A1(_01986_ ), .A2(fanout_net_42 ), .ZN(_01987_ ) );
INV_X1 _09572_ ( .A(\EX_LS_dest_csreg_mem [25] ), .ZN(_01988_ ) );
AND2_X4 _09573_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_01989_ ) );
NAND4_X1 _09574_ ( .A1(_01987_ ), .A2(_01988_ ), .A3(_01989_ ), .A4(_01952_ ), .ZN(_01990_ ) );
OAI211_X4 _09575_ ( .A(_01958_ ), .B(_01990_ ), .C1(\mylsu.araddr_tmp [25] ), .C2(_01961_ ), .ZN(_01991_ ) );
OAI21_X4 _09576_ ( .A(_01991_ ), .B1(_01836_ ), .B2(_01963_ ), .ZN(\io_master_araddr [25] ) );
NAND2_X1 _09577_ ( .A1(_01985_ ), .A2(\io_master_araddr [25] ), .ZN(_01992_ ) );
OR4_X1 _09578_ ( .A1(_01976_ ), .A2(\io_master_araddr [23] ), .A3(\io_master_araddr [17] ), .A4(_01992_ ), .ZN(_01993_ ) );
INV_X1 _09579_ ( .A(\EX_LS_dest_csreg_mem [24] ), .ZN(_01994_ ) );
NAND4_X1 _09580_ ( .A1(_01987_ ), .A2(_01994_ ), .A3(_01989_ ), .A4(_01952_ ), .ZN(_01995_ ) );
OAI211_X1 _09581_ ( .A(_01957_ ), .B(_01995_ ), .C1(\mylsu.araddr_tmp [24] ), .C2(_01961_ ), .ZN(_01996_ ) );
OAI221_X1 _09582_ ( .A(\IF_ID_pc [24] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01947_ ), .C2(_01948_ ), .ZN(_01997_ ) );
AND2_X1 _09583_ ( .A1(_01996_ ), .A2(_01997_ ), .ZN(_01998_ ) );
INV_X1 _09584_ ( .A(_01998_ ), .ZN(\io_master_araddr [24] ) );
OR3_X1 _09585_ ( .A1(_01967_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(fanout_net_42 ), .ZN(_01999_ ) );
OAI211_X1 _09586_ ( .A(_01958_ ), .B(_01999_ ), .C1(\mylsu.araddr_tmp [27] ), .C2(_01969_ ), .ZN(_02000_ ) );
INV_X1 _09587_ ( .A(\IF_ID_pc [27] ), .ZN(_02001_ ) );
OAI21_X1 _09588_ ( .A(_02000_ ), .B1(_02001_ ), .B2(_01972_ ), .ZN(\io_master_araddr [27] ) );
OR3_X1 _09589_ ( .A1(_01959_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(fanout_net_42 ), .ZN(_02002_ ) );
OAI211_X1 _09590_ ( .A(_01958_ ), .B(_02002_ ), .C1(\mylsu.araddr_tmp [26] ), .C2(_01961_ ), .ZN(_02003_ ) );
INV_X1 _09591_ ( .A(\IF_ID_pc [26] ), .ZN(_02004_ ) );
OAI21_X1 _09592_ ( .A(_02003_ ), .B1(_02004_ ), .B2(_01963_ ), .ZN(\io_master_araddr [26] ) );
OR3_X1 _09593_ ( .A1(_01967_ ), .A2(\EX_LS_dest_csreg_mem [22] ), .A3(fanout_net_42 ), .ZN(_02005_ ) );
OAI211_X1 _09594_ ( .A(_01958_ ), .B(_02005_ ), .C1(\mylsu.araddr_tmp [22] ), .C2(_01969_ ), .ZN(_02006_ ) );
INV_X1 _09595_ ( .A(\IF_ID_pc [22] ), .ZN(_02007_ ) );
OAI21_X1 _09596_ ( .A(_02006_ ), .B1(_02007_ ), .B2(_01972_ ), .ZN(\io_master_araddr [22] ) );
NOR4_X1 _09597_ ( .A1(\io_master_araddr [24] ), .A2(\io_master_araddr [27] ), .A3(\io_master_araddr [26] ), .A4(\io_master_araddr [22] ), .ZN(_02008_ ) );
OR3_X1 _09598_ ( .A1(_01959_ ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(fanout_net_42 ), .ZN(_02009_ ) );
OAI211_X1 _09599_ ( .A(_01957_ ), .B(_02009_ ), .C1(\mylsu.araddr_tmp [30] ), .C2(_01954_ ), .ZN(_02010_ ) );
OAI21_X1 _09600_ ( .A(_02010_ ), .B1(_01770_ ), .B2(_01963_ ), .ZN(\io_master_araddr [30] ) );
OR3_X1 _09601_ ( .A1(_01959_ ), .A2(\EX_LS_dest_csreg_mem [16] ), .A3(fanout_net_42 ), .ZN(_02011_ ) );
OAI211_X1 _09602_ ( .A(_01958_ ), .B(_02011_ ), .C1(\mylsu.araddr_tmp [16] ), .C2(_01961_ ), .ZN(_02012_ ) );
OAI21_X1 _09603_ ( .A(_02012_ ), .B1(_01851_ ), .B2(_01963_ ), .ZN(\io_master_araddr [16] ) );
OR3_X1 _09604_ ( .A1(_01953_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(fanout_net_42 ), .ZN(_02013_ ) );
OAI211_X1 _09605_ ( .A(_01957_ ), .B(_02013_ ), .C1(\mylsu.araddr_tmp [28] ), .C2(_01954_ ), .ZN(_02014_ ) );
OAI21_X1 _09606_ ( .A(_02014_ ), .B1(_01777_ ), .B2(_01963_ ), .ZN(\io_master_araddr [28] ) );
OR3_X1 _09607_ ( .A1(_01959_ ), .A2(\EX_LS_dest_csreg_mem [31] ), .A3(fanout_net_42 ), .ZN(_02015_ ) );
OAI211_X1 _09608_ ( .A(_01957_ ), .B(_02015_ ), .C1(\mylsu.araddr_tmp [31] ), .C2(_01961_ ), .ZN(_02016_ ) );
OAI221_X1 _09609_ ( .A(\IF_ID_pc [31] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01947_ ), .C2(_01948_ ), .ZN(_02017_ ) );
NAND2_X1 _09610_ ( .A1(_02016_ ), .A2(_02017_ ), .ZN(\io_master_araddr [31] ) );
NOR4_X1 _09611_ ( .A1(\io_master_araddr [30] ), .A2(\io_master_araddr [16] ), .A3(\io_master_araddr [28] ), .A4(\io_master_araddr [31] ), .ZN(_02018_ ) );
NAND2_X1 _09612_ ( .A1(_02008_ ), .A2(_02018_ ), .ZN(_02019_ ) );
CLKBUF_X2 _09613_ ( .A(_01951_ ), .Z(_02020_ ) );
CLKBUF_X2 _09614_ ( .A(_02020_ ), .Z(_02021_ ) );
CLKBUF_X2 _09615_ ( .A(_02021_ ), .Z(_02022_ ) );
AND2_X4 _09616_ ( .A1(_01989_ ), .A2(_01952_ ), .ZN(_02023_ ) );
NOR2_X1 _09617_ ( .A1(fanout_net_3 ), .A2(fanout_net_4 ), .ZN(_02024_ ) );
INV_X1 _09618_ ( .A(_02024_ ), .ZN(_02025_ ) );
INV_X1 _09619_ ( .A(\EX_LS_typ [1] ), .ZN(_02026_ ) );
INV_X1 _09620_ ( .A(\EX_LS_typ [3] ), .ZN(_02027_ ) );
NAND4_X1 _09621_ ( .A1(_02025_ ), .A2(_02026_ ), .A3(_02027_ ), .A4(\EX_LS_typ [2] ), .ZN(_02028_ ) );
AND2_X1 _09622_ ( .A1(fanout_net_3 ), .A2(\EX_LS_typ [1] ), .ZN(_02029_ ) );
NOR2_X1 _09623_ ( .A1(\EX_LS_typ [3] ), .A2(\EX_LS_typ [2] ), .ZN(_02030_ ) );
NAND2_X1 _09624_ ( .A1(_02029_ ), .A2(_02030_ ), .ZN(_02031_ ) );
AOI21_X1 _09625_ ( .A(\EX_LS_typ [0] ), .B1(_02028_ ), .B2(_02031_ ), .ZN(_02032_ ) );
AND3_X1 _09626_ ( .A1(_02029_ ), .A2(\EX_LS_typ [0] ), .A3(_02030_ ), .ZN(_02033_ ) );
OAI21_X1 _09627_ ( .A(_02023_ ), .B1(_02032_ ), .B2(_02033_ ), .ZN(_02034_ ) );
OR2_X1 _09628_ ( .A1(_02034_ ), .A2(\EX_LS_typ [4] ), .ZN(_02035_ ) );
NAND2_X1 _09629_ ( .A1(_01994_ ), .A2(_01988_ ), .ZN(_02036_ ) );
NOR3_X1 _09630_ ( .A1(_02036_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(\EX_LS_dest_csreg_mem [26] ), .ZN(_02037_ ) );
NOR4_X1 _09631_ ( .A1(\EX_LS_dest_csreg_mem [31] ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(\EX_LS_dest_csreg_mem [29] ), .A4(\EX_LS_dest_csreg_mem [28] ), .ZN(_02038_ ) );
AND2_X1 _09632_ ( .A1(_02037_ ), .A2(_02038_ ), .ZN(_02039_ ) );
NAND2_X1 _09633_ ( .A1(_02039_ ), .A2(_02023_ ), .ZN(_02040_ ) );
NAND2_X1 _09634_ ( .A1(_02035_ ), .A2(_02040_ ), .ZN(_02041_ ) );
INV_X32 _09635_ ( .A(\EX_LS_flag [1] ), .ZN(_02042_ ) );
NOR2_X4 _09636_ ( .A1(_02042_ ), .A2(\EX_LS_flag [0] ), .ZN(_02043_ ) );
BUF_X4 _09637_ ( .A(_02043_ ), .Z(_02044_ ) );
AND2_X2 _09638_ ( .A1(_02044_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02045_ ) );
AND2_X1 _09639_ ( .A1(_02039_ ), .A2(_02045_ ), .ZN(_02046_ ) );
NAND2_X1 _09640_ ( .A1(\EX_LS_typ [2] ), .A2(\EX_LS_typ [0] ), .ZN(_02047_ ) );
NOR3_X1 _09641_ ( .A1(_02047_ ), .A2(_02026_ ), .A3(_02027_ ), .ZN(_02048_ ) );
BUF_X4 _09642_ ( .A(_01952_ ), .Z(_02049_ ) );
NOR3_X1 _09643_ ( .A1(_02042_ ), .A2(\EX_LS_typ [4] ), .A3(\EX_LS_flag [0] ), .ZN(_02050_ ) );
NAND4_X1 _09644_ ( .A1(_02048_ ), .A2(_02049_ ), .A3(_02025_ ), .A4(_02050_ ), .ZN(_02051_ ) );
AND3_X1 _09645_ ( .A1(_02030_ ), .A2(\EX_LS_typ [1] ), .A3(\EX_LS_typ [0] ), .ZN(_02052_ ) );
NAND4_X1 _09646_ ( .A1(_02052_ ), .A2(fanout_net_3 ), .A3(_02049_ ), .A4(_02050_ ), .ZN(_02053_ ) );
NAND2_X1 _09647_ ( .A1(_02051_ ), .A2(_02053_ ), .ZN(_02054_ ) );
NOR2_X1 _09648_ ( .A1(_02046_ ), .A2(_02054_ ), .ZN(_02055_ ) );
INV_X1 _09649_ ( .A(_02055_ ), .ZN(_02056_ ) );
NOR2_X1 _09650_ ( .A1(_02041_ ), .A2(_02056_ ), .ZN(_02057_ ) );
AOI21_X1 _09651_ ( .A(_02022_ ), .B1(_01969_ ), .B2(_02057_ ), .ZN(_02058_ ) );
NOR2_X1 _09652_ ( .A1(fanout_net_2 ), .A2(\myidu.stall_quest_fencei ), .ZN(_02059_ ) );
AOI211_X1 _09653_ ( .A(_01950_ ), .B(_01949_ ), .C1(\myifu.state [0] ), .C2(_02059_ ), .ZN(_02060_ ) );
NOR4_X1 _09654_ ( .A1(_01993_ ), .A2(_02019_ ), .A3(_02058_ ), .A4(_02060_ ), .ZN(_02061_ ) );
OAI21_X1 _09655_ ( .A(_01592_ ), .B1(_02061_ ), .B2(\myclint.rvalid ), .ZN(_02062_ ) );
OR4_X2 _09656_ ( .A1(\io_master_araddr [31] ), .A2(\io_master_araddr [30] ), .A3(\io_master_araddr [28] ), .A4(\io_master_araddr [29] ), .ZN(_02063_ ) );
NAND2_X4 _09657_ ( .A1(_01998_ ), .A2(\io_master_araddr [25] ), .ZN(_02064_ ) );
NOR4_X4 _09658_ ( .A1(_02063_ ), .A2(\io_master_araddr [27] ), .A3(\io_master_araddr [26] ), .A4(_02064_ ), .ZN(_02065_ ) );
INV_X1 _09659_ ( .A(_01985_ ), .ZN(\io_master_araddr [19] ) );
NOR4_X1 _09660_ ( .A1(\io_master_araddr [19] ), .A2(\io_master_araddr [22] ), .A3(\io_master_araddr [16] ), .A4(\io_master_araddr [21] ), .ZN(_02066_ ) );
NOR4_X1 _09661_ ( .A1(\io_master_araddr [20] ), .A2(\io_master_araddr [18] ), .A3(\io_master_araddr [23] ), .A4(\io_master_araddr [17] ), .ZN(_02067_ ) );
AND2_X1 _09662_ ( .A1(_02066_ ), .A2(_02067_ ), .ZN(_02068_ ) );
NAND3_X1 _09663_ ( .A1(_02065_ ), .A2(\myclint.rvalid ), .A3(_02068_ ), .ZN(_02069_ ) );
AOI211_X1 _09664_ ( .A(_01955_ ), .B(_02022_ ), .C1(_01969_ ), .C2(_02057_ ), .ZN(_02070_ ) );
AND3_X1 _09665_ ( .A1(_01946_ ), .A2(\myifu.state [0] ), .A3(_02059_ ), .ZN(_02071_ ) );
NOR4_X1 _09666_ ( .A1(_01949_ ), .A2(_01948_ ), .A3(_01950_ ), .A4(_02071_ ), .ZN(_02072_ ) );
NOR3_X1 _09667_ ( .A1(_02069_ ), .A2(_02070_ ), .A3(_02072_ ), .ZN(_02073_ ) );
NOR2_X1 _09668_ ( .A1(_02062_ ), .A2(_02073_ ), .ZN(_00064_ ) );
INV_X1 _09669_ ( .A(\LS_WB_wen_csreg [6] ), .ZN(_02074_ ) );
CLKBUF_X2 _09670_ ( .A(_02074_ ), .Z(_02075_ ) );
AND2_X1 _09671_ ( .A1(_02075_ ), .A2(\LS_WB_wdata_csreg [31] ), .ZN(_00065_ ) );
AND2_X1 _09672_ ( .A1(_02075_ ), .A2(\LS_WB_wdata_csreg [30] ), .ZN(_00066_ ) );
AND2_X1 _09673_ ( .A1(_02075_ ), .A2(\LS_WB_wdata_csreg [21] ), .ZN(_00067_ ) );
AND2_X1 _09674_ ( .A1(_02075_ ), .A2(\LS_WB_wdata_csreg [20] ), .ZN(_00068_ ) );
AND2_X1 _09675_ ( .A1(_02075_ ), .A2(\LS_WB_wdata_csreg [19] ), .ZN(_00069_ ) );
AND2_X1 _09676_ ( .A1(_02075_ ), .A2(\LS_WB_wdata_csreg [18] ), .ZN(_00070_ ) );
AND2_X1 _09677_ ( .A1(_02075_ ), .A2(\LS_WB_wdata_csreg [17] ), .ZN(_00071_ ) );
AND2_X1 _09678_ ( .A1(_02075_ ), .A2(\LS_WB_wdata_csreg [16] ), .ZN(_00072_ ) );
AND2_X1 _09679_ ( .A1(_02075_ ), .A2(\LS_WB_wdata_csreg [15] ), .ZN(_00073_ ) );
AND2_X1 _09680_ ( .A1(_02075_ ), .A2(\LS_WB_wdata_csreg [14] ), .ZN(_00074_ ) );
CLKBUF_X2 _09681_ ( .A(_02074_ ), .Z(_02076_ ) );
AND2_X1 _09682_ ( .A1(_02076_ ), .A2(\LS_WB_wdata_csreg [13] ), .ZN(_00075_ ) );
AND2_X1 _09683_ ( .A1(_02076_ ), .A2(\LS_WB_wdata_csreg [12] ), .ZN(_00076_ ) );
AND2_X1 _09684_ ( .A1(_02076_ ), .A2(\LS_WB_wdata_csreg [29] ), .ZN(_00077_ ) );
INV_X1 _09685_ ( .A(\LS_WB_wdata_csreg [11] ), .ZN(_02077_ ) );
NOR2_X1 _09686_ ( .A1(_02077_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00078_ ) );
AND2_X1 _09687_ ( .A1(_02076_ ), .A2(\LS_WB_wdata_csreg [10] ), .ZN(_00079_ ) );
AND2_X1 _09688_ ( .A1(_02076_ ), .A2(\LS_WB_wdata_csreg [9] ), .ZN(_00080_ ) );
AND2_X1 _09689_ ( .A1(_02076_ ), .A2(\LS_WB_wdata_csreg [8] ), .ZN(_00081_ ) );
AND2_X1 _09690_ ( .A1(_02076_ ), .A2(\LS_WB_wdata_csreg [7] ), .ZN(_00082_ ) );
AND2_X1 _09691_ ( .A1(_02076_ ), .A2(\LS_WB_wdata_csreg [6] ), .ZN(_00083_ ) );
AND2_X1 _09692_ ( .A1(_02076_ ), .A2(\LS_WB_wdata_csreg [5] ), .ZN(_00084_ ) );
AND2_X1 _09693_ ( .A1(_02076_ ), .A2(\LS_WB_wdata_csreg [4] ), .ZN(_00085_ ) );
AND2_X1 _09694_ ( .A1(_02074_ ), .A2(\LS_WB_wdata_csreg [28] ), .ZN(_00086_ ) );
AND2_X1 _09695_ ( .A1(_02074_ ), .A2(\LS_WB_wdata_csreg [27] ), .ZN(_00087_ ) );
AND2_X1 _09696_ ( .A1(_02074_ ), .A2(\LS_WB_wdata_csreg [26] ), .ZN(_00088_ ) );
AND2_X1 _09697_ ( .A1(_02074_ ), .A2(\LS_WB_wdata_csreg [25] ), .ZN(_00089_ ) );
AND2_X1 _09698_ ( .A1(_02074_ ), .A2(\LS_WB_wdata_csreg [24] ), .ZN(_00090_ ) );
AND2_X1 _09699_ ( .A1(_02074_ ), .A2(\LS_WB_wdata_csreg [23] ), .ZN(_00091_ ) );
INV_X1 _09700_ ( .A(\LS_WB_wdata_csreg [22] ), .ZN(_02078_ ) );
NOR2_X1 _09701_ ( .A1(_02078_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00092_ ) );
BUF_X2 _09702_ ( .A(_02056_ ), .Z(_02079_ ) );
NOR2_X1 _09703_ ( .A1(\myec.state [0] ), .A2(\myec.state [1] ), .ZN(_02080_ ) );
NAND2_X1 _09704_ ( .A1(_02080_ ), .A2(_01548_ ), .ZN(_02081_ ) );
OR2_X1 _09705_ ( .A1(\myexu.pc_jump [27] ), .A2(\myexu.pc_jump [24] ), .ZN(_02082_ ) );
OR3_X1 _09706_ ( .A1(_02082_ ), .A2(\myexu.pc_jump [26] ), .A3(\myexu.pc_jump [25] ), .ZN(_02083_ ) );
OR4_X1 _09707_ ( .A1(\myexu.pc_jump [31] ), .A2(\myexu.pc_jump [30] ), .A3(\myexu.pc_jump [29] ), .A4(\myexu.pc_jump [28] ), .ZN(_02084_ ) );
NOR2_X1 _09708_ ( .A1(_02083_ ), .A2(_02084_ ), .ZN(_02085_ ) );
NOR2_X1 _09709_ ( .A1(\myexu.pc_jump [0] ), .A2(\myexu.pc_jump [1] ), .ZN(_02086_ ) );
INV_X1 _09710_ ( .A(_02086_ ), .ZN(_02087_ ) );
NOR3_X1 _09711_ ( .A1(_02085_ ), .A2(exception_quest_IDU ), .A3(_02087_ ), .ZN(_02088_ ) );
NOR4_X1 _09712_ ( .A1(_02041_ ), .A2(_02079_ ), .A3(_02081_ ), .A4(_02088_ ), .ZN(_00094_ ) );
AOI21_X1 _09713_ ( .A(_02081_ ), .B1(_02057_ ), .B2(exception_quest_IDU ), .ZN(_00095_ ) );
AND3_X1 _09714_ ( .A1(_02042_ ), .A2(\EX_LS_flag [0] ), .A3(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02089_ ) );
AND2_X1 _09715_ ( .A1(_02042_ ), .A2(\EX_LS_flag [0] ), .ZN(_02090_ ) );
AOI211_X2 _09716_ ( .A(_02089_ ), .B(_02023_ ), .C1(\EX_LS_flag [2] ), .C2(_02090_ ), .ZN(_02091_ ) );
AND2_X1 _09717_ ( .A1(_02043_ ), .A2(\EX_LS_flag [2] ), .ZN(_02092_ ) );
INV_X1 _09718_ ( .A(_02092_ ), .ZN(_02093_ ) );
NAND2_X4 _09719_ ( .A1(_02091_ ), .A2(_02093_ ), .ZN(_02094_ ) );
XNOR2_X1 _09720_ ( .A(\ID_EX_rs1 [0] ), .B(\EX_LS_dest_reg [0] ), .ZN(_02095_ ) );
OR3_X1 _09721_ ( .A1(\EX_LS_dest_reg [2] ), .A2(\EX_LS_dest_reg [1] ), .A3(\EX_LS_dest_reg [0] ), .ZN(_02096_ ) );
OR2_X1 _09722_ ( .A1(\EX_LS_dest_reg [4] ), .A2(\EX_LS_dest_reg [3] ), .ZN(_02097_ ) );
NOR2_X1 _09723_ ( .A1(_02096_ ), .A2(_02097_ ), .ZN(_02098_ ) );
INV_X1 _09724_ ( .A(_02098_ ), .ZN(_02099_ ) );
INV_X8 _09725_ ( .A(\EX_LS_dest_reg [1] ), .ZN(_02100_ ) );
NAND2_X1 _09726_ ( .A1(_02100_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_02101_ ) );
NAND4_X4 _09727_ ( .A1(_02094_ ), .A2(_02095_ ), .A3(_02099_ ), .A4(_02101_ ), .ZN(_02102_ ) );
BUF_X8 _09728_ ( .A(_02102_ ), .Z(_02103_ ) );
BUF_X2 _09729_ ( .A(_02103_ ), .Z(_02104_ ) );
BUF_X8 _09730_ ( .A(_02104_ ), .Z(_02105_ ) );
XOR2_X1 _09731_ ( .A(\ID_EX_rs1 [4] ), .B(\EX_LS_dest_reg [4] ), .Z(_02106_ ) );
XOR2_X2 _09732_ ( .A(\ID_EX_rs1 [2] ), .B(\EX_LS_dest_reg [2] ), .Z(_02107_ ) );
INV_X1 _09733_ ( .A(\ID_EX_rs1 [3] ), .ZN(_02108_ ) );
OAI22_X1 _09734_ ( .A1(_02108_ ), .A2(\EX_LS_dest_reg [3] ), .B1(_02100_ ), .B2(\ID_EX_rs1 [1] ), .ZN(_02109_ ) );
INV_X1 _09735_ ( .A(\EX_LS_dest_reg [3] ), .ZN(_02110_ ) );
OAI21_X1 _09736_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .B1(_02110_ ), .B2(\ID_EX_rs1 [3] ), .ZN(_02111_ ) );
OR4_X4 _09737_ ( .A1(_02106_ ), .A2(_02107_ ), .A3(_02109_ ), .A4(_02111_ ), .ZN(_02112_ ) );
BUF_X8 _09738_ ( .A(_02112_ ), .Z(_02113_ ) );
BUF_X8 _09739_ ( .A(_02113_ ), .Z(_02114_ ) );
BUF_X8 _09740_ ( .A(_02114_ ), .Z(_02115_ ) );
OR3_X1 _09741_ ( .A1(_02105_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02115_ ), .ZN(_02116_ ) );
INV_X1 _09742_ ( .A(fanout_net_27 ), .ZN(_02117_ ) );
BUF_X4 _09743_ ( .A(_02117_ ), .Z(_02118_ ) );
BUF_X4 _09744_ ( .A(_02118_ ), .Z(_02119_ ) );
BUF_X4 _09745_ ( .A(_02119_ ), .Z(_02120_ ) );
INV_X1 _09746_ ( .A(fanout_net_15 ), .ZN(_02121_ ) );
CLKBUF_X2 _09747_ ( .A(_02121_ ), .Z(_02122_ ) );
CLKBUF_X3 _09748_ ( .A(_02122_ ), .Z(_02123_ ) );
CLKBUF_X3 _09749_ ( .A(_02123_ ), .Z(_02124_ ) );
OR2_X1 _09750_ ( .A1(_02124_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02125_ ) );
INV_X1 _09751_ ( .A(fanout_net_23 ), .ZN(_02126_ ) );
BUF_X4 _09752_ ( .A(_02126_ ), .Z(_02127_ ) );
BUF_X4 _09753_ ( .A(_02127_ ), .Z(_02128_ ) );
BUF_X4 _09754_ ( .A(_02128_ ), .Z(_02129_ ) );
BUF_X4 _09755_ ( .A(_02129_ ), .Z(_02130_ ) );
OAI211_X1 _09756_ ( .A(_02125_ ), .B(_02130_ ), .C1(fanout_net_15 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02131_ ) );
INV_X1 _09757_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02132_ ) );
NAND2_X1 _09758_ ( .A1(_02132_ ), .A2(fanout_net_15 ), .ZN(_02133_ ) );
OAI211_X1 _09759_ ( .A(_02133_ ), .B(fanout_net_23 ), .C1(fanout_net_15 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02134_ ) );
INV_X2 _09760_ ( .A(fanout_net_26 ), .ZN(_02135_ ) );
BUF_X4 _09761_ ( .A(_02135_ ), .Z(_02136_ ) );
BUF_X4 _09762_ ( .A(_02136_ ), .Z(_02137_ ) );
BUF_X4 _09763_ ( .A(_02137_ ), .Z(_02138_ ) );
NAND3_X1 _09764_ ( .A1(_02131_ ), .A2(_02134_ ), .A3(_02138_ ), .ZN(_02139_ ) );
MUX2_X1 _09765_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02140_ ) );
MUX2_X1 _09766_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02141_ ) );
BUF_X4 _09767_ ( .A(_02127_ ), .Z(_02142_ ) );
BUF_X4 _09768_ ( .A(_02142_ ), .Z(_02143_ ) );
BUF_X4 _09769_ ( .A(_02143_ ), .Z(_02144_ ) );
MUX2_X1 _09770_ ( .A(_02140_ ), .B(_02141_ ), .S(_02144_ ), .Z(_02145_ ) );
BUF_X4 _09771_ ( .A(_02136_ ), .Z(_02146_ ) );
BUF_X4 _09772_ ( .A(_02146_ ), .Z(_02147_ ) );
OAI211_X1 _09773_ ( .A(_02120_ ), .B(_02139_ ), .C1(_02145_ ), .C2(_02147_ ), .ZN(_02148_ ) );
OR2_X1 _09774_ ( .A1(_02124_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02149_ ) );
OAI211_X1 _09775_ ( .A(_02149_ ), .B(_02130_ ), .C1(fanout_net_15 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02150_ ) );
OR2_X1 _09776_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02151_ ) );
BUF_X2 _09777_ ( .A(_02123_ ), .Z(_02152_ ) );
BUF_X2 _09778_ ( .A(_02152_ ), .Z(_02153_ ) );
OAI211_X1 _09779_ ( .A(_02151_ ), .B(fanout_net_23 ), .C1(_02153_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02154_ ) );
NAND3_X1 _09780_ ( .A1(_02150_ ), .A2(fanout_net_26 ), .A3(_02154_ ), .ZN(_02155_ ) );
MUX2_X1 _09781_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02156_ ) );
MUX2_X1 _09782_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02157_ ) );
MUX2_X1 _09783_ ( .A(_02156_ ), .B(_02157_ ), .S(fanout_net_23 ), .Z(_02158_ ) );
OAI211_X1 _09784_ ( .A(fanout_net_27 ), .B(_02155_ ), .C1(_02158_ ), .C2(fanout_net_26 ), .ZN(_02159_ ) );
BUF_X8 _09785_ ( .A(_02102_ ), .Z(_02160_ ) );
BUF_X2 _09786_ ( .A(_02160_ ), .Z(_02161_ ) );
BUF_X2 _09787_ ( .A(_02161_ ), .Z(_02162_ ) );
CLKBUF_X2 _09788_ ( .A(_02112_ ), .Z(_02163_ ) );
BUF_X2 _09789_ ( .A(_02163_ ), .Z(_02164_ ) );
BUF_X2 _09790_ ( .A(_02164_ ), .Z(_02165_ ) );
OAI211_X1 _09791_ ( .A(_02148_ ), .B(_02159_ ), .C1(_02162_ ), .C2(_02165_ ), .ZN(_02166_ ) );
NAND2_X2 _09792_ ( .A1(_02116_ ), .A2(_02166_ ), .ZN(_02167_ ) );
XNOR2_X1 _09793_ ( .A(_02167_ ), .B(\ID_EX_imm [28] ), .ZN(_02168_ ) );
CLKBUF_X2 _09794_ ( .A(_02121_ ), .Z(_02169_ ) );
CLKBUF_X2 _09795_ ( .A(_02169_ ), .Z(_02170_ ) );
BUF_X2 _09796_ ( .A(_02170_ ), .Z(_02171_ ) );
OR2_X1 _09797_ ( .A1(_02171_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02172_ ) );
BUF_X4 _09798_ ( .A(_02127_ ), .Z(_02173_ ) );
BUF_X4 _09799_ ( .A(_02173_ ), .Z(_02174_ ) );
BUF_X4 _09800_ ( .A(_02174_ ), .Z(_02175_ ) );
BUF_X4 _09801_ ( .A(_02175_ ), .Z(_02176_ ) );
OAI211_X1 _09802_ ( .A(_02172_ ), .B(_02176_ ), .C1(fanout_net_15 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02177_ ) );
OR2_X1 _09803_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02178_ ) );
BUF_X4 _09804_ ( .A(_02171_ ), .Z(_02179_ ) );
OAI211_X1 _09805_ ( .A(_02178_ ), .B(fanout_net_23 ), .C1(_02179_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02180_ ) );
NAND3_X1 _09806_ ( .A1(_02177_ ), .A2(fanout_net_26 ), .A3(_02180_ ), .ZN(_02181_ ) );
MUX2_X1 _09807_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02182_ ) );
MUX2_X1 _09808_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02183_ ) );
MUX2_X1 _09809_ ( .A(_02182_ ), .B(_02183_ ), .S(_02176_ ), .Z(_02184_ ) );
OAI211_X1 _09810_ ( .A(_02120_ ), .B(_02181_ ), .C1(_02184_ ), .C2(fanout_net_26 ), .ZN(_02185_ ) );
MUX2_X1 _09811_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02186_ ) );
AND2_X1 _09812_ ( .A1(_02186_ ), .A2(fanout_net_23 ), .ZN(_02187_ ) );
MUX2_X1 _09813_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02188_ ) );
AOI211_X1 _09814_ ( .A(fanout_net_26 ), .B(_02187_ ), .C1(_02176_ ), .C2(_02188_ ), .ZN(_02189_ ) );
MUX2_X1 _09815_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02190_ ) );
MUX2_X1 _09816_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02191_ ) );
MUX2_X1 _09817_ ( .A(_02190_ ), .B(_02191_ ), .S(fanout_net_23 ), .Z(_02192_ ) );
OAI21_X1 _09818_ ( .A(fanout_net_27 ), .B1(_02192_ ), .B2(_02147_ ), .ZN(_02193_ ) );
OAI221_X1 _09819_ ( .A(_02185_ ), .B1(_02189_ ), .B2(_02193_ ), .C1(_02162_ ), .C2(_02165_ ), .ZN(_02194_ ) );
OR3_X1 _09820_ ( .A1(_02105_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02115_ ), .ZN(_02195_ ) );
NAND2_X1 _09821_ ( .A1(_02194_ ), .A2(_02195_ ), .ZN(_02196_ ) );
INV_X1 _09822_ ( .A(\ID_EX_imm [26] ), .ZN(_02197_ ) );
XNOR2_X1 _09823_ ( .A(_02196_ ), .B(_02197_ ), .ZN(_02198_ ) );
OR3_X1 _09824_ ( .A1(_02105_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02115_ ), .ZN(_02199_ ) );
INV_X1 _09825_ ( .A(\ID_EX_imm [27] ), .ZN(_02200_ ) );
OR2_X1 _09826_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02201_ ) );
OAI211_X1 _09827_ ( .A(_02201_ ), .B(_02130_ ), .C1(_02153_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02202_ ) );
OR2_X1 _09828_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02203_ ) );
OAI211_X1 _09829_ ( .A(_02203_ ), .B(fanout_net_23 ), .C1(_02153_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02204_ ) );
NAND3_X1 _09830_ ( .A1(_02202_ ), .A2(_02204_ ), .A3(fanout_net_26 ), .ZN(_02205_ ) );
MUX2_X1 _09831_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02206_ ) );
MUX2_X1 _09832_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02207_ ) );
MUX2_X1 _09833_ ( .A(_02206_ ), .B(_02207_ ), .S(_02144_ ), .Z(_02208_ ) );
OAI211_X1 _09834_ ( .A(_02120_ ), .B(_02205_ ), .C1(_02208_ ), .C2(fanout_net_26 ), .ZN(_02209_ ) );
NOR2_X1 _09835_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02210_ ) );
OAI21_X1 _09836_ ( .A(_02144_ ), .B1(_02171_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02211_ ) );
INV_X1 _09837_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02212_ ) );
INV_X1 _09838_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02213_ ) );
MUX2_X1 _09839_ ( .A(_02212_ ), .B(_02213_ ), .S(fanout_net_15 ), .Z(_02214_ ) );
OAI221_X1 _09840_ ( .A(_02138_ ), .B1(_02210_ ), .B2(_02211_ ), .C1(_02214_ ), .C2(_02176_ ), .ZN(_02215_ ) );
MUX2_X1 _09841_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02216_ ) );
MUX2_X1 _09842_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02217_ ) );
MUX2_X1 _09843_ ( .A(_02216_ ), .B(_02217_ ), .S(fanout_net_23 ), .Z(_02218_ ) );
OAI211_X1 _09844_ ( .A(fanout_net_27 ), .B(_02215_ ), .C1(_02218_ ), .C2(_02147_ ), .ZN(_02219_ ) );
OAI211_X1 _09845_ ( .A(_02209_ ), .B(_02219_ ), .C1(_02162_ ), .C2(_02165_ ), .ZN(_02220_ ) );
AND3_X1 _09846_ ( .A1(_02199_ ), .A2(_02200_ ), .A3(_02220_ ), .ZN(_02221_ ) );
AOI21_X1 _09847_ ( .A(_02200_ ), .B1(_02199_ ), .B2(_02220_ ), .ZN(_02222_ ) );
NOR2_X1 _09848_ ( .A1(_02221_ ), .A2(_02222_ ), .ZN(_02223_ ) );
AND2_X1 _09849_ ( .A1(_02198_ ), .A2(_02223_ ), .ZN(_02224_ ) );
OR3_X1 _09850_ ( .A1(_02161_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02164_ ), .ZN(_02225_ ) );
BUF_X2 _09851_ ( .A(_02122_ ), .Z(_02226_ ) );
BUF_X2 _09852_ ( .A(_02226_ ), .Z(_02227_ ) );
OR2_X1 _09853_ ( .A1(_02227_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02228_ ) );
OAI211_X1 _09854_ ( .A(_02228_ ), .B(_02175_ ), .C1(fanout_net_15 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02229_ ) );
OR2_X1 _09855_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02230_ ) );
OAI211_X1 _09856_ ( .A(_02230_ ), .B(fanout_net_23 ), .C1(_02171_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02231_ ) );
NAND3_X1 _09857_ ( .A1(_02229_ ), .A2(_02146_ ), .A3(_02231_ ), .ZN(_02232_ ) );
MUX2_X1 _09858_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02233_ ) );
MUX2_X1 _09859_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02234_ ) );
MUX2_X1 _09860_ ( .A(_02233_ ), .B(_02234_ ), .S(_02175_ ), .Z(_02235_ ) );
OAI211_X1 _09861_ ( .A(_02119_ ), .B(_02232_ ), .C1(_02235_ ), .C2(_02138_ ), .ZN(_02236_ ) );
OR2_X1 _09862_ ( .A1(_02227_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02237_ ) );
OAI211_X1 _09863_ ( .A(_02237_ ), .B(fanout_net_23 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02238_ ) );
OR2_X1 _09864_ ( .A1(_02227_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02239_ ) );
OAI211_X1 _09865_ ( .A(_02239_ ), .B(_02175_ ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02240_ ) );
NAND3_X1 _09866_ ( .A1(_02238_ ), .A2(_02240_ ), .A3(fanout_net_26 ), .ZN(_02241_ ) );
MUX2_X1 _09867_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02242_ ) );
MUX2_X1 _09868_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02243_ ) );
MUX2_X1 _09869_ ( .A(_02242_ ), .B(_02243_ ), .S(fanout_net_23 ), .Z(_02244_ ) );
OAI211_X1 _09870_ ( .A(fanout_net_27 ), .B(_02241_ ), .C1(_02244_ ), .C2(fanout_net_26 ), .ZN(_02245_ ) );
OAI211_X1 _09871_ ( .A(_02236_ ), .B(_02245_ ), .C1(_02105_ ), .C2(_02115_ ), .ZN(_02246_ ) );
NAND2_X2 _09872_ ( .A1(_02225_ ), .A2(_02246_ ), .ZN(_02247_ ) );
INV_X1 _09873_ ( .A(\ID_EX_imm [23] ), .ZN(_02248_ ) );
XNOR2_X1 _09874_ ( .A(_02247_ ), .B(_02248_ ), .ZN(_02249_ ) );
OR3_X1 _09875_ ( .A1(_02105_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02115_ ), .ZN(_02250_ ) );
OR2_X1 _09876_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02251_ ) );
OAI211_X1 _09877_ ( .A(_02251_ ), .B(_02176_ ), .C1(_02179_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02252_ ) );
OR2_X1 _09878_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02253_ ) );
OAI211_X1 _09879_ ( .A(_02253_ ), .B(fanout_net_23 ), .C1(_02179_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02254_ ) );
NAND3_X1 _09880_ ( .A1(_02252_ ), .A2(_02254_ ), .A3(fanout_net_26 ), .ZN(_02255_ ) );
MUX2_X1 _09881_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02256_ ) );
MUX2_X1 _09882_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02257_ ) );
MUX2_X1 _09883_ ( .A(_02256_ ), .B(_02257_ ), .S(_02176_ ), .Z(_02258_ ) );
OAI211_X1 _09884_ ( .A(_02120_ ), .B(_02255_ ), .C1(_02258_ ), .C2(fanout_net_26 ), .ZN(_02259_ ) );
NOR2_X1 _09885_ ( .A1(_02179_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02260_ ) );
OAI21_X1 _09886_ ( .A(fanout_net_23 ), .B1(fanout_net_16 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02261_ ) );
NOR2_X1 _09887_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02262_ ) );
OAI21_X1 _09888_ ( .A(_02130_ ), .B1(_02179_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02263_ ) );
OAI221_X1 _09889_ ( .A(_02138_ ), .B1(_02260_ ), .B2(_02261_ ), .C1(_02262_ ), .C2(_02263_ ), .ZN(_02264_ ) );
MUX2_X1 _09890_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02265_ ) );
MUX2_X1 _09891_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02266_ ) );
MUX2_X1 _09892_ ( .A(_02265_ ), .B(_02266_ ), .S(fanout_net_23 ), .Z(_02267_ ) );
OAI211_X1 _09893_ ( .A(fanout_net_27 ), .B(_02264_ ), .C1(_02267_ ), .C2(_02147_ ), .ZN(_02268_ ) );
OAI211_X1 _09894_ ( .A(_02259_ ), .B(_02268_ ), .C1(_02162_ ), .C2(_02165_ ), .ZN(_02269_ ) );
NAND2_X2 _09895_ ( .A1(_02250_ ), .A2(_02269_ ), .ZN(_02270_ ) );
INV_X1 _09896_ ( .A(\ID_EX_imm [22] ), .ZN(_02271_ ) );
XNOR2_X1 _09897_ ( .A(_02270_ ), .B(_02271_ ), .ZN(_02272_ ) );
AND2_X1 _09898_ ( .A1(_02249_ ), .A2(_02272_ ), .ZN(_02273_ ) );
OR3_X4 _09899_ ( .A1(_02105_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02115_ ), .ZN(_02274_ ) );
OR2_X1 _09900_ ( .A1(_02171_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02275_ ) );
OAI211_X1 _09901_ ( .A(_02275_ ), .B(_02176_ ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02276_ ) );
OR2_X1 _09902_ ( .A1(_02171_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02277_ ) );
OAI211_X1 _09903_ ( .A(_02277_ ), .B(fanout_net_23 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02278_ ) );
NAND3_X1 _09904_ ( .A1(_02276_ ), .A2(_02278_ ), .A3(_02138_ ), .ZN(_02279_ ) );
MUX2_X1 _09905_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02280_ ) );
MUX2_X1 _09906_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02281_ ) );
MUX2_X1 _09907_ ( .A(_02280_ ), .B(_02281_ ), .S(_02130_ ), .Z(_02282_ ) );
OAI211_X1 _09908_ ( .A(fanout_net_27 ), .B(_02279_ ), .C1(_02282_ ), .C2(_02147_ ), .ZN(_02283_ ) );
OR2_X1 _09909_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02284_ ) );
OAI211_X1 _09910_ ( .A(_02284_ ), .B(_02130_ ), .C1(_02153_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02285_ ) );
NOR2_X1 _09911_ ( .A1(_02179_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02286_ ) );
OAI21_X1 _09912_ ( .A(fanout_net_23 ), .B1(fanout_net_16 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02287_ ) );
OAI211_X1 _09913_ ( .A(_02285_ ), .B(_02138_ ), .C1(_02286_ ), .C2(_02287_ ), .ZN(_02288_ ) );
MUX2_X1 _09914_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02289_ ) );
MUX2_X1 _09915_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02290_ ) );
MUX2_X1 _09916_ ( .A(_02289_ ), .B(_02290_ ), .S(_02130_ ), .Z(_02291_ ) );
OAI211_X1 _09917_ ( .A(_02120_ ), .B(_02288_ ), .C1(_02291_ ), .C2(_02147_ ), .ZN(_02292_ ) );
OAI211_X1 _09918_ ( .A(_02283_ ), .B(_02292_ ), .C1(_02162_ ), .C2(_02165_ ), .ZN(_02293_ ) );
NAND2_X2 _09919_ ( .A1(_02274_ ), .A2(_02293_ ), .ZN(_02294_ ) );
INV_X1 _09920_ ( .A(\ID_EX_imm [20] ), .ZN(_02295_ ) );
XNOR2_X1 _09921_ ( .A(_02294_ ), .B(_02295_ ), .ZN(_02296_ ) );
OR3_X1 _09922_ ( .A1(_02105_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02115_ ), .ZN(_02297_ ) );
INV_X1 _09923_ ( .A(\ID_EX_imm [21] ), .ZN(_02298_ ) );
OR2_X1 _09924_ ( .A1(_02171_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02299_ ) );
OAI211_X1 _09925_ ( .A(_02299_ ), .B(fanout_net_23 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02300_ ) );
OR2_X1 _09926_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02301_ ) );
OAI211_X1 _09927_ ( .A(_02301_ ), .B(_02130_ ), .C1(_02179_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02302_ ) );
NAND3_X1 _09928_ ( .A1(_02300_ ), .A2(fanout_net_26 ), .A3(_02302_ ), .ZN(_02303_ ) );
MUX2_X1 _09929_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02304_ ) );
MUX2_X1 _09930_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02305_ ) );
MUX2_X1 _09931_ ( .A(_02304_ ), .B(_02305_ ), .S(_02144_ ), .Z(_02306_ ) );
OAI211_X1 _09932_ ( .A(_02120_ ), .B(_02303_ ), .C1(_02306_ ), .C2(fanout_net_26 ), .ZN(_02307_ ) );
NOR2_X1 _09933_ ( .A1(_02153_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02308_ ) );
OAI21_X1 _09934_ ( .A(fanout_net_23 ), .B1(fanout_net_16 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02309_ ) );
NOR2_X1 _09935_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02310_ ) );
OAI21_X1 _09936_ ( .A(_02144_ ), .B1(_02153_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02311_ ) );
OAI221_X1 _09937_ ( .A(_02138_ ), .B1(_02308_ ), .B2(_02309_ ), .C1(_02310_ ), .C2(_02311_ ), .ZN(_02312_ ) );
MUX2_X1 _09938_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02313_ ) );
MUX2_X1 _09939_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02314_ ) );
MUX2_X1 _09940_ ( .A(_02313_ ), .B(_02314_ ), .S(fanout_net_23 ), .Z(_02315_ ) );
OAI211_X1 _09941_ ( .A(fanout_net_27 ), .B(_02312_ ), .C1(_02315_ ), .C2(_02147_ ), .ZN(_02316_ ) );
OAI211_X1 _09942_ ( .A(_02307_ ), .B(_02316_ ), .C1(_02162_ ), .C2(_02165_ ), .ZN(_02317_ ) );
AND3_X1 _09943_ ( .A1(_02297_ ), .A2(_02298_ ), .A3(_02317_ ), .ZN(_02318_ ) );
AOI21_X1 _09944_ ( .A(_02298_ ), .B1(_02297_ ), .B2(_02317_ ), .ZN(_02319_ ) );
NOR2_X1 _09945_ ( .A1(_02318_ ), .A2(_02319_ ), .ZN(_02320_ ) );
AND2_X1 _09946_ ( .A1(_02296_ ), .A2(_02320_ ), .ZN(_02321_ ) );
AND2_X1 _09947_ ( .A1(_02273_ ), .A2(_02321_ ), .ZN(_02322_ ) );
INV_X1 _09948_ ( .A(_02322_ ), .ZN(_02323_ ) );
OR3_X1 _09949_ ( .A1(_02160_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02163_ ), .ZN(_02324_ ) );
OR2_X1 _09950_ ( .A1(_02123_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02325_ ) );
OAI211_X1 _09951_ ( .A(_02325_ ), .B(fanout_net_23 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02326_ ) );
BUF_X4 _09952_ ( .A(_02135_ ), .Z(_02327_ ) );
BUF_X4 _09953_ ( .A(_02327_ ), .Z(_02328_ ) );
OR2_X1 _09954_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02329_ ) );
OAI211_X1 _09955_ ( .A(_02329_ ), .B(_02174_ ), .C1(_02227_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02330_ ) );
NAND3_X1 _09956_ ( .A1(_02326_ ), .A2(_02328_ ), .A3(_02330_ ), .ZN(_02331_ ) );
MUX2_X1 _09957_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02332_ ) );
MUX2_X1 _09958_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02333_ ) );
MUX2_X1 _09959_ ( .A(_02332_ ), .B(_02333_ ), .S(_02174_ ), .Z(_02334_ ) );
OAI211_X1 _09960_ ( .A(_02118_ ), .B(_02331_ ), .C1(_02334_ ), .C2(_02137_ ), .ZN(_02335_ ) );
OR2_X1 _09961_ ( .A1(_02123_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02336_ ) );
OAI211_X1 _09962_ ( .A(_02336_ ), .B(fanout_net_23 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02337_ ) );
OR2_X1 _09963_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02338_ ) );
OAI211_X1 _09964_ ( .A(_02338_ ), .B(_02174_ ), .C1(_02227_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02339_ ) );
NAND3_X1 _09965_ ( .A1(_02337_ ), .A2(fanout_net_26 ), .A3(_02339_ ), .ZN(_02340_ ) );
MUX2_X1 _09966_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02341_ ) );
MUX2_X1 _09967_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02342_ ) );
MUX2_X1 _09968_ ( .A(_02341_ ), .B(_02342_ ), .S(fanout_net_23 ), .Z(_02343_ ) );
OAI211_X1 _09969_ ( .A(fanout_net_27 ), .B(_02340_ ), .C1(_02343_ ), .C2(fanout_net_26 ), .ZN(_02344_ ) );
OAI211_X1 _09970_ ( .A(_02335_ ), .B(_02344_ ), .C1(_02104_ ), .C2(_02114_ ), .ZN(_02345_ ) );
NAND2_X2 _09971_ ( .A1(_02324_ ), .A2(_02345_ ), .ZN(_02346_ ) );
INV_X1 _09972_ ( .A(\ID_EX_imm [18] ), .ZN(_02347_ ) );
XNOR2_X1 _09973_ ( .A(_02346_ ), .B(_02347_ ), .ZN(_02348_ ) );
OR3_X1 _09974_ ( .A1(_02160_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02163_ ), .ZN(_02349_ ) );
CLKBUF_X2 _09975_ ( .A(_02169_ ), .Z(_02350_ ) );
OR2_X1 _09976_ ( .A1(_02350_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02351_ ) );
OAI211_X1 _09977_ ( .A(_02351_ ), .B(fanout_net_23 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02352_ ) );
OR2_X1 _09978_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02353_ ) );
OAI211_X1 _09979_ ( .A(_02353_ ), .B(_02143_ ), .C1(_02152_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02354_ ) );
NAND3_X1 _09980_ ( .A1(_02352_ ), .A2(_02328_ ), .A3(_02354_ ), .ZN(_02355_ ) );
MUX2_X1 _09981_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02356_ ) );
MUX2_X1 _09982_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02357_ ) );
MUX2_X1 _09983_ ( .A(_02356_ ), .B(_02357_ ), .S(_02174_ ), .Z(_02358_ ) );
OAI211_X1 _09984_ ( .A(_02119_ ), .B(_02355_ ), .C1(_02358_ ), .C2(_02137_ ), .ZN(_02359_ ) );
OR2_X1 _09985_ ( .A1(_02123_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02360_ ) );
OAI211_X1 _09986_ ( .A(_02360_ ), .B(fanout_net_23 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02361_ ) );
OR2_X1 _09987_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02362_ ) );
OAI211_X1 _09988_ ( .A(_02362_ ), .B(_02143_ ), .C1(_02152_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02363_ ) );
NAND3_X1 _09989_ ( .A1(_02361_ ), .A2(fanout_net_26 ), .A3(_02363_ ), .ZN(_02364_ ) );
MUX2_X1 _09990_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02365_ ) );
MUX2_X1 _09991_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02366_ ) );
MUX2_X1 _09992_ ( .A(_02365_ ), .B(_02366_ ), .S(fanout_net_23 ), .Z(_02367_ ) );
OAI211_X1 _09993_ ( .A(fanout_net_27 ), .B(_02364_ ), .C1(_02367_ ), .C2(fanout_net_26 ), .ZN(_02368_ ) );
OAI211_X2 _09994_ ( .A(_02359_ ), .B(_02368_ ), .C1(_02104_ ), .C2(_02114_ ), .ZN(_02369_ ) );
NAND2_X2 _09995_ ( .A1(_02349_ ), .A2(_02369_ ), .ZN(_02370_ ) );
INV_X1 _09996_ ( .A(\ID_EX_imm [19] ), .ZN(_02371_ ) );
XNOR2_X1 _09997_ ( .A(_02370_ ), .B(_02371_ ), .ZN(_02372_ ) );
AND2_X1 _09998_ ( .A1(_02348_ ), .A2(_02372_ ), .ZN(_02373_ ) );
OR3_X1 _09999_ ( .A1(_02104_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02114_ ), .ZN(_02374_ ) );
OR2_X1 _10000_ ( .A1(_02350_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02375_ ) );
OAI211_X1 _10001_ ( .A(_02375_ ), .B(fanout_net_23 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02376_ ) );
OR2_X1 _10002_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02377_ ) );
OAI211_X1 _10003_ ( .A(_02377_ ), .B(_02129_ ), .C1(_02152_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02378_ ) );
NAND3_X1 _10004_ ( .A1(_02376_ ), .A2(_02328_ ), .A3(_02378_ ), .ZN(_02379_ ) );
MUX2_X1 _10005_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02380_ ) );
MUX2_X1 _10006_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02381_ ) );
MUX2_X1 _10007_ ( .A(_02380_ ), .B(_02381_ ), .S(_02143_ ), .Z(_02382_ ) );
OAI211_X1 _10008_ ( .A(_02119_ ), .B(_02379_ ), .C1(_02382_ ), .C2(_02146_ ), .ZN(_02383_ ) );
OR2_X1 _10009_ ( .A1(_02350_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02384_ ) );
OAI211_X1 _10010_ ( .A(_02384_ ), .B(fanout_net_23 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02385_ ) );
OR2_X1 _10011_ ( .A1(_02350_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02386_ ) );
OAI211_X1 _10012_ ( .A(_02386_ ), .B(_02129_ ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02387_ ) );
NAND3_X1 _10013_ ( .A1(_02385_ ), .A2(_02387_ ), .A3(fanout_net_26 ), .ZN(_02388_ ) );
MUX2_X1 _10014_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02389_ ) );
MUX2_X1 _10015_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02390_ ) );
MUX2_X1 _10016_ ( .A(_02389_ ), .B(_02390_ ), .S(fanout_net_23 ), .Z(_02391_ ) );
OAI211_X1 _10017_ ( .A(fanout_net_27 ), .B(_02388_ ), .C1(_02391_ ), .C2(fanout_net_26 ), .ZN(_02392_ ) );
OAI211_X1 _10018_ ( .A(_02383_ ), .B(_02392_ ), .C1(_02161_ ), .C2(_02164_ ), .ZN(_02393_ ) );
NAND2_X4 _10019_ ( .A1(_02374_ ), .A2(_02393_ ), .ZN(_02394_ ) );
INV_X1 _10020_ ( .A(\ID_EX_imm [17] ), .ZN(_02395_ ) );
XNOR2_X1 _10021_ ( .A(_02394_ ), .B(_02395_ ), .ZN(_02396_ ) );
OR3_X1 _10022_ ( .A1(_02161_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02164_ ), .ZN(_02397_ ) );
OR2_X1 _10023_ ( .A1(_02124_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02398_ ) );
OAI211_X1 _10024_ ( .A(_02398_ ), .B(_02144_ ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02399_ ) );
OR2_X1 _10025_ ( .A1(_02152_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02400_ ) );
OAI211_X1 _10026_ ( .A(_02400_ ), .B(fanout_net_23 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02401_ ) );
NAND3_X1 _10027_ ( .A1(_02399_ ), .A2(_02401_ ), .A3(fanout_net_26 ), .ZN(_02402_ ) );
MUX2_X1 _10028_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02403_ ) );
MUX2_X1 _10029_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02404_ ) );
MUX2_X1 _10030_ ( .A(_02403_ ), .B(_02404_ ), .S(_02144_ ), .Z(_02405_ ) );
OAI211_X1 _10031_ ( .A(_02120_ ), .B(_02402_ ), .C1(_02405_ ), .C2(fanout_net_26 ), .ZN(_02406_ ) );
NOR2_X1 _10032_ ( .A1(_02171_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02407_ ) );
OAI21_X1 _10033_ ( .A(fanout_net_24 ), .B1(fanout_net_17 ), .B2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02408_ ) );
NOR2_X1 _10034_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02409_ ) );
OAI21_X1 _10035_ ( .A(_02144_ ), .B1(_02171_ ), .B2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02410_ ) );
OAI221_X1 _10036_ ( .A(_02146_ ), .B1(_02407_ ), .B2(_02408_ ), .C1(_02409_ ), .C2(_02410_ ), .ZN(_02411_ ) );
MUX2_X1 _10037_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02412_ ) );
MUX2_X1 _10038_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02413_ ) );
MUX2_X1 _10039_ ( .A(_02412_ ), .B(_02413_ ), .S(fanout_net_24 ), .Z(_02414_ ) );
OAI211_X1 _10040_ ( .A(fanout_net_27 ), .B(_02411_ ), .C1(_02414_ ), .C2(_02138_ ), .ZN(_02415_ ) );
OAI211_X1 _10041_ ( .A(_02406_ ), .B(_02415_ ), .C1(_02105_ ), .C2(_02115_ ), .ZN(_02416_ ) );
NAND2_X2 _10042_ ( .A1(_02397_ ), .A2(_02416_ ), .ZN(_02417_ ) );
INV_X1 _10043_ ( .A(\ID_EX_imm [16] ), .ZN(_02418_ ) );
XNOR2_X1 _10044_ ( .A(_02417_ ), .B(_02418_ ), .ZN(_02419_ ) );
NAND3_X1 _10045_ ( .A1(_02373_ ), .A2(_02396_ ), .A3(_02419_ ), .ZN(_02420_ ) );
OR3_X1 _10046_ ( .A1(_02102_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02112_ ), .ZN(_02421_ ) );
OR2_X1 _10047_ ( .A1(_02122_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02422_ ) );
OAI211_X1 _10048_ ( .A(_02422_ ), .B(_02173_ ), .C1(fanout_net_18 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02423_ ) );
OR2_X1 _10049_ ( .A1(fanout_net_18 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02424_ ) );
OAI211_X1 _10050_ ( .A(_02424_ ), .B(fanout_net_24 ), .C1(_02226_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02425_ ) );
NAND3_X1 _10051_ ( .A1(_02423_ ), .A2(_02327_ ), .A3(_02425_ ), .ZN(_02426_ ) );
MUX2_X1 _10052_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02427_ ) );
MUX2_X1 _10053_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02428_ ) );
MUX2_X1 _10054_ ( .A(_02427_ ), .B(_02428_ ), .S(_02127_ ), .Z(_02429_ ) );
OAI211_X1 _10055_ ( .A(_02117_ ), .B(_02426_ ), .C1(_02429_ ), .C2(_02327_ ), .ZN(_02430_ ) );
OR2_X1 _10056_ ( .A1(_02122_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02431_ ) );
OAI211_X1 _10057_ ( .A(_02431_ ), .B(fanout_net_24 ), .C1(fanout_net_18 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02432_ ) );
OR2_X1 _10058_ ( .A1(_02122_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02433_ ) );
OAI211_X1 _10059_ ( .A(_02433_ ), .B(_02127_ ), .C1(fanout_net_18 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02434_ ) );
NAND3_X1 _10060_ ( .A1(_02432_ ), .A2(_02434_ ), .A3(fanout_net_26 ), .ZN(_02435_ ) );
MUX2_X1 _10061_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02436_ ) );
MUX2_X1 _10062_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02437_ ) );
MUX2_X1 _10063_ ( .A(_02436_ ), .B(_02437_ ), .S(fanout_net_24 ), .Z(_02438_ ) );
OAI211_X1 _10064_ ( .A(fanout_net_27 ), .B(_02435_ ), .C1(_02438_ ), .C2(fanout_net_26 ), .ZN(_02439_ ) );
OAI211_X1 _10065_ ( .A(_02430_ ), .B(_02439_ ), .C1(_02103_ ), .C2(_02113_ ), .ZN(_02440_ ) );
NAND2_X2 _10066_ ( .A1(_02421_ ), .A2(_02440_ ), .ZN(_02441_ ) );
INV_X1 _10067_ ( .A(\ID_EX_imm [2] ), .ZN(_02442_ ) );
XNOR2_X1 _10068_ ( .A(_02441_ ), .B(_02442_ ), .ZN(_02443_ ) );
OR3_X4 _10069_ ( .A1(_02102_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02112_ ), .ZN(_02444_ ) );
OR2_X1 _10070_ ( .A1(_02121_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02445_ ) );
OAI211_X1 _10071_ ( .A(_02445_ ), .B(_02126_ ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02446_ ) );
OR2_X1 _10072_ ( .A1(_02121_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02447_ ) );
OAI211_X1 _10073_ ( .A(_02447_ ), .B(fanout_net_24 ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02448_ ) );
NAND3_X1 _10074_ ( .A1(_02446_ ), .A2(_02448_ ), .A3(_02135_ ), .ZN(_02449_ ) );
MUX2_X1 _10075_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02450_ ) );
MUX2_X1 _10076_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02451_ ) );
MUX2_X1 _10077_ ( .A(_02450_ ), .B(_02451_ ), .S(_02126_ ), .Z(_02452_ ) );
OAI211_X1 _10078_ ( .A(fanout_net_27 ), .B(_02449_ ), .C1(_02452_ ), .C2(_02135_ ), .ZN(_02453_ ) );
OR2_X1 _10079_ ( .A1(_02121_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02454_ ) );
OAI211_X1 _10080_ ( .A(_02454_ ), .B(_02126_ ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02455_ ) );
OR2_X1 _10081_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02456_ ) );
OAI211_X1 _10082_ ( .A(_02456_ ), .B(fanout_net_24 ), .C1(_02121_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02457_ ) );
NAND3_X1 _10083_ ( .A1(_02455_ ), .A2(_02135_ ), .A3(_02457_ ), .ZN(_02458_ ) );
MUX2_X1 _10084_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02459_ ) );
MUX2_X1 _10085_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02460_ ) );
MUX2_X1 _10086_ ( .A(_02459_ ), .B(_02460_ ), .S(_02126_ ), .Z(_02461_ ) );
OAI211_X1 _10087_ ( .A(_02117_ ), .B(_02458_ ), .C1(_02461_ ), .C2(_02135_ ), .ZN(_02462_ ) );
OAI211_X1 _10088_ ( .A(_02453_ ), .B(_02462_ ), .C1(_02102_ ), .C2(_02112_ ), .ZN(_02463_ ) );
NAND2_X2 _10089_ ( .A1(_02444_ ), .A2(_02463_ ), .ZN(_02464_ ) );
INV_X1 _10090_ ( .A(\ID_EX_imm [1] ), .ZN(_02465_ ) );
XNOR2_X1 _10091_ ( .A(_02464_ ), .B(_02465_ ), .ZN(_02466_ ) );
NOR2_X1 _10092_ ( .A1(_02102_ ), .A2(_02112_ ), .ZN(_02467_ ) );
NAND2_X1 _10093_ ( .A1(_02467_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_02468_ ) );
OR2_X1 _10094_ ( .A1(_02121_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02469_ ) );
OAI211_X1 _10095_ ( .A(_02469_ ), .B(fanout_net_24 ), .C1(fanout_net_18 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02470_ ) );
OR2_X1 _10096_ ( .A1(fanout_net_18 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02471_ ) );
OAI211_X1 _10097_ ( .A(_02471_ ), .B(_02127_ ), .C1(_02169_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02472_ ) );
NAND3_X1 _10098_ ( .A1(_02470_ ), .A2(_02135_ ), .A3(_02472_ ), .ZN(_02473_ ) );
MUX2_X1 _10099_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02474_ ) );
MUX2_X1 _10100_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02475_ ) );
MUX2_X1 _10101_ ( .A(_02474_ ), .B(_02475_ ), .S(_02127_ ), .Z(_02476_ ) );
OAI211_X1 _10102_ ( .A(fanout_net_27 ), .B(_02473_ ), .C1(_02476_ ), .C2(_02327_ ), .ZN(_02477_ ) );
OR2_X1 _10103_ ( .A1(_02121_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02478_ ) );
OAI211_X1 _10104_ ( .A(_02478_ ), .B(_02127_ ), .C1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C2(fanout_net_18 ), .ZN(_02479_ ) );
OR2_X1 _10105_ ( .A1(fanout_net_18 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02480_ ) );
OAI211_X1 _10106_ ( .A(_02480_ ), .B(fanout_net_24 ), .C1(_02169_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02481_ ) );
NAND3_X1 _10107_ ( .A1(_02479_ ), .A2(_02135_ ), .A3(_02481_ ), .ZN(_02482_ ) );
MUX2_X1 _10108_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02483_ ) );
MUX2_X1 _10109_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02484_ ) );
MUX2_X1 _10110_ ( .A(_02483_ ), .B(_02484_ ), .S(_02127_ ), .Z(_02485_ ) );
OAI211_X1 _10111_ ( .A(_02117_ ), .B(_02482_ ), .C1(_02485_ ), .C2(_02135_ ), .ZN(_02486_ ) );
NAND2_X1 _10112_ ( .A1(_02477_ ), .A2(_02486_ ), .ZN(_02487_ ) );
OAI21_X1 _10113_ ( .A(_02487_ ), .B1(_02102_ ), .B2(_02113_ ), .ZN(_02488_ ) );
AND3_X1 _10114_ ( .A1(_02468_ ), .A2(\ID_EX_imm [0] ), .A3(_02488_ ), .ZN(_02489_ ) );
AND2_X1 _10115_ ( .A1(_02466_ ), .A2(_02489_ ), .ZN(_02490_ ) );
AOI21_X1 _10116_ ( .A(_02465_ ), .B1(_02444_ ), .B2(_02463_ ), .ZN(_02491_ ) );
OAI21_X1 _10117_ ( .A(_02443_ ), .B1(_02490_ ), .B2(_02491_ ), .ZN(_02492_ ) );
INV_X1 _10118_ ( .A(_02441_ ), .ZN(_02493_ ) );
OAI21_X1 _10119_ ( .A(_02492_ ), .B1(_02442_ ), .B2(_02493_ ), .ZN(_02494_ ) );
OR3_X1 _10120_ ( .A1(_02160_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02163_ ), .ZN(_02495_ ) );
OR2_X1 _10121_ ( .A1(_02350_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02496_ ) );
OAI211_X1 _10122_ ( .A(_02496_ ), .B(_02143_ ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02497_ ) );
INV_X1 _10123_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02498_ ) );
NAND2_X1 _10124_ ( .A1(_02498_ ), .A2(fanout_net_18 ), .ZN(_02499_ ) );
OAI211_X1 _10125_ ( .A(_02499_ ), .B(fanout_net_24 ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02500_ ) );
NAND3_X1 _10126_ ( .A1(_02497_ ), .A2(_02500_ ), .A3(_02328_ ), .ZN(_02501_ ) );
MUX2_X1 _10127_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02502_ ) );
MUX2_X1 _10128_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02503_ ) );
MUX2_X1 _10129_ ( .A(_02502_ ), .B(_02503_ ), .S(_02174_ ), .Z(_02504_ ) );
OAI211_X1 _10130_ ( .A(_02119_ ), .B(_02501_ ), .C1(_02504_ ), .C2(_02146_ ), .ZN(_02505_ ) );
OR2_X1 _10131_ ( .A1(_02123_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02506_ ) );
OAI211_X1 _10132_ ( .A(_02506_ ), .B(_02143_ ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02507_ ) );
OR2_X1 _10133_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02508_ ) );
OAI211_X1 _10134_ ( .A(_02508_ ), .B(fanout_net_24 ), .C1(_02152_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02509_ ) );
NAND3_X1 _10135_ ( .A1(_02507_ ), .A2(fanout_net_26 ), .A3(_02509_ ), .ZN(_02510_ ) );
MUX2_X1 _10136_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02511_ ) );
MUX2_X1 _10137_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02512_ ) );
MUX2_X1 _10138_ ( .A(_02511_ ), .B(_02512_ ), .S(fanout_net_24 ), .Z(_02513_ ) );
OAI211_X1 _10139_ ( .A(fanout_net_27 ), .B(_02510_ ), .C1(_02513_ ), .C2(fanout_net_26 ), .ZN(_02514_ ) );
OAI211_X1 _10140_ ( .A(_02505_ ), .B(_02514_ ), .C1(_02104_ ), .C2(_02164_ ), .ZN(_02515_ ) );
NAND2_X1 _10141_ ( .A1(_02495_ ), .A2(_02515_ ), .ZN(_02516_ ) );
XNOR2_X1 _10142_ ( .A(_02516_ ), .B(\ID_EX_imm [3] ), .ZN(_02517_ ) );
INV_X1 _10143_ ( .A(_02517_ ), .ZN(_02518_ ) );
NAND2_X1 _10144_ ( .A1(_02494_ ), .A2(_02518_ ), .ZN(_02519_ ) );
INV_X1 _10145_ ( .A(_02516_ ), .ZN(_02520_ ) );
OR2_X1 _10146_ ( .A1(_02520_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_02521_ ) );
AND2_X1 _10147_ ( .A1(_02519_ ), .A2(_02521_ ), .ZN(_02522_ ) );
OR3_X1 _10148_ ( .A1(_02103_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02112_ ), .ZN(_02523_ ) );
OR2_X1 _10149_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02524_ ) );
OAI211_X1 _10150_ ( .A(_02524_ ), .B(_02142_ ), .C1(_02123_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02525_ ) );
OR2_X1 _10151_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02526_ ) );
OAI211_X1 _10152_ ( .A(_02526_ ), .B(fanout_net_24 ), .C1(_02123_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02527_ ) );
NAND3_X1 _10153_ ( .A1(_02525_ ), .A2(_02527_ ), .A3(_02327_ ), .ZN(_02528_ ) );
MUX2_X1 _10154_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02529_ ) );
MUX2_X1 _10155_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02530_ ) );
MUX2_X1 _10156_ ( .A(_02529_ ), .B(_02530_ ), .S(_02173_ ), .Z(_02531_ ) );
OAI211_X1 _10157_ ( .A(_02118_ ), .B(_02528_ ), .C1(_02531_ ), .C2(_02136_ ), .ZN(_02532_ ) );
OR2_X1 _10158_ ( .A1(_02169_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02533_ ) );
OAI211_X1 _10159_ ( .A(_02533_ ), .B(_02142_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02534_ ) );
OR2_X1 _10160_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02535_ ) );
OAI211_X1 _10161_ ( .A(_02535_ ), .B(fanout_net_24 ), .C1(_02226_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02536_ ) );
NAND3_X1 _10162_ ( .A1(_02534_ ), .A2(fanout_net_26 ), .A3(_02536_ ), .ZN(_02537_ ) );
MUX2_X1 _10163_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02538_ ) );
MUX2_X1 _10164_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02539_ ) );
MUX2_X1 _10165_ ( .A(_02538_ ), .B(_02539_ ), .S(fanout_net_24 ), .Z(_02540_ ) );
OAI211_X1 _10166_ ( .A(fanout_net_27 ), .B(_02537_ ), .C1(_02540_ ), .C2(fanout_net_26 ), .ZN(_02541_ ) );
OAI211_X1 _10167_ ( .A(_02532_ ), .B(_02541_ ), .C1(_02103_ ), .C2(_02113_ ), .ZN(_02542_ ) );
NAND2_X2 _10168_ ( .A1(_02523_ ), .A2(_02542_ ), .ZN(_02543_ ) );
XNOR2_X1 _10169_ ( .A(_02543_ ), .B(\ID_EX_imm [7] ), .ZN(_02544_ ) );
OR3_X1 _10170_ ( .A1(_02102_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02112_ ), .ZN(_02545_ ) );
OR2_X1 _10171_ ( .A1(fanout_net_19 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02546_ ) );
OAI211_X1 _10172_ ( .A(_02546_ ), .B(_02173_ ), .C1(_02226_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02547_ ) );
OR2_X1 _10173_ ( .A1(fanout_net_19 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02548_ ) );
OAI211_X1 _10174_ ( .A(_02548_ ), .B(fanout_net_24 ), .C1(_02226_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02549_ ) );
NAND3_X1 _10175_ ( .A1(_02547_ ), .A2(_02549_ ), .A3(_02327_ ), .ZN(_02550_ ) );
MUX2_X1 _10176_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02551_ ) );
MUX2_X1 _10177_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02552_ ) );
MUX2_X1 _10178_ ( .A(_02551_ ), .B(_02552_ ), .S(_02173_ ), .Z(_02553_ ) );
OAI211_X1 _10179_ ( .A(_02118_ ), .B(_02550_ ), .C1(_02553_ ), .C2(_02136_ ), .ZN(_02554_ ) );
OR2_X1 _10180_ ( .A1(_02122_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02555_ ) );
OAI211_X1 _10181_ ( .A(_02555_ ), .B(fanout_net_24 ), .C1(fanout_net_19 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02556_ ) );
OR2_X1 _10182_ ( .A1(_02122_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02557_ ) );
OAI211_X1 _10183_ ( .A(_02557_ ), .B(_02173_ ), .C1(fanout_net_19 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02558_ ) );
NAND3_X1 _10184_ ( .A1(_02556_ ), .A2(_02558_ ), .A3(fanout_net_26 ), .ZN(_02559_ ) );
MUX2_X1 _10185_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02560_ ) );
MUX2_X1 _10186_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02561_ ) );
MUX2_X1 _10187_ ( .A(_02560_ ), .B(_02561_ ), .S(fanout_net_24 ), .Z(_02562_ ) );
OAI211_X1 _10188_ ( .A(fanout_net_27 ), .B(_02559_ ), .C1(_02562_ ), .C2(fanout_net_26 ), .ZN(_02563_ ) );
OAI211_X1 _10189_ ( .A(_02554_ ), .B(_02563_ ), .C1(_02103_ ), .C2(_02113_ ), .ZN(_02564_ ) );
NAND2_X2 _10190_ ( .A1(_02545_ ), .A2(_02564_ ), .ZN(_02565_ ) );
XOR2_X1 _10191_ ( .A(_02565_ ), .B(\ID_EX_imm [6] ), .Z(_02566_ ) );
INV_X1 _10192_ ( .A(_02566_ ), .ZN(_02567_ ) );
OR3_X1 _10193_ ( .A1(_02102_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02112_ ), .ZN(_02568_ ) );
OR2_X1 _10194_ ( .A1(_02122_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02569_ ) );
OAI211_X1 _10195_ ( .A(_02569_ ), .B(_02173_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02570_ ) );
INV_X1 _10196_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02571_ ) );
INV_X1 _10197_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02572_ ) );
MUX2_X1 _10198_ ( .A(_02571_ ), .B(_02572_ ), .S(fanout_net_19 ), .Z(_02573_ ) );
OAI211_X1 _10199_ ( .A(_02570_ ), .B(_02327_ ), .C1(_02573_ ), .C2(_02142_ ), .ZN(_02574_ ) );
MUX2_X1 _10200_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02575_ ) );
MUX2_X1 _10201_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02576_ ) );
MUX2_X1 _10202_ ( .A(_02575_ ), .B(_02576_ ), .S(_02173_ ), .Z(_02577_ ) );
OAI211_X1 _10203_ ( .A(_02574_ ), .B(fanout_net_27 ), .C1(_02577_ ), .C2(_02136_ ), .ZN(_02578_ ) );
OR2_X1 _10204_ ( .A1(_02122_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02579_ ) );
OAI211_X1 _10205_ ( .A(_02579_ ), .B(_02173_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02580_ ) );
OR2_X1 _10206_ ( .A1(_02122_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02581_ ) );
OAI211_X1 _10207_ ( .A(_02581_ ), .B(fanout_net_24 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02582_ ) );
NAND3_X1 _10208_ ( .A1(_02580_ ), .A2(_02582_ ), .A3(_02327_ ), .ZN(_02583_ ) );
MUX2_X1 _10209_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02584_ ) );
MUX2_X1 _10210_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02585_ ) );
MUX2_X1 _10211_ ( .A(_02584_ ), .B(_02585_ ), .S(_02127_ ), .Z(_02586_ ) );
OAI211_X1 _10212_ ( .A(_02117_ ), .B(_02583_ ), .C1(_02586_ ), .C2(_02327_ ), .ZN(_02587_ ) );
OAI211_X1 _10213_ ( .A(_02578_ ), .B(_02587_ ), .C1(_02103_ ), .C2(_02113_ ), .ZN(_02588_ ) );
NAND2_X1 _10214_ ( .A1(_02568_ ), .A2(_02588_ ), .ZN(_02589_ ) );
XNOR2_X1 _10215_ ( .A(_02589_ ), .B(\ID_EX_imm [5] ), .ZN(_02590_ ) );
OR3_X1 _10216_ ( .A1(_02160_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02163_ ), .ZN(_02591_ ) );
OR2_X1 _10217_ ( .A1(_02226_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02592_ ) );
OAI211_X1 _10218_ ( .A(_02592_ ), .B(_02128_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02593_ ) );
OR2_X1 _10219_ ( .A1(_02226_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02594_ ) );
OAI211_X1 _10220_ ( .A(_02594_ ), .B(fanout_net_24 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02595_ ) );
NAND3_X1 _10221_ ( .A1(_02593_ ), .A2(_02595_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02596_ ) );
MUX2_X1 _10222_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02597_ ) );
MUX2_X1 _10223_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02598_ ) );
MUX2_X1 _10224_ ( .A(_02597_ ), .B(_02598_ ), .S(_02128_ ), .Z(_02599_ ) );
OAI211_X1 _10225_ ( .A(_02118_ ), .B(_02596_ ), .C1(_02599_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02600_ ) );
NOR2_X1 _10226_ ( .A1(_02170_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02601_ ) );
OAI21_X1 _10227_ ( .A(fanout_net_24 ), .B1(fanout_net_20 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02602_ ) );
NOR2_X1 _10228_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02603_ ) );
OAI21_X1 _10229_ ( .A(_02128_ ), .B1(_02170_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02604_ ) );
OAI221_X1 _10230_ ( .A(_02136_ ), .B1(_02601_ ), .B2(_02602_ ), .C1(_02603_ ), .C2(_02604_ ), .ZN(_02605_ ) );
MUX2_X1 _10231_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02606_ ) );
MUX2_X1 _10232_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02607_ ) );
MUX2_X1 _10233_ ( .A(_02606_ ), .B(_02607_ ), .S(fanout_net_24 ), .Z(_02608_ ) );
OAI211_X1 _10234_ ( .A(fanout_net_27 ), .B(_02605_ ), .C1(_02608_ ), .C2(_02328_ ), .ZN(_02609_ ) );
OAI211_X4 _10235_ ( .A(_02600_ ), .B(_02609_ ), .C1(_02160_ ), .C2(_02114_ ), .ZN(_02610_ ) );
NAND2_X4 _10236_ ( .A1(_02591_ ), .A2(_02610_ ), .ZN(_02611_ ) );
INV_X1 _10237_ ( .A(\ID_EX_imm [4] ), .ZN(_02612_ ) );
XNOR2_X2 _10238_ ( .A(_02611_ ), .B(_02612_ ), .ZN(_02613_ ) );
INV_X1 _10239_ ( .A(_02613_ ), .ZN(_02614_ ) );
OR4_X1 _10240_ ( .A1(_02544_ ), .A2(_02567_ ), .A3(_02590_ ), .A4(_02614_ ), .ZN(_02615_ ) );
OR2_X2 _10241_ ( .A1(_02522_ ), .A2(_02615_ ), .ZN(_02616_ ) );
NAND2_X1 _10242_ ( .A1(_02565_ ), .A2(\ID_EX_imm [6] ), .ZN(_02617_ ) );
NOR2_X1 _10243_ ( .A1(_02544_ ), .A2(_02617_ ), .ZN(_02618_ ) );
AOI21_X1 _10244_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02568_ ), .B2(_02588_ ), .ZN(_02619_ ) );
INV_X1 _10245_ ( .A(_02590_ ), .ZN(_02620_ ) );
AOI21_X1 _10246_ ( .A(_02612_ ), .B1(_02591_ ), .B2(_02610_ ), .ZN(_02621_ ) );
AOI21_X1 _10247_ ( .A(_02619_ ), .B1(_02620_ ), .B2(_02621_ ), .ZN(_02622_ ) );
NOR3_X1 _10248_ ( .A1(_02622_ ), .A2(_02544_ ), .A3(_02567_ ), .ZN(_02623_ ) );
AOI211_X1 _10249_ ( .A(_02618_ ), .B(_02623_ ), .C1(\ID_EX_imm [7] ), .C2(_02543_ ), .ZN(_02624_ ) );
AND2_X2 _10250_ ( .A1(_02616_ ), .A2(_02624_ ), .ZN(_02625_ ) );
INV_X1 _10251_ ( .A(_02625_ ), .ZN(_02626_ ) );
OR3_X1 _10252_ ( .A1(_02104_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02163_ ), .ZN(_02627_ ) );
OR2_X1 _10253_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02628_ ) );
OAI211_X1 _10254_ ( .A(_02628_ ), .B(_02143_ ), .C1(_02152_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02629_ ) );
OR2_X1 _10255_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02630_ ) );
OAI211_X1 _10256_ ( .A(_02630_ ), .B(fanout_net_24 ), .C1(_02152_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02631_ ) );
NAND3_X1 _10257_ ( .A1(_02629_ ), .A2(_02631_ ), .A3(_02328_ ), .ZN(_02632_ ) );
MUX2_X1 _10258_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02633_ ) );
MUX2_X1 _10259_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02634_ ) );
MUX2_X1 _10260_ ( .A(_02633_ ), .B(_02634_ ), .S(_02174_ ), .Z(_02635_ ) );
OAI211_X1 _10261_ ( .A(_02119_ ), .B(_02632_ ), .C1(_02635_ ), .C2(_02146_ ), .ZN(_02636_ ) );
OR2_X1 _10262_ ( .A1(_02350_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02637_ ) );
OAI211_X1 _10263_ ( .A(_02637_ ), .B(_02143_ ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02638_ ) );
OR2_X1 _10264_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02639_ ) );
OAI211_X1 _10265_ ( .A(_02639_ ), .B(fanout_net_24 ), .C1(_02152_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02640_ ) );
NAND3_X1 _10266_ ( .A1(_02638_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02640_ ), .ZN(_02641_ ) );
MUX2_X1 _10267_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02642_ ) );
MUX2_X1 _10268_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02643_ ) );
MUX2_X1 _10269_ ( .A(_02642_ ), .B(_02643_ ), .S(fanout_net_24 ), .Z(_02644_ ) );
OAI211_X1 _10270_ ( .A(fanout_net_27 ), .B(_02641_ ), .C1(_02644_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02645_ ) );
OAI211_X1 _10271_ ( .A(_02636_ ), .B(_02645_ ), .C1(_02161_ ), .C2(_02164_ ), .ZN(_02646_ ) );
NAND2_X2 _10272_ ( .A1(_02627_ ), .A2(_02646_ ), .ZN(_02647_ ) );
INV_X1 _10273_ ( .A(\ID_EX_imm [12] ), .ZN(_02648_ ) );
XNOR2_X1 _10274_ ( .A(_02647_ ), .B(_02648_ ), .ZN(_02649_ ) );
OR2_X1 _10275_ ( .A1(_02226_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02650_ ) );
OAI211_X1 _10276_ ( .A(_02650_ ), .B(_02174_ ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02651_ ) );
OR2_X1 _10277_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02652_ ) );
OAI211_X1 _10278_ ( .A(_02652_ ), .B(fanout_net_24 ), .C1(_02227_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02653_ ) );
NAND3_X1 _10279_ ( .A1(_02651_ ), .A2(_02136_ ), .A3(_02653_ ), .ZN(_02654_ ) );
MUX2_X1 _10280_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02655_ ) );
MUX2_X1 _10281_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02656_ ) );
MUX2_X1 _10282_ ( .A(_02655_ ), .B(_02656_ ), .S(_02128_ ), .Z(_02657_ ) );
OAI211_X1 _10283_ ( .A(fanout_net_27 ), .B(_02654_ ), .C1(_02657_ ), .C2(_02137_ ), .ZN(_02658_ ) );
MUX2_X1 _10284_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02659_ ) );
AND2_X1 _10285_ ( .A1(_02659_ ), .A2(_02128_ ), .ZN(_02660_ ) );
MUX2_X1 _10286_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02661_ ) );
AOI211_X1 _10287_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_02660_ ), .C1(fanout_net_24 ), .C2(_02661_ ), .ZN(_02662_ ) );
MUX2_X1 _10288_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02663_ ) );
MUX2_X1 _10289_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02664_ ) );
MUX2_X1 _10290_ ( .A(_02663_ ), .B(_02664_ ), .S(_02142_ ), .Z(_02665_ ) );
OAI21_X1 _10291_ ( .A(_02118_ ), .B1(_02665_ ), .B2(_02328_ ), .ZN(_02666_ ) );
OAI221_X1 _10292_ ( .A(_02658_ ), .B1(_02662_ ), .B2(_02666_ ), .C1(_02104_ ), .C2(_02114_ ), .ZN(_02667_ ) );
OR3_X1 _10293_ ( .A1(_02160_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02163_ ), .ZN(_02668_ ) );
INV_X1 _10294_ ( .A(\ID_EX_imm [13] ), .ZN(_02669_ ) );
AND3_X1 _10295_ ( .A1(_02667_ ), .A2(_02668_ ), .A3(_02669_ ), .ZN(_02670_ ) );
AOI21_X1 _10296_ ( .A(_02669_ ), .B1(_02667_ ), .B2(_02668_ ), .ZN(_02671_ ) );
NOR2_X1 _10297_ ( .A1(_02670_ ), .A2(_02671_ ), .ZN(_02672_ ) );
AND2_X1 _10298_ ( .A1(_02649_ ), .A2(_02672_ ), .ZN(_02673_ ) );
OR3_X1 _10299_ ( .A1(_02104_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02114_ ), .ZN(_02674_ ) );
OR2_X1 _10300_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02675_ ) );
OAI211_X1 _10301_ ( .A(_02675_ ), .B(_02129_ ), .C1(_02124_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02676_ ) );
OR2_X1 _10302_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02677_ ) );
OAI211_X1 _10303_ ( .A(_02677_ ), .B(fanout_net_24 ), .C1(_02124_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02678_ ) );
NAND3_X1 _10304_ ( .A1(_02676_ ), .A2(_02678_ ), .A3(_02137_ ), .ZN(_02679_ ) );
MUX2_X1 _10305_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02680_ ) );
MUX2_X1 _10306_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02681_ ) );
MUX2_X1 _10307_ ( .A(_02680_ ), .B(_02681_ ), .S(_02143_ ), .Z(_02682_ ) );
OAI211_X1 _10308_ ( .A(_02119_ ), .B(_02679_ ), .C1(_02682_ ), .C2(_02146_ ), .ZN(_02683_ ) );
OR2_X1 _10309_ ( .A1(_02350_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02684_ ) );
OAI211_X1 _10310_ ( .A(_02684_ ), .B(fanout_net_24 ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02685_ ) );
OR2_X1 _10311_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02686_ ) );
OAI211_X1 _10312_ ( .A(_02686_ ), .B(_02129_ ), .C1(_02124_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02687_ ) );
NAND3_X1 _10313_ ( .A1(_02685_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02687_ ), .ZN(_02688_ ) );
MUX2_X1 _10314_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02689_ ) );
MUX2_X1 _10315_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02690_ ) );
MUX2_X1 _10316_ ( .A(_02689_ ), .B(_02690_ ), .S(fanout_net_24 ), .Z(_02691_ ) );
OAI211_X1 _10317_ ( .A(fanout_net_27 ), .B(_02688_ ), .C1(_02691_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02692_ ) );
OAI211_X1 _10318_ ( .A(_02683_ ), .B(_02692_ ), .C1(_02161_ ), .C2(_02164_ ), .ZN(_02693_ ) );
NAND2_X2 _10319_ ( .A1(_02674_ ), .A2(_02693_ ), .ZN(_02694_ ) );
INV_X1 _10320_ ( .A(\ID_EX_imm [15] ), .ZN(_02695_ ) );
XNOR2_X1 _10321_ ( .A(_02694_ ), .B(_02695_ ), .ZN(_02696_ ) );
OR3_X1 _10322_ ( .A1(_02161_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02114_ ), .ZN(_02697_ ) );
OR2_X1 _10323_ ( .A1(_02170_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02698_ ) );
OAI211_X1 _10324_ ( .A(_02698_ ), .B(_02175_ ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02699_ ) );
OR2_X1 _10325_ ( .A1(_02170_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02700_ ) );
OAI211_X1 _10326_ ( .A(_02700_ ), .B(fanout_net_25 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02701_ ) );
NAND3_X1 _10327_ ( .A1(_02699_ ), .A2(_02701_ ), .A3(_02137_ ), .ZN(_02702_ ) );
MUX2_X1 _10328_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02703_ ) );
MUX2_X1 _10329_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02704_ ) );
MUX2_X1 _10330_ ( .A(_02703_ ), .B(_02704_ ), .S(_02129_ ), .Z(_02705_ ) );
OAI211_X1 _10331_ ( .A(_02119_ ), .B(_02702_ ), .C1(_02705_ ), .C2(_02146_ ), .ZN(_02706_ ) );
OR2_X1 _10332_ ( .A1(_02170_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02707_ ) );
OAI211_X1 _10333_ ( .A(_02707_ ), .B(_02175_ ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02708_ ) );
OR2_X1 _10334_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02709_ ) );
OAI211_X1 _10335_ ( .A(_02709_ ), .B(fanout_net_25 ), .C1(_02124_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02710_ ) );
NAND3_X1 _10336_ ( .A1(_02708_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02710_ ), .ZN(_02711_ ) );
MUX2_X1 _10337_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02712_ ) );
MUX2_X1 _10338_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02713_ ) );
MUX2_X1 _10339_ ( .A(_02712_ ), .B(_02713_ ), .S(fanout_net_25 ), .Z(_02714_ ) );
OAI211_X1 _10340_ ( .A(fanout_net_27 ), .B(_02711_ ), .C1(_02714_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02715_ ) );
OAI211_X1 _10341_ ( .A(_02706_ ), .B(_02715_ ), .C1(_02161_ ), .C2(_02164_ ), .ZN(_02716_ ) );
NAND2_X1 _10342_ ( .A1(_02697_ ), .A2(_02716_ ), .ZN(_02717_ ) );
BUF_X4 _10343_ ( .A(_02717_ ), .Z(_02718_ ) );
XOR2_X1 _10344_ ( .A(_02718_ ), .B(\ID_EX_imm [14] ), .Z(_02719_ ) );
AND3_X1 _10345_ ( .A1(_02673_ ), .A2(_02696_ ), .A3(_02719_ ), .ZN(_02720_ ) );
OR3_X1 _10346_ ( .A1(_02103_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02113_ ), .ZN(_02721_ ) );
OR2_X1 _10347_ ( .A1(_02169_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02722_ ) );
OAI211_X1 _10348_ ( .A(_02722_ ), .B(fanout_net_25 ), .C1(fanout_net_21 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02723_ ) );
OR2_X1 _10349_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02724_ ) );
OAI211_X1 _10350_ ( .A(_02724_ ), .B(_02142_ ), .C1(_02123_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02725_ ) );
NAND3_X1 _10351_ ( .A1(_02723_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02725_ ), .ZN(_02726_ ) );
MUX2_X1 _10352_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02727_ ) );
MUX2_X1 _10353_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02728_ ) );
MUX2_X1 _10354_ ( .A(_02727_ ), .B(_02728_ ), .S(_02142_ ), .Z(_02729_ ) );
OAI211_X1 _10355_ ( .A(_02118_ ), .B(_02726_ ), .C1(_02729_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02730_ ) );
NOR2_X1 _10356_ ( .A1(_02226_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02731_ ) );
OAI21_X1 _10357_ ( .A(fanout_net_25 ), .B1(fanout_net_21 ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02732_ ) );
NOR2_X1 _10358_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02733_ ) );
OAI21_X1 _10359_ ( .A(_02173_ ), .B1(_02226_ ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02734_ ) );
OAI221_X1 _10360_ ( .A(_02327_ ), .B1(_02731_ ), .B2(_02732_ ), .C1(_02733_ ), .C2(_02734_ ), .ZN(_02735_ ) );
MUX2_X1 _10361_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02736_ ) );
MUX2_X1 _10362_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02737_ ) );
MUX2_X1 _10363_ ( .A(_02736_ ), .B(_02737_ ), .S(fanout_net_25 ), .Z(_02738_ ) );
OAI211_X1 _10364_ ( .A(fanout_net_27 ), .B(_02735_ ), .C1(_02738_ ), .C2(_02136_ ), .ZN(_02739_ ) );
OAI211_X1 _10365_ ( .A(_02730_ ), .B(_02739_ ), .C1(_02103_ ), .C2(_02113_ ), .ZN(_02740_ ) );
NAND2_X1 _10366_ ( .A1(_02721_ ), .A2(_02740_ ), .ZN(_02741_ ) );
BUF_X4 _10367_ ( .A(_02741_ ), .Z(_02742_ ) );
INV_X1 _10368_ ( .A(\ID_EX_imm [10] ), .ZN(_02743_ ) );
XNOR2_X1 _10369_ ( .A(_02742_ ), .B(_02743_ ), .ZN(_02744_ ) );
OR3_X1 _10370_ ( .A1(_02103_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_02113_ ), .ZN(_02745_ ) );
OR2_X1 _10371_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02746_ ) );
OAI211_X1 _10372_ ( .A(_02746_ ), .B(_02128_ ), .C1(_02170_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02747_ ) );
OR2_X1 _10373_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02748_ ) );
OAI211_X1 _10374_ ( .A(_02748_ ), .B(fanout_net_25 ), .C1(_02350_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02749_ ) );
NAND3_X1 _10375_ ( .A1(_02747_ ), .A2(_02749_ ), .A3(_02136_ ), .ZN(_02750_ ) );
MUX2_X1 _10376_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02751_ ) );
MUX2_X1 _10377_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02752_ ) );
MUX2_X1 _10378_ ( .A(_02751_ ), .B(_02752_ ), .S(_02142_ ), .Z(_02753_ ) );
OAI211_X1 _10379_ ( .A(_02118_ ), .B(_02750_ ), .C1(_02753_ ), .C2(_02328_ ), .ZN(_02754_ ) );
OR2_X1 _10380_ ( .A1(_02169_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02755_ ) );
OAI211_X1 _10381_ ( .A(_02755_ ), .B(_02128_ ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02756_ ) );
OR2_X1 _10382_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02757_ ) );
OAI211_X1 _10383_ ( .A(_02757_ ), .B(fanout_net_25 ), .C1(_02350_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02758_ ) );
NAND3_X1 _10384_ ( .A1(_02756_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02758_ ), .ZN(_02759_ ) );
MUX2_X1 _10385_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02760_ ) );
MUX2_X1 _10386_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02761_ ) );
MUX2_X1 _10387_ ( .A(_02760_ ), .B(_02761_ ), .S(fanout_net_25 ), .Z(_02762_ ) );
OAI211_X1 _10388_ ( .A(fanout_net_27 ), .B(_02759_ ), .C1(_02762_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02763_ ) );
OAI211_X1 _10389_ ( .A(_02754_ ), .B(_02763_ ), .C1(_02160_ ), .C2(_02163_ ), .ZN(_02764_ ) );
NAND2_X2 _10390_ ( .A1(_02745_ ), .A2(_02764_ ), .ZN(_02765_ ) );
INV_X1 _10391_ ( .A(\ID_EX_imm [11] ), .ZN(_02766_ ) );
XNOR2_X1 _10392_ ( .A(_02765_ ), .B(_02766_ ), .ZN(_02767_ ) );
AND2_X1 _10393_ ( .A1(_02744_ ), .A2(_02767_ ), .ZN(_02768_ ) );
OR3_X1 _10394_ ( .A1(_02160_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02163_ ), .ZN(_02769_ ) );
OR2_X1 _10395_ ( .A1(_02123_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02770_ ) );
OAI211_X1 _10396_ ( .A(_02770_ ), .B(_02174_ ), .C1(fanout_net_21 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02771_ ) );
OR2_X1 _10397_ ( .A1(fanout_net_21 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02772_ ) );
OAI211_X1 _10398_ ( .A(_02772_ ), .B(fanout_net_25 ), .C1(_02227_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02773_ ) );
NAND3_X1 _10399_ ( .A1(_02771_ ), .A2(_02328_ ), .A3(_02773_ ), .ZN(_02774_ ) );
MUX2_X1 _10400_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02775_ ) );
MUX2_X1 _10401_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02776_ ) );
MUX2_X1 _10402_ ( .A(_02775_ ), .B(_02776_ ), .S(_02128_ ), .Z(_02777_ ) );
OAI211_X1 _10403_ ( .A(_02118_ ), .B(_02774_ ), .C1(_02777_ ), .C2(_02137_ ), .ZN(_02778_ ) );
OR2_X1 _10404_ ( .A1(fanout_net_21 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02779_ ) );
OAI211_X1 _10405_ ( .A(_02779_ ), .B(fanout_net_25 ), .C1(_02227_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02780_ ) );
OR2_X1 _10406_ ( .A1(fanout_net_21 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02781_ ) );
OAI211_X1 _10407_ ( .A(_02781_ ), .B(_02174_ ), .C1(_02227_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02782_ ) );
NAND3_X1 _10408_ ( .A1(_02780_ ), .A2(_02782_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02783_ ) );
MUX2_X1 _10409_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02784_ ) );
MUX2_X1 _10410_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02785_ ) );
MUX2_X1 _10411_ ( .A(_02784_ ), .B(_02785_ ), .S(fanout_net_25 ), .Z(_02786_ ) );
OAI211_X1 _10412_ ( .A(fanout_net_27 ), .B(_02783_ ), .C1(_02786_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02787_ ) );
OAI211_X1 _10413_ ( .A(_02778_ ), .B(_02787_ ), .C1(_02104_ ), .C2(_02114_ ), .ZN(_02788_ ) );
NAND2_X2 _10414_ ( .A1(_02769_ ), .A2(_02788_ ), .ZN(_02789_ ) );
INV_X1 _10415_ ( .A(\ID_EX_imm [8] ), .ZN(_02790_ ) );
XNOR2_X1 _10416_ ( .A(_02789_ ), .B(_02790_ ), .ZN(_02791_ ) );
OR3_X1 _10417_ ( .A1(_02103_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02113_ ), .ZN(_02792_ ) );
OR2_X1 _10418_ ( .A1(_02169_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02793_ ) );
OAI211_X1 _10419_ ( .A(_02793_ ), .B(_02128_ ), .C1(fanout_net_22 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02794_ ) );
OR2_X1 _10420_ ( .A1(fanout_net_22 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02795_ ) );
OAI211_X1 _10421_ ( .A(_02795_ ), .B(fanout_net_25 ), .C1(_02350_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02796_ ) );
NAND3_X1 _10422_ ( .A1(_02794_ ), .A2(_02136_ ), .A3(_02796_ ), .ZN(_02797_ ) );
MUX2_X1 _10423_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02798_ ) );
MUX2_X1 _10424_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02799_ ) );
MUX2_X1 _10425_ ( .A(_02798_ ), .B(_02799_ ), .S(_02142_ ), .Z(_02800_ ) );
OAI211_X1 _10426_ ( .A(_02118_ ), .B(_02797_ ), .C1(_02800_ ), .C2(_02328_ ), .ZN(_02801_ ) );
OR2_X1 _10427_ ( .A1(_02169_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02802_ ) );
OAI211_X1 _10428_ ( .A(_02802_ ), .B(fanout_net_25 ), .C1(fanout_net_22 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02803_ ) );
OR2_X1 _10429_ ( .A1(_02169_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02804_ ) );
OAI211_X1 _10430_ ( .A(_02804_ ), .B(_02142_ ), .C1(fanout_net_22 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02805_ ) );
NAND3_X1 _10431_ ( .A1(_02803_ ), .A2(_02805_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02806_ ) );
MUX2_X1 _10432_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02807_ ) );
MUX2_X1 _10433_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02808_ ) );
MUX2_X1 _10434_ ( .A(_02807_ ), .B(_02808_ ), .S(fanout_net_25 ), .Z(_02809_ ) );
OAI211_X1 _10435_ ( .A(fanout_net_27 ), .B(_02806_ ), .C1(_02809_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02810_ ) );
OAI211_X1 _10436_ ( .A(_02801_ ), .B(_02810_ ), .C1(_02160_ ), .C2(_02163_ ), .ZN(_02811_ ) );
NAND2_X2 _10437_ ( .A1(_02792_ ), .A2(_02811_ ), .ZN(_02812_ ) );
INV_X1 _10438_ ( .A(\ID_EX_imm [9] ), .ZN(_02813_ ) );
XNOR2_X1 _10439_ ( .A(_02812_ ), .B(_02813_ ), .ZN(_02814_ ) );
AND2_X1 _10440_ ( .A1(_02791_ ), .A2(_02814_ ), .ZN(_02815_ ) );
AND2_X1 _10441_ ( .A1(_02768_ ), .A2(_02815_ ), .ZN(_02816_ ) );
AND3_X1 _10442_ ( .A1(_02626_ ), .A2(_02720_ ), .A3(_02816_ ), .ZN(_02817_ ) );
INV_X1 _10443_ ( .A(_02817_ ), .ZN(_02818_ ) );
AND2_X1 _10444_ ( .A1(_02789_ ), .A2(\ID_EX_imm [8] ), .ZN(_02819_ ) );
AND2_X1 _10445_ ( .A1(_02814_ ), .A2(_02819_ ), .ZN(_02820_ ) );
AOI21_X1 _10446_ ( .A(_02820_ ), .B1(\ID_EX_imm [9] ), .B2(_02812_ ), .ZN(_02821_ ) );
INV_X1 _10447_ ( .A(_02821_ ), .ZN(_02822_ ) );
AND2_X1 _10448_ ( .A1(_02822_ ), .A2(_02768_ ), .ZN(_02823_ ) );
AOI21_X1 _10449_ ( .A(_02766_ ), .B1(_02745_ ), .B2(_02764_ ), .ZN(_02824_ ) );
AND2_X1 _10450_ ( .A1(_02742_ ), .A2(\ID_EX_imm [10] ), .ZN(_02825_ ) );
AND2_X1 _10451_ ( .A1(_02767_ ), .A2(_02825_ ), .ZN(_02826_ ) );
NOR3_X1 _10452_ ( .A1(_02823_ ), .A2(_02824_ ), .A3(_02826_ ), .ZN(_02827_ ) );
INV_X1 _10453_ ( .A(_02827_ ), .ZN(_02828_ ) );
NAND2_X1 _10454_ ( .A1(_02828_ ), .A2(_02720_ ), .ZN(_02829_ ) );
OAI211_X1 _10455_ ( .A(\ID_EX_imm [14] ), .B(_02718_ ), .C1(_02694_ ), .C2(\ID_EX_imm [15] ), .ZN(_02830_ ) );
NAND2_X1 _10456_ ( .A1(_02647_ ), .A2(\ID_EX_imm [12] ), .ZN(_02831_ ) );
NOR3_X1 _10457_ ( .A1(_02831_ ), .A2(_02670_ ), .A3(_02671_ ), .ZN(_02832_ ) );
OR2_X1 _10458_ ( .A1(_02832_ ), .A2(_02671_ ), .ZN(_02833_ ) );
AND2_X1 _10459_ ( .A1(_02719_ ), .A2(_02696_ ), .ZN(_02834_ ) );
AOI22_X1 _10460_ ( .A1(_02833_ ), .A2(_02834_ ), .B1(\ID_EX_imm [15] ), .B2(_02694_ ), .ZN(_02835_ ) );
AND3_X1 _10461_ ( .A1(_02829_ ), .A2(_02830_ ), .A3(_02835_ ), .ZN(_02836_ ) );
AOI211_X1 _10462_ ( .A(_02323_ ), .B(_02420_ ), .C1(_02818_ ), .C2(_02836_ ), .ZN(_02837_ ) );
INV_X1 _10463_ ( .A(_02837_ ), .ZN(_02838_ ) );
AND2_X1 _10464_ ( .A1(_02417_ ), .A2(\ID_EX_imm [16] ), .ZN(_02839_ ) );
AND2_X1 _10465_ ( .A1(_02396_ ), .A2(_02839_ ), .ZN(_02840_ ) );
AOI21_X1 _10466_ ( .A(_02840_ ), .B1(\ID_EX_imm [17] ), .B2(_02394_ ), .ZN(_02841_ ) );
INV_X1 _10467_ ( .A(_02841_ ), .ZN(_02842_ ) );
AND2_X1 _10468_ ( .A1(_02842_ ), .A2(_02373_ ), .ZN(_02843_ ) );
AOI21_X1 _10469_ ( .A(_02371_ ), .B1(_02349_ ), .B2(_02369_ ), .ZN(_02844_ ) );
AND2_X1 _10470_ ( .A1(_02346_ ), .A2(\ID_EX_imm [18] ), .ZN(_02845_ ) );
AND2_X1 _10471_ ( .A1(_02372_ ), .A2(_02845_ ), .ZN(_02846_ ) );
NOR3_X1 _10472_ ( .A1(_02843_ ), .A2(_02844_ ), .A3(_02846_ ), .ZN(_02847_ ) );
OR2_X1 _10473_ ( .A1(_02847_ ), .A2(_02323_ ), .ZN(_02848_ ) );
OAI211_X1 _10474_ ( .A(\ID_EX_imm [22] ), .B(_02270_ ), .C1(_02247_ ), .C2(\ID_EX_imm [23] ), .ZN(_02849_ ) );
NAND2_X1 _10475_ ( .A1(_02294_ ), .A2(\ID_EX_imm [20] ), .ZN(_02850_ ) );
NOR3_X1 _10476_ ( .A1(_02850_ ), .A2(_02318_ ), .A3(_02319_ ), .ZN(_02851_ ) );
OR2_X1 _10477_ ( .A1(_02851_ ), .A2(_02319_ ), .ZN(_02852_ ) );
AOI22_X1 _10478_ ( .A1(_02852_ ), .A2(_02273_ ), .B1(\ID_EX_imm [23] ), .B2(_02247_ ), .ZN(_02853_ ) );
AND3_X1 _10479_ ( .A1(_02848_ ), .A2(_02849_ ), .A3(_02853_ ), .ZN(_02854_ ) );
NAND2_X2 _10480_ ( .A1(_02838_ ), .A2(_02854_ ), .ZN(_02855_ ) );
OR3_X1 _10481_ ( .A1(_02162_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02165_ ), .ZN(_02856_ ) );
OR2_X1 _10482_ ( .A1(_02153_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02857_ ) );
OAI211_X1 _10483_ ( .A(_02857_ ), .B(fanout_net_25 ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02858_ ) );
OR2_X1 _10484_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02859_ ) );
OAI211_X1 _10485_ ( .A(_02859_ ), .B(_02176_ ), .C1(_02179_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02860_ ) );
NAND3_X1 _10486_ ( .A1(_02858_ ), .A2(_02147_ ), .A3(_02860_ ), .ZN(_02861_ ) );
MUX2_X1 _10487_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02862_ ) );
MUX2_X1 _10488_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02863_ ) );
MUX2_X1 _10489_ ( .A(_02862_ ), .B(_02863_ ), .S(_02176_ ), .Z(_02864_ ) );
OAI211_X1 _10490_ ( .A(_02120_ ), .B(_02861_ ), .C1(_02864_ ), .C2(_02147_ ), .ZN(_02865_ ) );
OR2_X1 _10491_ ( .A1(_02171_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02866_ ) );
OAI211_X1 _10492_ ( .A(_02866_ ), .B(_02176_ ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02867_ ) );
NOR2_X1 _10493_ ( .A1(_02179_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02868_ ) );
OAI21_X1 _10494_ ( .A(fanout_net_25 ), .B1(fanout_net_22 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02869_ ) );
OAI211_X1 _10495_ ( .A(_02867_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .C1(_02868_ ), .C2(_02869_ ), .ZN(_02870_ ) );
MUX2_X1 _10496_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02871_ ) );
MUX2_X1 _10497_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02872_ ) );
MUX2_X1 _10498_ ( .A(_02871_ ), .B(_02872_ ), .S(fanout_net_25 ), .Z(_02873_ ) );
OAI211_X1 _10499_ ( .A(_02870_ ), .B(fanout_net_27 ), .C1(_02873_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02874_ ) );
OAI211_X1 _10500_ ( .A(_02865_ ), .B(_02874_ ), .C1(_02162_ ), .C2(_02165_ ), .ZN(_02875_ ) );
NAND2_X2 _10501_ ( .A1(_02856_ ), .A2(_02875_ ), .ZN(_02876_ ) );
INV_X1 _10502_ ( .A(\ID_EX_imm [24] ), .ZN(_02877_ ) );
XNOR2_X1 _10503_ ( .A(_02876_ ), .B(_02877_ ), .ZN(_02878_ ) );
OR3_X1 _10504_ ( .A1(_02161_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02164_ ), .ZN(_02879_ ) );
OR2_X1 _10505_ ( .A1(_02152_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02880_ ) );
OAI211_X1 _10506_ ( .A(_02880_ ), .B(_02144_ ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02881_ ) );
OR2_X1 _10507_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02882_ ) );
OAI211_X1 _10508_ ( .A(_02882_ ), .B(fanout_net_25 ), .C1(_02153_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02883_ ) );
NAND3_X1 _10509_ ( .A1(_02881_ ), .A2(_02883_ ), .A3(_02146_ ), .ZN(_02884_ ) );
MUX2_X1 _10510_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02885_ ) );
MUX2_X1 _10511_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02886_ ) );
MUX2_X1 _10512_ ( .A(_02885_ ), .B(_02886_ ), .S(_02175_ ), .Z(_02887_ ) );
OAI211_X1 _10513_ ( .A(_02120_ ), .B(_02884_ ), .C1(_02887_ ), .C2(_02138_ ), .ZN(_02888_ ) );
OR2_X1 _10514_ ( .A1(_02227_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02889_ ) );
OAI211_X1 _10515_ ( .A(_02889_ ), .B(_02175_ ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02890_ ) );
NOR2_X1 _10516_ ( .A1(_02153_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02891_ ) );
OAI21_X1 _10517_ ( .A(fanout_net_25 ), .B1(fanout_net_22 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02892_ ) );
OAI211_X1 _10518_ ( .A(_02890_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .C1(_02891_ ), .C2(_02892_ ), .ZN(_02893_ ) );
MUX2_X1 _10519_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02894_ ) );
MUX2_X1 _10520_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02895_ ) );
MUX2_X1 _10521_ ( .A(_02894_ ), .B(_02895_ ), .S(fanout_net_25 ), .Z(_02896_ ) );
OAI211_X1 _10522_ ( .A(_02893_ ), .B(fanout_net_27 ), .C1(_02896_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02897_ ) );
OAI211_X1 _10523_ ( .A(_02888_ ), .B(_02897_ ), .C1(_02105_ ), .C2(_02115_ ), .ZN(_02898_ ) );
NAND2_X2 _10524_ ( .A1(_02879_ ), .A2(_02898_ ), .ZN(_02899_ ) );
INV_X1 _10525_ ( .A(\ID_EX_imm [25] ), .ZN(_02900_ ) );
XNOR2_X1 _10526_ ( .A(_02899_ ), .B(_02900_ ), .ZN(_02901_ ) );
AND3_X2 _10527_ ( .A1(_02855_ ), .A2(_02878_ ), .A3(_02901_ ), .ZN(_02902_ ) );
AND2_X1 _10528_ ( .A1(_02899_ ), .A2(\ID_EX_imm [25] ), .ZN(_02903_ ) );
AND3_X1 _10529_ ( .A1(_02879_ ), .A2(_02900_ ), .A3(_02898_ ), .ZN(_02904_ ) );
NAND2_X1 _10530_ ( .A1(_02876_ ), .A2(\ID_EX_imm [24] ), .ZN(_02905_ ) );
OR3_X1 _10531_ ( .A1(_02903_ ), .A2(_02904_ ), .A3(_02905_ ), .ZN(_02906_ ) );
INV_X1 _10532_ ( .A(_02899_ ), .ZN(_02907_ ) );
OAI21_X1 _10533_ ( .A(_02906_ ), .B1(_02900_ ), .B2(_02907_ ), .ZN(_02908_ ) );
OAI21_X2 _10534_ ( .A(_02224_ ), .B1(_02902_ ), .B2(_02908_ ), .ZN(_02909_ ) );
NAND2_X1 _10535_ ( .A1(_02196_ ), .A2(\ID_EX_imm [26] ), .ZN(_02910_ ) );
NOR3_X1 _10536_ ( .A1(_02910_ ), .A2(_02221_ ), .A3(_02222_ ), .ZN(_02911_ ) );
NOR2_X1 _10537_ ( .A1(_02911_ ), .A2(_02222_ ), .ZN(_02912_ ) );
AOI21_X2 _10538_ ( .A(_02168_ ), .B1(_02909_ ), .B2(_02912_ ), .ZN(_02913_ ) );
OR3_X1 _10539_ ( .A1(_02104_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02114_ ), .ZN(_02914_ ) );
OR2_X1 _10540_ ( .A1(_02170_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02915_ ) );
OAI211_X1 _10541_ ( .A(_02915_ ), .B(fanout_net_25 ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02916_ ) );
OR2_X1 _10542_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02917_ ) );
OAI211_X1 _10543_ ( .A(_02917_ ), .B(_02129_ ), .C1(_02124_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02918_ ) );
NAND3_X1 _10544_ ( .A1(_02916_ ), .A2(_02137_ ), .A3(_02918_ ), .ZN(_02919_ ) );
MUX2_X1 _10545_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02920_ ) );
MUX2_X1 _10546_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02921_ ) );
MUX2_X1 _10547_ ( .A(_02920_ ), .B(_02921_ ), .S(_02143_ ), .Z(_02922_ ) );
OAI211_X1 _10548_ ( .A(_02119_ ), .B(_02919_ ), .C1(_02922_ ), .C2(_02146_ ), .ZN(_02923_ ) );
OR2_X1 _10549_ ( .A1(_02170_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02924_ ) );
OAI211_X1 _10550_ ( .A(_02924_ ), .B(fanout_net_25 ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02925_ ) );
OR2_X1 _10551_ ( .A1(_02170_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02926_ ) );
OAI211_X1 _10552_ ( .A(_02926_ ), .B(_02129_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02927_ ) );
NAND3_X1 _10553_ ( .A1(_02925_ ), .A2(_02927_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02928_ ) );
MUX2_X1 _10554_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02929_ ) );
MUX2_X1 _10555_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02930_ ) );
MUX2_X1 _10556_ ( .A(_02929_ ), .B(_02930_ ), .S(fanout_net_25 ), .Z(_02931_ ) );
OAI211_X1 _10557_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02928_ ), .C1(_02931_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02932_ ) );
OAI211_X1 _10558_ ( .A(_02923_ ), .B(_02932_ ), .C1(_02161_ ), .C2(_02164_ ), .ZN(_02933_ ) );
NAND2_X1 _10559_ ( .A1(_02914_ ), .A2(_02933_ ), .ZN(_02934_ ) );
INV_X1 _10560_ ( .A(\ID_EX_imm [29] ), .ZN(_02935_ ) );
XNOR2_X1 _10561_ ( .A(_02934_ ), .B(_02935_ ), .ZN(_02936_ ) );
AND2_X1 _10562_ ( .A1(_02913_ ), .A2(_02936_ ), .ZN(_02937_ ) );
AOI21_X1 _10563_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02116_ ), .B2(_02166_ ), .ZN(_02938_ ) );
NAND2_X1 _10564_ ( .A1(_02936_ ), .A2(_02938_ ), .ZN(_02939_ ) );
INV_X1 _10565_ ( .A(_02934_ ), .ZN(_02940_ ) );
OAI21_X1 _10566_ ( .A(_02939_ ), .B1(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_02940_ ), .ZN(_02941_ ) );
NOR2_X1 _10567_ ( .A1(_02937_ ), .A2(_02941_ ), .ZN(_02942_ ) );
MUX2_X1 _10568_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02943_ ) );
AND2_X1 _10569_ ( .A1(_02943_ ), .A2(_02175_ ), .ZN(_02944_ ) );
MUX2_X1 _10570_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02945_ ) );
AOI211_X1 _10571_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_02944_ ), .C1(fanout_net_25 ), .C2(_02945_ ), .ZN(_02946_ ) );
MUX2_X1 _10572_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02947_ ) );
AND2_X1 _10573_ ( .A1(_02947_ ), .A2(_02129_ ), .ZN(_02948_ ) );
MUX2_X1 _10574_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02949_ ) );
AOI211_X1 _10575_ ( .A(_02137_ ), .B(_02948_ ), .C1(fanout_net_25 ), .C2(_02949_ ), .ZN(_02950_ ) );
OR3_X1 _10576_ ( .A1(_02946_ ), .A2(_02950_ ), .A3(_02119_ ), .ZN(_02951_ ) );
MUX2_X1 _10577_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02952_ ) );
AND2_X1 _10578_ ( .A1(_02952_ ), .A2(_02175_ ), .ZN(_02953_ ) );
MUX2_X1 _10579_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02954_ ) );
AOI211_X1 _10580_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_02953_ ), .C1(fanout_net_25 ), .C2(_02954_ ), .ZN(_02955_ ) );
MUX2_X1 _10581_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02956_ ) );
AND2_X1 _10582_ ( .A1(_02956_ ), .A2(_02129_ ), .ZN(_02957_ ) );
MUX2_X1 _10583_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02958_ ) );
AOI211_X1 _10584_ ( .A(_02137_ ), .B(_02957_ ), .C1(fanout_net_25 ), .C2(_02958_ ), .ZN(_02959_ ) );
OR3_X1 _10585_ ( .A1(_02955_ ), .A2(_02959_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .ZN(_02960_ ) );
OAI211_X1 _10586_ ( .A(_02951_ ), .B(_02960_ ), .C1(_02165_ ), .C2(_02162_ ), .ZN(_02961_ ) );
OR3_X4 _10587_ ( .A1(_02105_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02115_ ), .ZN(_02962_ ) );
AND2_X2 _10588_ ( .A1(_02961_ ), .A2(_02962_ ), .ZN(_02963_ ) );
INV_X1 _10589_ ( .A(\ID_EX_imm [30] ), .ZN(_02964_ ) );
XNOR2_X1 _10590_ ( .A(_02963_ ), .B(_02964_ ), .ZN(_02965_ ) );
OR2_X1 _10591_ ( .A1(_02942_ ), .A2(_02965_ ), .ZN(_02966_ ) );
OR2_X1 _10592_ ( .A1(_02963_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02967_ ) );
AND2_X1 _10593_ ( .A1(_02966_ ), .A2(_02967_ ), .ZN(_02968_ ) );
NAND2_X1 _10594_ ( .A1(_02467_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_02969_ ) );
OR2_X1 _10595_ ( .A1(_02124_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02970_ ) );
OAI211_X1 _10596_ ( .A(_02970_ ), .B(_02130_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02971_ ) );
NOR2_X1 _10597_ ( .A1(_02179_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02972_ ) );
OAI21_X1 _10598_ ( .A(fanout_net_25 ), .B1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02973_ ) );
OAI211_X1 _10599_ ( .A(_02971_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .C1(_02972_ ), .C2(_02973_ ), .ZN(_02974_ ) );
MUX2_X1 _10600_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02975_ ) );
MUX2_X1 _10601_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02976_ ) );
MUX2_X1 _10602_ ( .A(_02975_ ), .B(_02976_ ), .S(fanout_net_25 ), .Z(_02977_ ) );
OAI211_X1 _10603_ ( .A(_02974_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .C1(_02977_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02978_ ) );
OR2_X1 _10604_ ( .A1(_02124_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02979_ ) );
OAI211_X1 _10605_ ( .A(_02979_ ), .B(_02130_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02980_ ) );
OR2_X1 _10606_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02981_ ) );
OAI211_X1 _10607_ ( .A(_02981_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02153_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02982_ ) );
NAND3_X1 _10608_ ( .A1(_02980_ ), .A2(_02138_ ), .A3(_02982_ ), .ZN(_02983_ ) );
MUX2_X1 _10609_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02984_ ) );
MUX2_X1 _10610_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02985_ ) );
MUX2_X1 _10611_ ( .A(_02984_ ), .B(_02985_ ), .S(_02144_ ), .Z(_02986_ ) );
OAI211_X1 _10612_ ( .A(_02120_ ), .B(_02983_ ), .C1(_02986_ ), .C2(_02147_ ), .ZN(_02987_ ) );
NAND2_X1 _10613_ ( .A1(_02978_ ), .A2(_02987_ ), .ZN(_02988_ ) );
OAI21_X1 _10614_ ( .A(_02988_ ), .B1(_02162_ ), .B2(_02165_ ), .ZN(_02989_ ) );
AND2_X2 _10615_ ( .A1(_02969_ ), .A2(_02989_ ), .ZN(_02990_ ) );
XNOR2_X1 _10616_ ( .A(_02990_ ), .B(\ID_EX_imm [31] ), .ZN(_02991_ ) );
XNOR2_X1 _10617_ ( .A(_02968_ ), .B(_02991_ ), .ZN(_02992_ ) );
AND2_X2 _10618_ ( .A1(\ID_EX_typ [7] ), .A2(\ID_EX_typ [6] ), .ZN(_02993_ ) );
BUF_X4 _10619_ ( .A(_02993_ ), .Z(_02994_ ) );
NOR2_X1 _10620_ ( .A1(_02992_ ), .A2(_02994_ ), .ZN(_00097_ ) );
XNOR2_X1 _10621_ ( .A(_02942_ ), .B(_02965_ ), .ZN(_02995_ ) );
NOR2_X1 _10622_ ( .A1(_02995_ ), .A2(_02994_ ), .ZN(_00098_ ) );
AOI21_X1 _10623_ ( .A(_02420_ ), .B1(_02818_ ), .B2(_02836_ ), .ZN(_02996_ ) );
INV_X1 _10624_ ( .A(_02847_ ), .ZN(_02997_ ) );
OAI21_X1 _10625_ ( .A(_02296_ ), .B1(_02996_ ), .B2(_02997_ ), .ZN(_02998_ ) );
NAND2_X1 _10626_ ( .A1(_02998_ ), .A2(_02850_ ), .ZN(_02999_ ) );
XNOR2_X1 _10627_ ( .A(_02999_ ), .B(_02320_ ), .ZN(_03000_ ) );
NOR2_X1 _10628_ ( .A1(_03000_ ), .A2(_02994_ ), .ZN(_00099_ ) );
OR3_X1 _10629_ ( .A1(_02996_ ), .A2(_02296_ ), .A3(_02997_ ), .ZN(_03001_ ) );
INV_X1 _10630_ ( .A(_02993_ ), .ZN(_03002_ ) );
CLKBUF_X2 _10631_ ( .A(_03002_ ), .Z(_03003_ ) );
AND3_X1 _10632_ ( .A1(_03001_ ), .A2(_03003_ ), .A3(_02998_ ), .ZN(_00100_ ) );
INV_X1 _10633_ ( .A(_02419_ ), .ZN(_03004_ ) );
AOI21_X1 _10634_ ( .A(_03004_ ), .B1(_02818_ ), .B2(_02836_ ), .ZN(_03005_ ) );
AND2_X1 _10635_ ( .A1(_03005_ ), .A2(_02396_ ), .ZN(_03006_ ) );
OAI21_X1 _10636_ ( .A(_02348_ ), .B1(_03006_ ), .B2(_02842_ ), .ZN(_03007_ ) );
INV_X1 _10637_ ( .A(_02845_ ), .ZN(_03008_ ) );
NAND2_X1 _10638_ ( .A1(_03007_ ), .A2(_03008_ ), .ZN(_03009_ ) );
XNOR2_X1 _10639_ ( .A(_03009_ ), .B(_02372_ ), .ZN(_03010_ ) );
NOR2_X1 _10640_ ( .A1(_03010_ ), .A2(_02994_ ), .ZN(_00101_ ) );
NOR2_X1 _10641_ ( .A1(_03006_ ), .A2(_02842_ ), .ZN(_03011_ ) );
XNOR2_X1 _10642_ ( .A(_03011_ ), .B(_02348_ ), .ZN(_03012_ ) );
AND2_X1 _10643_ ( .A1(_03012_ ), .A2(_03003_ ), .ZN(_00102_ ) );
OR2_X1 _10644_ ( .A1(_03005_ ), .A2(_02839_ ), .ZN(_03013_ ) );
XNOR2_X1 _10645_ ( .A(_03013_ ), .B(_02396_ ), .ZN(_03014_ ) );
NOR2_X1 _10646_ ( .A1(_03014_ ), .A2(_02994_ ), .ZN(_00103_ ) );
AND3_X1 _10647_ ( .A1(_02818_ ), .A2(_02836_ ), .A3(_03004_ ), .ZN(_03015_ ) );
NOR3_X1 _10648_ ( .A1(_03015_ ), .A2(_03005_ ), .A3(_02993_ ), .ZN(_00104_ ) );
INV_X1 _10649_ ( .A(_02673_ ), .ZN(_03016_ ) );
INV_X1 _10650_ ( .A(_02816_ ), .ZN(_03017_ ) );
AOI21_X1 _10651_ ( .A(_03017_ ), .B1(_02616_ ), .B2(_02624_ ), .ZN(_03018_ ) );
INV_X1 _10652_ ( .A(_03018_ ), .ZN(_03019_ ) );
AOI21_X1 _10653_ ( .A(_03016_ ), .B1(_03019_ ), .B2(_02827_ ), .ZN(_03020_ ) );
OR2_X1 _10654_ ( .A1(_03020_ ), .A2(_02833_ ), .ZN(_03021_ ) );
AND2_X1 _10655_ ( .A1(_03021_ ), .A2(_02719_ ), .ZN(_03022_ ) );
AND2_X1 _10656_ ( .A1(_02718_ ), .A2(\ID_EX_imm [14] ), .ZN(_03023_ ) );
OR2_X1 _10657_ ( .A1(_03022_ ), .A2(_03023_ ), .ZN(_03024_ ) );
XNOR2_X1 _10658_ ( .A(_03024_ ), .B(_02696_ ), .ZN(_03025_ ) );
NOR2_X1 _10659_ ( .A1(_03025_ ), .A2(_02994_ ), .ZN(_00105_ ) );
XOR2_X1 _10660_ ( .A(_03021_ ), .B(_02719_ ), .Z(_03026_ ) );
AND2_X1 _10661_ ( .A1(_03026_ ), .A2(_03003_ ), .ZN(_00106_ ) );
OAI21_X1 _10662_ ( .A(_02649_ ), .B1(_03018_ ), .B2(_02828_ ), .ZN(_03027_ ) );
NAND2_X1 _10663_ ( .A1(_03027_ ), .A2(_02831_ ), .ZN(_03028_ ) );
XNOR2_X1 _10664_ ( .A(_03028_ ), .B(_02672_ ), .ZN(_03029_ ) );
NOR2_X1 _10665_ ( .A1(_03029_ ), .A2(_02994_ ), .ZN(_00107_ ) );
OR3_X1 _10666_ ( .A1(_03018_ ), .A2(_02649_ ), .A3(_02828_ ), .ZN(_03030_ ) );
AND3_X1 _10667_ ( .A1(_03030_ ), .A2(_03003_ ), .A3(_03027_ ), .ZN(_00108_ ) );
OR2_X1 _10668_ ( .A1(_02913_ ), .A2(_02938_ ), .ZN(_03031_ ) );
XNOR2_X1 _10669_ ( .A(_03031_ ), .B(_02936_ ), .ZN(_03032_ ) );
NOR2_X1 _10670_ ( .A1(_03032_ ), .A2(_02994_ ), .ZN(_00109_ ) );
AND3_X1 _10671_ ( .A1(_02909_ ), .A2(_02912_ ), .A3(_02168_ ), .ZN(_03033_ ) );
NOR3_X1 _10672_ ( .A1(_03033_ ), .A2(_02913_ ), .A3(_02993_ ), .ZN(_00110_ ) );
OAI21_X1 _10673_ ( .A(_02198_ ), .B1(_02902_ ), .B2(_02908_ ), .ZN(_03034_ ) );
NAND2_X1 _10674_ ( .A1(_03034_ ), .A2(_02910_ ), .ZN(_03035_ ) );
XNOR2_X1 _10675_ ( .A(_03035_ ), .B(_02223_ ), .ZN(_03036_ ) );
NOR2_X1 _10676_ ( .A1(_03036_ ), .A2(_02994_ ), .ZN(_00111_ ) );
OR3_X1 _10677_ ( .A1(_02902_ ), .A2(_02198_ ), .A3(_02908_ ), .ZN(_03037_ ) );
AND3_X1 _10678_ ( .A1(_03037_ ), .A2(_03003_ ), .A3(_03034_ ), .ZN(_00112_ ) );
NAND2_X1 _10679_ ( .A1(_02855_ ), .A2(_02878_ ), .ZN(_03038_ ) );
NAND2_X1 _10680_ ( .A1(_03038_ ), .A2(_02905_ ), .ZN(_03039_ ) );
XNOR2_X1 _10681_ ( .A(_03039_ ), .B(_02901_ ), .ZN(_03040_ ) );
NOR2_X1 _10682_ ( .A1(_03040_ ), .A2(_02994_ ), .ZN(_00113_ ) );
XOR2_X1 _10683_ ( .A(_02855_ ), .B(_02878_ ), .Z(_03041_ ) );
AND2_X1 _10684_ ( .A1(_03041_ ), .A2(_03003_ ), .ZN(_00114_ ) );
OAI21_X1 _10685_ ( .A(_02321_ ), .B1(_02996_ ), .B2(_02997_ ), .ZN(_03042_ ) );
INV_X1 _10686_ ( .A(_03042_ ), .ZN(_03043_ ) );
OR2_X1 _10687_ ( .A1(_03043_ ), .A2(_02852_ ), .ZN(_03044_ ) );
AND2_X1 _10688_ ( .A1(_03044_ ), .A2(_02272_ ), .ZN(_03045_ ) );
AND2_X1 _10689_ ( .A1(_02270_ ), .A2(\ID_EX_imm [22] ), .ZN(_03046_ ) );
OR2_X1 _10690_ ( .A1(_03045_ ), .A2(_03046_ ), .ZN(_03047_ ) );
XNOR2_X1 _10691_ ( .A(_03047_ ), .B(_02249_ ), .ZN(_03048_ ) );
NOR2_X1 _10692_ ( .A1(_03048_ ), .A2(_02993_ ), .ZN(_00115_ ) );
XOR2_X1 _10693_ ( .A(_03044_ ), .B(_02272_ ), .Z(_03049_ ) );
AND2_X1 _10694_ ( .A1(_03049_ ), .A2(_03003_ ), .ZN(_00116_ ) );
AND2_X1 _10695_ ( .A1(\IF_ID_inst [0] ), .A2(\IF_ID_inst [1] ), .ZN(_03050_ ) );
NOR2_X1 _10696_ ( .A1(\IF_ID_inst [3] ), .A2(\IF_ID_inst [2] ), .ZN(_03051_ ) );
AND2_X2 _10697_ ( .A1(_03050_ ), .A2(_03051_ ), .ZN(_03052_ ) );
CLKBUF_X2 _10698_ ( .A(_03052_ ), .Z(_03053_ ) );
INV_X1 _10699_ ( .A(_03053_ ), .ZN(_03054_ ) );
AND2_X1 _10700_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03055_ ) );
CLKBUF_X2 _10701_ ( .A(_03055_ ), .Z(_03056_ ) );
INV_X1 _10702_ ( .A(\IF_ID_inst [12] ), .ZN(_03057_ ) );
NAND4_X1 _10703_ ( .A1(_03056_ ), .A2(\IF_ID_inst [13] ), .A3(_03057_ ), .A4(\IF_ID_inst [6] ), .ZN(_03058_ ) );
NOR2_X1 _10704_ ( .A1(_03054_ ), .A2(_03058_ ), .ZN(_03059_ ) );
AND4_X1 _10705_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [6] ), .ZN(_03060_ ) );
AND2_X2 _10706_ ( .A1(_03053_ ), .A2(_03060_ ), .ZN(_03061_ ) );
NOR2_X1 _10707_ ( .A1(_03059_ ), .A2(_03061_ ), .ZN(_03062_ ) );
BUF_X4 _10708_ ( .A(_03062_ ), .Z(_03063_ ) );
INV_X1 _10709_ ( .A(\IF_ID_inst [31] ), .ZN(_03064_ ) );
NOR2_X1 _10710_ ( .A1(fanout_net_2 ), .A2(excp_written ), .ZN(_03065_ ) );
AND2_X2 _10711_ ( .A1(_02080_ ), .A2(_03065_ ), .ZN(_03066_ ) );
INV_X2 _10712_ ( .A(_03066_ ), .ZN(_03067_ ) );
BUF_X4 _10713_ ( .A(_03067_ ), .Z(_03068_ ) );
NOR3_X1 _10714_ ( .A1(_03063_ ), .A2(_03064_ ), .A3(_03068_ ), .ZN(_00195_ ) );
INV_X1 _10715_ ( .A(\IF_ID_inst [30] ), .ZN(_03069_ ) );
NOR3_X1 _10716_ ( .A1(_03063_ ), .A2(_03069_ ), .A3(_03068_ ), .ZN(_00196_ ) );
INV_X1 _10717_ ( .A(\IF_ID_inst [21] ), .ZN(_03070_ ) );
NOR3_X1 _10718_ ( .A1(_03063_ ), .A2(_03070_ ), .A3(_03068_ ), .ZN(_00197_ ) );
BUF_X4 _10719_ ( .A(_03067_ ), .Z(_03071_ ) );
INV_X1 _10720_ ( .A(_03062_ ), .ZN(_03072_ ) );
INV_X1 _10721_ ( .A(\IF_ID_inst [20] ), .ZN(_03073_ ) );
AOI21_X1 _10722_ ( .A(_03071_ ), .B1(_03072_ ), .B2(_03073_ ), .ZN(_00198_ ) );
INV_X1 _10723_ ( .A(\IF_ID_inst [29] ), .ZN(_03074_ ) );
AOI21_X1 _10724_ ( .A(_03071_ ), .B1(_03072_ ), .B2(_03074_ ), .ZN(_00199_ ) );
INV_X1 _10725_ ( .A(\IF_ID_inst [28] ), .ZN(_03075_ ) );
AOI21_X1 _10726_ ( .A(_03071_ ), .B1(_03072_ ), .B2(_03075_ ), .ZN(_00200_ ) );
INV_X1 _10727_ ( .A(\IF_ID_inst [27] ), .ZN(_03076_ ) );
NOR3_X1 _10728_ ( .A1(_03063_ ), .A2(_03076_ ), .A3(_03068_ ), .ZN(_00201_ ) );
INV_X1 _10729_ ( .A(\IF_ID_inst [26] ), .ZN(_03077_ ) );
AOI21_X1 _10730_ ( .A(_03071_ ), .B1(_03072_ ), .B2(_03077_ ), .ZN(_00202_ ) );
INV_X1 _10731_ ( .A(\IF_ID_inst [25] ), .ZN(_03078_ ) );
BUF_X4 _10732_ ( .A(_03067_ ), .Z(_03079_ ) );
NOR3_X1 _10733_ ( .A1(_03063_ ), .A2(_03078_ ), .A3(_03079_ ), .ZN(_00203_ ) );
INV_X1 _10734_ ( .A(\IF_ID_inst [24] ), .ZN(_03080_ ) );
NOR3_X1 _10735_ ( .A1(_03063_ ), .A2(_03080_ ), .A3(_03079_ ), .ZN(_00204_ ) );
INV_X1 _10736_ ( .A(\IF_ID_inst [23] ), .ZN(_03081_ ) );
NOR3_X1 _10737_ ( .A1(_03063_ ), .A2(_03081_ ), .A3(_03079_ ), .ZN(_00205_ ) );
INV_X1 _10738_ ( .A(\IF_ID_inst [22] ), .ZN(_03082_ ) );
NOR3_X1 _10739_ ( .A1(_03063_ ), .A2(_03082_ ), .A3(_03079_ ), .ZN(_00206_ ) );
CLKBUF_X2 _10740_ ( .A(_03065_ ), .Z(_03083_ ) );
AND3_X1 _10741_ ( .A1(_02080_ ), .A2(_03083_ ), .A3(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ), .ZN(_00207_ ) );
AND3_X1 _10742_ ( .A1(_02080_ ), .A2(_03083_ ), .A3(\myidu.state [2] ), .ZN(_00208_ ) );
AND3_X1 _10743_ ( .A1(_03050_ ), .A2(\IF_ID_inst [3] ), .A3(\IF_ID_inst [2] ), .ZN(_03084_ ) );
INV_X1 _10744_ ( .A(_03084_ ), .ZN(_03085_ ) );
NOR2_X1 _10745_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_03086_ ) );
NOR2_X1 _10746_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03087_ ) );
INV_X1 _10747_ ( .A(\IF_ID_inst [6] ), .ZN(_03088_ ) );
NAND4_X1 _10748_ ( .A1(_03086_ ), .A2(_03087_ ), .A3(\IF_ID_inst [12] ), .A4(_03088_ ), .ZN(_03089_ ) );
NOR2_X1 _10749_ ( .A1(_03085_ ), .A2(_03089_ ), .ZN(_03090_ ) );
INV_X1 _10750_ ( .A(_03090_ ), .ZN(_03091_ ) );
INV_X1 _10751_ ( .A(\IF_ID_inst [7] ), .ZN(_03092_ ) );
INV_X1 _10752_ ( .A(\IF_ID_inst [15] ), .ZN(_03093_ ) );
AND4_X1 _10753_ ( .A1(_03057_ ), .A2(_03092_ ), .A3(_03093_ ), .A4(\IF_ID_inst [6] ), .ZN(_03094_ ) );
AND3_X1 _10754_ ( .A1(_03094_ ), .A2(_03055_ ), .A3(_03086_ ), .ZN(_03095_ ) );
INV_X1 _10755_ ( .A(\IF_ID_inst [11] ), .ZN(_03096_ ) );
INV_X1 _10756_ ( .A(\IF_ID_inst [10] ), .ZN(_03097_ ) );
INV_X1 _10757_ ( .A(\IF_ID_inst [9] ), .ZN(_03098_ ) );
NAND3_X1 _10758_ ( .A1(_03096_ ), .A2(_03097_ ), .A3(_03098_ ), .ZN(_03099_ ) );
NOR2_X1 _10759_ ( .A1(_03099_ ), .A2(\IF_ID_inst [8] ), .ZN(_03100_ ) );
NAND3_X1 _10760_ ( .A1(_03095_ ), .A2(_03053_ ), .A3(_03100_ ), .ZN(_03101_ ) );
INV_X1 _10761_ ( .A(_03101_ ), .ZN(_03102_ ) );
NOR2_X1 _10762_ ( .A1(\IF_ID_inst [19] ), .A2(\IF_ID_inst [18] ), .ZN(_03103_ ) );
NOR2_X1 _10763_ ( .A1(\IF_ID_inst [17] ), .A2(\IF_ID_inst [16] ), .ZN(_03104_ ) );
NOR2_X1 _10764_ ( .A1(\IF_ID_inst [23] ), .A2(\IF_ID_inst [22] ), .ZN(_03105_ ) );
AND3_X1 _10765_ ( .A1(_03103_ ), .A2(_03104_ ), .A3(_03105_ ), .ZN(_03106_ ) );
AND3_X1 _10766_ ( .A1(_03106_ ), .A2(_03070_ ), .A3(\IF_ID_inst [20] ), .ZN(_03107_ ) );
NOR2_X1 _10767_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .ZN(_03108_ ) );
NAND4_X1 _10768_ ( .A1(_03108_ ), .A2(_03076_ ), .A3(_03080_ ), .A4(_03064_ ), .ZN(_03109_ ) );
NAND3_X1 _10769_ ( .A1(_03069_ ), .A2(_03074_ ), .A3(_03075_ ), .ZN(_03110_ ) );
NOR2_X1 _10770_ ( .A1(_03109_ ), .A2(_03110_ ), .ZN(_03111_ ) );
NAND3_X1 _10771_ ( .A1(_03102_ ), .A2(_03107_ ), .A3(_03111_ ), .ZN(_03112_ ) );
INV_X1 _10772_ ( .A(\IF_ID_inst [5] ), .ZN(_03113_ ) );
NOR2_X1 _10773_ ( .A1(_03113_ ), .A2(\IF_ID_inst [4] ), .ZN(_03114_ ) );
NOR2_X1 _10774_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_03115_ ) );
AND3_X1 _10775_ ( .A1(_03052_ ), .A2(_03114_ ), .A3(_03115_ ), .ZN(_03116_ ) );
INV_X1 _10776_ ( .A(\IF_ID_inst [13] ), .ZN(_03117_ ) );
NOR2_X1 _10777_ ( .A1(_03117_ ), .A2(\IF_ID_inst [14] ), .ZN(_03118_ ) );
AND2_X1 _10778_ ( .A1(_03116_ ), .A2(_03118_ ), .ZN(_03119_ ) );
INV_X1 _10779_ ( .A(_03119_ ), .ZN(_03120_ ) );
NOR2_X1 _10780_ ( .A1(_03057_ ), .A2(\IF_ID_inst [6] ), .ZN(_03121_ ) );
BUF_X2 _10781_ ( .A(_03086_ ), .Z(_03122_ ) );
NAND3_X1 _10782_ ( .A1(_03114_ ), .A2(_03121_ ), .A3(_03122_ ), .ZN(_03123_ ) );
NOR2_X1 _10783_ ( .A1(_03054_ ), .A2(_03123_ ), .ZN(_03124_ ) );
AOI21_X1 _10784_ ( .A(_03124_ ), .B1(_03122_ ), .B2(_03116_ ), .ZN(_03125_ ) );
AND4_X1 _10785_ ( .A1(_03091_ ), .A2(_03112_ ), .A3(_03120_ ), .A4(_03125_ ), .ZN(_03126_ ) );
BUF_X2 _10786_ ( .A(_03066_ ), .Z(_03127_ ) );
INV_X1 _10787_ ( .A(\IF_ID_inst [4] ), .ZN(_03128_ ) );
NAND4_X1 _10788_ ( .A1(_03128_ ), .A2(\IF_ID_inst [5] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [6] ), .ZN(_03129_ ) );
NOR2_X1 _10789_ ( .A1(_03054_ ), .A2(_03129_ ), .ZN(_03130_ ) );
AND2_X1 _10790_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_03131_ ) );
NAND2_X1 _10791_ ( .A1(_03130_ ), .A2(_03131_ ), .ZN(_03132_ ) );
NOR2_X1 _10792_ ( .A1(_03088_ ), .A2(\IF_ID_inst [12] ), .ZN(_03133_ ) );
AND2_X1 _10793_ ( .A1(_03133_ ), .A2(_03114_ ), .ZN(_03134_ ) );
AND2_X1 _10794_ ( .A1(_03134_ ), .A2(_03053_ ), .ZN(_03135_ ) );
AND2_X1 _10795_ ( .A1(_03135_ ), .A2(\IF_ID_inst [14] ), .ZN(_03136_ ) );
NOR3_X1 _10796_ ( .A1(_03054_ ), .A2(\IF_ID_inst [13] ), .A3(_03129_ ), .ZN(_03137_ ) );
NOR2_X1 _10797_ ( .A1(_03136_ ), .A2(_03137_ ), .ZN(_03138_ ) );
AND2_X1 _10798_ ( .A1(_03103_ ), .A2(_03104_ ), .ZN(_03139_ ) );
NAND3_X1 _10799_ ( .A1(_03077_ ), .A2(_03078_ ), .A3(_03080_ ), .ZN(_03140_ ) );
NOR2_X1 _10800_ ( .A1(_03140_ ), .A2(\IF_ID_inst [27] ), .ZN(_03141_ ) );
NAND2_X1 _10801_ ( .A1(_03069_ ), .A2(\IF_ID_inst [29] ), .ZN(_03142_ ) );
NOR3_X1 _10802_ ( .A1(_03142_ ), .A2(_03075_ ), .A3(\IF_ID_inst [31] ), .ZN(_03143_ ) );
AND3_X1 _10803_ ( .A1(_03105_ ), .A2(\IF_ID_inst [21] ), .A3(_03073_ ), .ZN(_03144_ ) );
AND4_X1 _10804_ ( .A1(_03139_ ), .A2(_03141_ ), .A3(_03143_ ), .A4(_03144_ ), .ZN(_03145_ ) );
NAND2_X1 _10805_ ( .A1(_03102_ ), .A2(_03145_ ), .ZN(_03146_ ) );
NAND3_X1 _10806_ ( .A1(_03134_ ), .A2(_03053_ ), .A3(_03122_ ), .ZN(_03147_ ) );
AND4_X1 _10807_ ( .A1(_03132_ ), .A2(_03138_ ), .A3(_03146_ ), .A4(_03147_ ), .ZN(_03148_ ) );
AND4_X1 _10808_ ( .A1(\IF_ID_inst [11] ), .A2(_03126_ ), .A3(_03127_ ), .A4(_03148_ ), .ZN(_00209_ ) );
AND4_X1 _10809_ ( .A1(\IF_ID_inst [10] ), .A2(_03126_ ), .A3(_03127_ ), .A4(_03148_ ), .ZN(_00210_ ) );
AND4_X1 _10810_ ( .A1(\IF_ID_inst [9] ), .A2(_03126_ ), .A3(_03127_ ), .A4(_03148_ ), .ZN(_00211_ ) );
AND4_X1 _10811_ ( .A1(\IF_ID_inst [8] ), .A2(_03126_ ), .A3(_03066_ ), .A4(_03148_ ), .ZN(_00212_ ) );
AND4_X1 _10812_ ( .A1(\IF_ID_inst [7] ), .A2(_03126_ ), .A3(_03066_ ), .A4(_03148_ ), .ZN(_00213_ ) );
AND4_X1 _10813_ ( .A1(\IF_ID_inst [6] ), .A2(_03052_ ), .A3(_03092_ ), .A4(_03055_ ), .ZN(_03149_ ) );
NOR4_X1 _10814_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [15] ), .ZN(_03150_ ) );
AND3_X1 _10815_ ( .A1(_03149_ ), .A2(_03100_ ), .A3(_03150_ ), .ZN(_03151_ ) );
AND4_X1 _10816_ ( .A1(_03070_ ), .A2(_03111_ ), .A3(\IF_ID_inst [20] ), .A4(_03106_ ), .ZN(_03152_ ) );
AND2_X1 _10817_ ( .A1(_03151_ ), .A2(_03152_ ), .ZN(_03153_ ) );
AND3_X1 _10818_ ( .A1(_03087_ ), .A2(\IF_ID_inst [12] ), .A3(_03088_ ), .ZN(_03154_ ) );
AND2_X1 _10819_ ( .A1(_03084_ ), .A2(_03154_ ), .ZN(_03155_ ) );
AOI21_X1 _10820_ ( .A(_03153_ ), .B1(_03086_ ), .B2(_03155_ ), .ZN(_03156_ ) );
INV_X1 _10821_ ( .A(_03156_ ), .ZN(_03157_ ) );
INV_X1 _10822_ ( .A(\IF_ID_inst [19] ), .ZN(_03158_ ) );
INV_X1 _10823_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03159_ ) );
AND2_X1 _10824_ ( .A1(_03114_ ), .A2(_03159_ ), .ZN(_03160_ ) );
AND2_X1 _10825_ ( .A1(_03160_ ), .A2(_03084_ ), .ZN(_03161_ ) );
CLKBUF_X2 _10826_ ( .A(_03161_ ), .Z(_03162_ ) );
BUF_X2 _10827_ ( .A(_03162_ ), .Z(_03163_ ) );
NAND3_X1 _10828_ ( .A1(\IF_ID_inst [2] ), .A2(\IF_ID_inst [0] ), .A3(\IF_ID_inst [1] ), .ZN(_03164_ ) );
NOR2_X1 _10829_ ( .A1(_03164_ ), .A2(\IF_ID_inst [3] ), .ZN(_03165_ ) );
NOR2_X1 _10830_ ( .A1(_03128_ ), .A2(\IF_ID_inst [6] ), .ZN(_03166_ ) );
AND2_X1 _10831_ ( .A1(_03165_ ), .A2(_03166_ ), .ZN(_03167_ ) );
NOR2_X2 _10832_ ( .A1(_03163_ ), .A2(_03167_ ), .ZN(_03168_ ) );
INV_X1 _10833_ ( .A(_03145_ ), .ZN(_03169_ ) );
OAI21_X1 _10834_ ( .A(_03168_ ), .B1(_03169_ ), .B2(_03101_ ), .ZN(_03170_ ) );
NOR4_X1 _10835_ ( .A1(_03157_ ), .A2(_03158_ ), .A3(_03079_ ), .A4(_03170_ ), .ZN(_00214_ ) );
INV_X1 _10836_ ( .A(\IF_ID_inst [18] ), .ZN(_03171_ ) );
NOR4_X1 _10837_ ( .A1(_03157_ ), .A2(_03171_ ), .A3(_03079_ ), .A4(_03170_ ), .ZN(_00215_ ) );
INV_X1 _10838_ ( .A(\IF_ID_inst [17] ), .ZN(_03172_ ) );
NOR4_X1 _10839_ ( .A1(_03157_ ), .A2(_03172_ ), .A3(_03079_ ), .A4(_03170_ ), .ZN(_00216_ ) );
XNOR2_X1 _10840_ ( .A(\IF_ID_pc [14] ), .B(\myexu.pc_jump [14] ), .ZN(_03173_ ) );
XNOR2_X1 _10841_ ( .A(\IF_ID_pc [15] ), .B(\myexu.pc_jump [15] ), .ZN(_03174_ ) );
XNOR2_X1 _10842_ ( .A(\IF_ID_pc [10] ), .B(\myexu.pc_jump [10] ), .ZN(_03175_ ) );
XNOR2_X1 _10843_ ( .A(\IF_ID_pc [11] ), .B(\myexu.pc_jump [11] ), .ZN(_03176_ ) );
AND4_X1 _10844_ ( .A1(_03173_ ), .A2(_03174_ ), .A3(_03175_ ), .A4(_03176_ ), .ZN(_03177_ ) );
XNOR2_X1 _10845_ ( .A(\IF_ID_pc [5] ), .B(\myexu.pc_jump [5] ), .ZN(_03178_ ) );
XNOR2_X1 _10846_ ( .A(\myexu.pc_jump [0] ), .B(\IF_ID_pc [0] ), .ZN(_03179_ ) );
XNOR2_X1 _10847_ ( .A(\myexu.pc_jump [1] ), .B(\IF_ID_pc [1] ), .ZN(_03180_ ) );
XNOR2_X1 _10848_ ( .A(fanout_net_11 ), .B(\myexu.pc_jump [4] ), .ZN(_03181_ ) );
AND4_X1 _10849_ ( .A1(_03178_ ), .A2(_03179_ ), .A3(_03180_ ), .A4(_03181_ ), .ZN(_03182_ ) );
XNOR2_X1 _10850_ ( .A(\IF_ID_pc [20] ), .B(\myexu.pc_jump [20] ), .ZN(_03183_ ) );
XNOR2_X1 _10851_ ( .A(\IF_ID_pc [16] ), .B(\myexu.pc_jump [16] ), .ZN(_03184_ ) );
XNOR2_X1 _10852_ ( .A(\IF_ID_pc [17] ), .B(\myexu.pc_jump [17] ), .ZN(_03185_ ) );
XNOR2_X1 _10853_ ( .A(\IF_ID_pc [21] ), .B(\myexu.pc_jump [21] ), .ZN(_03186_ ) );
AND4_X1 _10854_ ( .A1(_03183_ ), .A2(_03184_ ), .A3(_03185_ ), .A4(_03186_ ), .ZN(_03187_ ) );
XNOR2_X1 _10855_ ( .A(\IF_ID_pc [30] ), .B(\myexu.pc_jump [30] ), .ZN(_03188_ ) );
XNOR2_X1 _10856_ ( .A(\IF_ID_pc [31] ), .B(\myexu.pc_jump [31] ), .ZN(_03189_ ) );
XNOR2_X1 _10857_ ( .A(\IF_ID_pc [26] ), .B(\myexu.pc_jump [26] ), .ZN(_03190_ ) );
XNOR2_X1 _10858_ ( .A(\IF_ID_pc [27] ), .B(\myexu.pc_jump [27] ), .ZN(_03191_ ) );
AND4_X1 _10859_ ( .A1(_03188_ ), .A2(_03189_ ), .A3(_03190_ ), .A4(_03191_ ), .ZN(_03192_ ) );
NAND4_X1 _10860_ ( .A1(_03177_ ), .A2(_03182_ ), .A3(_03187_ ), .A4(_03192_ ), .ZN(_03193_ ) );
XNOR2_X1 _10861_ ( .A(\IF_ID_pc [18] ), .B(\myexu.pc_jump [18] ), .ZN(_03194_ ) );
XNOR2_X1 _10862_ ( .A(\IF_ID_pc [19] ), .B(\myexu.pc_jump [19] ), .ZN(_03195_ ) );
XNOR2_X1 _10863_ ( .A(\IF_ID_pc [23] ), .B(\myexu.pc_jump [23] ), .ZN(_03196_ ) );
XNOR2_X1 _10864_ ( .A(\IF_ID_pc [22] ), .B(\myexu.pc_jump [22] ), .ZN(_03197_ ) );
NAND4_X1 _10865_ ( .A1(_03194_ ), .A2(_03195_ ), .A3(_03196_ ), .A4(_03197_ ), .ZN(_03198_ ) );
XNOR2_X1 _10866_ ( .A(\IF_ID_pc [24] ), .B(\myexu.pc_jump [24] ), .ZN(_03199_ ) );
XNOR2_X1 _10867_ ( .A(\IF_ID_pc [28] ), .B(\myexu.pc_jump [28] ), .ZN(_03200_ ) );
XNOR2_X1 _10868_ ( .A(\IF_ID_pc [29] ), .B(\myexu.pc_jump [29] ), .ZN(_03201_ ) );
XNOR2_X1 _10869_ ( .A(\IF_ID_pc [25] ), .B(\myexu.pc_jump [25] ), .ZN(_03202_ ) );
NAND4_X1 _10870_ ( .A1(_03199_ ), .A2(_03200_ ), .A3(_03201_ ), .A4(_03202_ ), .ZN(_03203_ ) );
NOR3_X1 _10871_ ( .A1(_03193_ ), .A2(_03198_ ), .A3(_03203_ ), .ZN(_03204_ ) );
XNOR2_X1 _10872_ ( .A(\IF_ID_pc [8] ), .B(\myexu.pc_jump [8] ), .ZN(_03205_ ) );
XNOR2_X1 _10873_ ( .A(\IF_ID_pc [13] ), .B(\myexu.pc_jump [13] ), .ZN(_03206_ ) );
XNOR2_X1 _10874_ ( .A(\IF_ID_pc [9] ), .B(\myexu.pc_jump [9] ), .ZN(_03207_ ) );
XNOR2_X1 _10875_ ( .A(\IF_ID_pc [12] ), .B(\myexu.pc_jump [12] ), .ZN(_03208_ ) );
AND4_X1 _10876_ ( .A1(_03205_ ), .A2(_03206_ ), .A3(_03207_ ), .A4(_03208_ ), .ZN(_03209_ ) );
XNOR2_X1 _10877_ ( .A(\IF_ID_pc [6] ), .B(\myexu.pc_jump [6] ), .ZN(_03210_ ) );
XNOR2_X1 _10878_ ( .A(\IF_ID_pc [7] ), .B(\myexu.pc_jump [7] ), .ZN(_03211_ ) );
XNOR2_X1 _10879_ ( .A(fanout_net_7 ), .B(\myexu.pc_jump [3] ), .ZN(_03212_ ) );
XNOR2_X1 _10880_ ( .A(\myexu.pc_jump [2] ), .B(\IF_ID_pc [2] ), .ZN(_03213_ ) );
AND4_X1 _10881_ ( .A1(_03210_ ), .A2(_03211_ ), .A3(_03212_ ), .A4(_03213_ ), .ZN(_03214_ ) );
AND3_X1 _10882_ ( .A1(_03204_ ), .A2(_03209_ ), .A3(_03214_ ), .ZN(_03215_ ) );
INV_X1 _10883_ ( .A(check_quest ), .ZN(_03216_ ) );
NOR2_X1 _10884_ ( .A1(_03215_ ), .A2(_03216_ ), .ZN(_03217_ ) );
INV_X1 _10885_ ( .A(\myifu.state [1] ), .ZN(_03218_ ) );
NOR2_X1 _10886_ ( .A1(_03218_ ), .A2(fanout_net_41 ), .ZN(_03219_ ) );
INV_X1 _10887_ ( .A(_03219_ ), .ZN(_03220_ ) );
NOR2_X1 _10888_ ( .A1(_03217_ ), .A2(_03220_ ), .ZN(_03221_ ) );
AND2_X2 _10889_ ( .A1(_03221_ ), .A2(IDU_ready_IFU ), .ZN(_03222_ ) );
INV_X1 _10890_ ( .A(_03222_ ), .ZN(_03223_ ) );
BUF_X4 _10891_ ( .A(_03223_ ), .Z(_03224_ ) );
NOR2_X1 _10892_ ( .A1(_03157_ ), .A2(_03170_ ), .ZN(_03225_ ) );
AND2_X2 _10893_ ( .A1(_03052_ ), .A2(_03115_ ), .ZN(_03226_ ) );
NAND3_X1 _10894_ ( .A1(_03226_ ), .A2(_03117_ ), .A3(_03087_ ), .ZN(_03227_ ) );
AND2_X1 _10895_ ( .A1(_03154_ ), .A2(_03052_ ), .ZN(_03228_ ) );
NAND2_X1 _10896_ ( .A1(_03228_ ), .A2(_03117_ ), .ZN(_03229_ ) );
AND2_X1 _10897_ ( .A1(_03227_ ), .A2(_03229_ ), .ZN(_03230_ ) );
NOR2_X1 _10898_ ( .A1(_03110_ ), .A2(\IF_ID_inst [27] ), .ZN(_03231_ ) );
INV_X1 _10899_ ( .A(_03231_ ), .ZN(_03232_ ) );
INV_X1 _10900_ ( .A(\IF_ID_inst [14] ), .ZN(_03233_ ) );
NAND4_X1 _10901_ ( .A1(_03108_ ), .A2(_03233_ ), .A3(\IF_ID_inst [13] ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03234_ ) );
NOR2_X1 _10902_ ( .A1(_03232_ ), .A2(_03234_ ), .ZN(_03235_ ) );
NAND3_X1 _10903_ ( .A1(_03235_ ), .A2(_03056_ ), .A3(_03226_ ), .ZN(_03236_ ) );
AND2_X1 _10904_ ( .A1(_03086_ ), .A2(_03108_ ), .ZN(_03237_ ) );
NOR2_X1 _10905_ ( .A1(_03069_ ), .A2(\IF_ID_inst [29] ), .ZN(_03238_ ) );
NOR2_X1 _10906_ ( .A1(\IF_ID_inst [28] ), .A2(\IF_ID_inst [27] ), .ZN(_03239_ ) );
AND3_X1 _10907_ ( .A1(_03238_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_03239_ ), .ZN(_03240_ ) );
NAND4_X1 _10908_ ( .A1(_03226_ ), .A2(_03056_ ), .A3(_03237_ ), .A4(_03240_ ), .ZN(_03241_ ) );
AND2_X1 _10909_ ( .A1(_03236_ ), .A2(_03241_ ), .ZN(_03242_ ) );
NOR2_X1 _10910_ ( .A1(_03128_ ), .A2(\IF_ID_inst [5] ), .ZN(_03243_ ) );
AND2_X1 _10911_ ( .A1(_03226_ ), .A2(_03243_ ), .ZN(_03244_ ) );
NAND2_X1 _10912_ ( .A1(_03244_ ), .A2(_03118_ ), .ZN(_03245_ ) );
AND4_X1 _10913_ ( .A1(\IF_ID_inst [4] ), .A2(_03113_ ), .A3(_03088_ ), .A4(\IF_ID_inst [12] ), .ZN(_03246_ ) );
AND3_X1 _10914_ ( .A1(_03053_ ), .A2(_03246_ ), .A3(\IF_ID_inst [13] ), .ZN(_03247_ ) );
INV_X1 _10915_ ( .A(_03247_ ), .ZN(_03248_ ) );
OAI21_X1 _10916_ ( .A(_03245_ ), .B1(\IF_ID_inst [14] ), .B2(_03248_ ), .ZN(_03249_ ) );
INV_X1 _10917_ ( .A(_03118_ ), .ZN(_03250_ ) );
NAND2_X1 _10918_ ( .A1(_03244_ ), .A2(_03250_ ), .ZN(_03251_ ) );
AND3_X1 _10919_ ( .A1(_03243_ ), .A2(_03050_ ), .A3(_03051_ ), .ZN(_03252_ ) );
NAND3_X1 _10920_ ( .A1(_03252_ ), .A2(_03131_ ), .A3(_03121_ ), .ZN(_03253_ ) );
NAND2_X1 _10921_ ( .A1(_03251_ ), .A2(_03253_ ), .ZN(_03254_ ) );
NOR2_X1 _10922_ ( .A1(_03249_ ), .A2(_03254_ ), .ZN(_03255_ ) );
AND4_X1 _10923_ ( .A1(_03225_ ), .A2(_03230_ ), .A3(_03242_ ), .A4(_03255_ ), .ZN(_03256_ ) );
AND2_X1 _10924_ ( .A1(_03226_ ), .A2(_03087_ ), .ZN(_03257_ ) );
AND2_X1 _10925_ ( .A1(_03257_ ), .A2(_03118_ ), .ZN(_03258_ ) );
AOI21_X1 _10926_ ( .A(_03258_ ), .B1(_03122_ ), .B2(_03135_ ), .ZN(_03259_ ) );
AND3_X1 _10927_ ( .A1(_03052_ ), .A2(_03114_ ), .A3(_03121_ ), .ZN(_03260_ ) );
OAI21_X1 _10928_ ( .A(_03086_ ), .B1(_03116_ ), .B2(_03260_ ), .ZN(_03261_ ) );
AND2_X1 _10929_ ( .A1(_03120_ ), .A2(_03261_ ), .ZN(_03262_ ) );
AND4_X1 _10930_ ( .A1(_03062_ ), .A2(_03259_ ), .A3(_03138_ ), .A4(_03262_ ), .ZN(_03263_ ) );
AND2_X1 _10931_ ( .A1(_03053_ ), .A2(_03246_ ), .ZN(_03264_ ) );
NOR2_X1 _10932_ ( .A1(_03233_ ), .A2(\IF_ID_inst [13] ), .ZN(_03265_ ) );
AND2_X1 _10933_ ( .A1(_03265_ ), .A2(_03108_ ), .ZN(_03266_ ) );
INV_X1 _10934_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03267_ ) );
NOR3_X1 _10935_ ( .A1(_03110_ ), .A2(\IF_ID_inst [27] ), .A3(_03267_ ), .ZN(_03268_ ) );
OAI211_X1 _10936_ ( .A(_03264_ ), .B(_03266_ ), .C1(_03240_ ), .C2(_03268_ ), .ZN(_03269_ ) );
AND3_X1 _10937_ ( .A1(_03134_ ), .A2(_03165_ ), .A3(_03086_ ), .ZN(_03270_ ) );
INV_X1 _10938_ ( .A(_03270_ ), .ZN(_03271_ ) );
NAND3_X1 _10939_ ( .A1(_03264_ ), .A2(_03237_ ), .A3(_03268_ ), .ZN(_03272_ ) );
AND4_X1 _10940_ ( .A1(_03132_ ), .A2(_03269_ ), .A3(_03271_ ), .A4(_03272_ ), .ZN(_03273_ ) );
AND3_X1 _10941_ ( .A1(_03256_ ), .A2(_03263_ ), .A3(_03273_ ), .ZN(_03274_ ) );
AND3_X1 _10942_ ( .A1(_03266_ ), .A2(_03231_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03275_ ) );
AND3_X1 _10943_ ( .A1(_03275_ ), .A2(_03056_ ), .A3(_03226_ ), .ZN(_03276_ ) );
AND4_X1 _10944_ ( .A1(_03056_ ), .A2(_03226_ ), .A3(_03237_ ), .A4(_03268_ ), .ZN(_03277_ ) );
NAND3_X1 _10945_ ( .A1(_03131_ ), .A2(_03108_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03278_ ) );
NOR3_X1 _10946_ ( .A1(_03278_ ), .A2(\IF_ID_inst [27] ), .A3(_03110_ ), .ZN(_03279_ ) );
AND3_X1 _10947_ ( .A1(_03226_ ), .A2(_03056_ ), .A3(_03279_ ), .ZN(_03280_ ) );
AND3_X1 _10948_ ( .A1(_03050_ ), .A2(\IF_ID_inst [12] ), .A3(_03051_ ), .ZN(_03281_ ) );
AND3_X1 _10949_ ( .A1(_03088_ ), .A2(\IF_ID_inst [4] ), .A3(\IF_ID_inst [5] ), .ZN(_03282_ ) );
AND3_X1 _10950_ ( .A1(_03279_ ), .A2(_03281_ ), .A3(_03282_ ), .ZN(_03283_ ) );
NOR4_X1 _10951_ ( .A1(_03276_ ), .A2(_03277_ ), .A3(_03280_ ), .A4(_03283_ ), .ZN(_03284_ ) );
AND2_X1 _10952_ ( .A1(_03240_ ), .A2(_03266_ ), .ZN(_03285_ ) );
AND2_X1 _10953_ ( .A1(_03281_ ), .A2(_03282_ ), .ZN(_03286_ ) );
NAND2_X1 _10954_ ( .A1(_03285_ ), .A2(_03286_ ), .ZN(_03287_ ) );
INV_X1 _10955_ ( .A(_03286_ ), .ZN(_03288_ ) );
AND4_X1 _10956_ ( .A1(\IF_ID_inst [14] ), .A2(_03108_ ), .A3(_03117_ ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03289_ ) );
AND2_X1 _10957_ ( .A1(_03289_ ), .A2(_03231_ ), .ZN(_03290_ ) );
NOR2_X1 _10958_ ( .A1(_03235_ ), .A2(_03290_ ), .ZN(_03291_ ) );
AND3_X1 _10959_ ( .A1(_03086_ ), .A2(_03108_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03292_ ) );
AND2_X1 _10960_ ( .A1(_03231_ ), .A2(_03292_ ), .ZN(_03293_ ) );
INV_X1 _10961_ ( .A(_03293_ ), .ZN(_03294_ ) );
AOI21_X1 _10962_ ( .A(_03288_ ), .B1(_03291_ ), .B2(_03294_ ), .ZN(_03295_ ) );
INV_X1 _10963_ ( .A(_03295_ ), .ZN(_03296_ ) );
AND3_X2 _10964_ ( .A1(_03284_ ), .A2(_03287_ ), .A3(_03296_ ), .ZN(_03297_ ) );
AOI221_X4 _10965_ ( .A(_03224_ ), .B1(\IF_ID_inst [18] ), .B2(_03225_ ), .C1(_03274_ ), .C2(_03297_ ), .ZN(_03298_ ) );
AND2_X1 _10966_ ( .A1(_03274_ ), .A2(_03297_ ), .ZN(_03299_ ) );
BUF_X4 _10967_ ( .A(_03299_ ), .Z(_03300_ ) );
NOR2_X1 _10968_ ( .A1(_03300_ ), .A2(_03224_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _10969_ ( .A(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_03301_ ) );
AOI211_X1 _10970_ ( .A(_03067_ ), .B(_03298_ ), .C1(_03301_ ), .C2(_02108_ ), .ZN(_00217_ ) );
INV_X1 _10971_ ( .A(\IF_ID_inst [16] ), .ZN(_03302_ ) );
NOR4_X1 _10972_ ( .A1(_03157_ ), .A2(_03302_ ), .A3(_03079_ ), .A4(_03170_ ), .ZN(_00218_ ) );
INV_X1 _10973_ ( .A(_03300_ ), .ZN(_03303_ ) );
NAND4_X1 _10974_ ( .A1(_03303_ ), .A2(\IF_ID_inst [17] ), .A3(_03225_ ), .A4(_03222_ ), .ZN(_03304_ ) );
OAI21_X1 _10975_ ( .A(\ID_EX_rs1 [2] ), .B1(_03300_ ), .B2(_03224_ ), .ZN(_03305_ ) );
AOI21_X1 _10976_ ( .A(_03071_ ), .B1(_03304_ ), .B2(_03305_ ), .ZN(_00219_ ) );
NOR4_X1 _10977_ ( .A1(_03157_ ), .A2(_03093_ ), .A3(_03079_ ), .A4(_03170_ ), .ZN(_00220_ ) );
NAND4_X1 _10978_ ( .A1(_03303_ ), .A2(\IF_ID_inst [16] ), .A3(_03225_ ), .A4(_03222_ ), .ZN(_03306_ ) );
OAI21_X1 _10979_ ( .A(\ID_EX_rs1 [1] ), .B1(_03300_ ), .B2(_03224_ ), .ZN(_03307_ ) );
AOI21_X1 _10980_ ( .A(_03071_ ), .B1(_03306_ ), .B2(_03307_ ), .ZN(_00221_ ) );
INV_X1 _10981_ ( .A(_03258_ ), .ZN(_03308_ ) );
NOR2_X1 _10982_ ( .A1(_03270_ ), .A2(_03163_ ), .ZN(_03309_ ) );
AND3_X1 _10983_ ( .A1(_03308_ ), .A2(_03230_ ), .A3(_03309_ ), .ZN(_03310_ ) );
AND3_X1 _10984_ ( .A1(_03095_ ), .A2(_03053_ ), .A3(_03100_ ), .ZN(_03311_ ) );
AND2_X1 _10985_ ( .A1(_03311_ ), .A2(_03111_ ), .ZN(_03312_ ) );
NAND2_X1 _10986_ ( .A1(_03312_ ), .A2(_03107_ ), .ZN(_03313_ ) );
NAND2_X1 _10987_ ( .A1(_03251_ ), .A2(_03248_ ), .ZN(_03314_ ) );
AND4_X1 _10988_ ( .A1(_03139_ ), .A2(_03141_ ), .A3(_03143_ ), .A4(_03144_ ), .ZN(_03315_ ) );
AND2_X1 _10989_ ( .A1(_03311_ ), .A2(_03315_ ), .ZN(_03316_ ) );
NOR3_X1 _10990_ ( .A1(_03314_ ), .A2(_03316_ ), .A3(_03090_ ), .ZN(_03317_ ) );
AND4_X1 _10991_ ( .A1(_03062_ ), .A2(_03310_ ), .A3(_03313_ ), .A4(_03317_ ), .ZN(_03318_ ) );
INV_X1 _10992_ ( .A(_03167_ ), .ZN(_03319_ ) );
AND2_X1 _10993_ ( .A1(_03245_ ), .A2(_03319_ ), .ZN(_03320_ ) );
AND2_X1 _10994_ ( .A1(_03269_ ), .A2(_03272_ ), .ZN(_03321_ ) );
AND2_X2 _10995_ ( .A1(_03320_ ), .A2(_03321_ ), .ZN(_03322_ ) );
AND4_X1 _10996_ ( .A1(\IF_ID_inst [24] ), .A2(_03318_ ), .A3(_03066_ ), .A4(_03322_ ), .ZN(_00222_ ) );
OAI21_X1 _10997_ ( .A(_03127_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs1 [0] ), .ZN(_03323_ ) );
AOI221_X4 _10998_ ( .A(_03224_ ), .B1(\IF_ID_inst [15] ), .B2(_03225_ ), .C1(_03274_ ), .C2(_03297_ ), .ZN(_03324_ ) );
NOR2_X1 _10999_ ( .A1(_03323_ ), .A2(_03324_ ), .ZN(_00223_ ) );
AND4_X1 _11000_ ( .A1(\IF_ID_inst [23] ), .A2(_03318_ ), .A3(_03066_ ), .A4(_03322_ ), .ZN(_00224_ ) );
AND4_X1 _11001_ ( .A1(\IF_ID_inst [22] ), .A2(_03318_ ), .A3(_03066_ ), .A4(_03322_ ), .ZN(_00225_ ) );
AND2_X1 _11002_ ( .A1(_03318_ ), .A2(_03322_ ), .ZN(_03325_ ) );
AOI221_X4 _11003_ ( .A(_03223_ ), .B1(\IF_ID_inst [23] ), .B2(_03325_ ), .C1(_03274_ ), .C2(_03297_ ), .ZN(_03326_ ) );
INV_X1 _11004_ ( .A(\ID_EX_rs2 [3] ), .ZN(_03327_ ) );
AOI211_X1 _11005_ ( .A(_03067_ ), .B(_03326_ ), .C1(_03301_ ), .C2(_03327_ ), .ZN(_00226_ ) );
AND4_X1 _11006_ ( .A1(\IF_ID_inst [21] ), .A2(_03318_ ), .A3(_03066_ ), .A4(_03322_ ), .ZN(_00227_ ) );
NAND4_X1 _11007_ ( .A1(_03303_ ), .A2(\IF_ID_inst [22] ), .A3(_03222_ ), .A4(_03325_ ), .ZN(_03328_ ) );
OAI21_X1 _11008_ ( .A(\ID_EX_rs2 [2] ), .B1(_03300_ ), .B2(_03224_ ), .ZN(_03329_ ) );
AOI21_X1 _11009_ ( .A(_03071_ ), .B1(_03328_ ), .B2(_03329_ ), .ZN(_00228_ ) );
AND4_X1 _11010_ ( .A1(\IF_ID_inst [20] ), .A2(_03318_ ), .A3(_03066_ ), .A4(_03322_ ), .ZN(_00229_ ) );
AOI221_X4 _11011_ ( .A(_03223_ ), .B1(\IF_ID_inst [21] ), .B2(_03325_ ), .C1(_03274_ ), .C2(_03297_ ), .ZN(_03330_ ) );
INV_X1 _11012_ ( .A(\ID_EX_rs2 [1] ), .ZN(_03331_ ) );
AOI211_X1 _11013_ ( .A(_03067_ ), .B(_03330_ ), .C1(_03301_ ), .C2(_03331_ ), .ZN(_00230_ ) );
NOR4_X1 _11014_ ( .A1(_03085_ ), .A2(_03079_ ), .A3(IDU_valid_EXU ), .A4(_03089_ ), .ZN(_00231_ ) );
NAND4_X1 _11015_ ( .A1(_03303_ ), .A2(\IF_ID_inst [20] ), .A3(_03222_ ), .A4(_03325_ ), .ZN(_03332_ ) );
OAI21_X1 _11016_ ( .A(\ID_EX_rs2 [0] ), .B1(_03300_ ), .B2(_03224_ ), .ZN(_03333_ ) );
AOI21_X1 _11017_ ( .A(_03071_ ), .B1(_03332_ ), .B2(_03333_ ), .ZN(_00232_ ) );
INV_X1 _11018_ ( .A(_03249_ ), .ZN(_03334_ ) );
OAI21_X1 _11019_ ( .A(_03257_ ), .B1(_03233_ ), .B2(_03117_ ), .ZN(_03335_ ) );
NAND4_X1 _11020_ ( .A1(_03334_ ), .A2(_03229_ ), .A3(_03271_ ), .A4(_03335_ ), .ZN(_03336_ ) );
NOR2_X1 _11021_ ( .A1(_03336_ ), .A2(_03254_ ), .ZN(_03337_ ) );
BUF_X2 _11022_ ( .A(_03337_ ), .Z(_03338_ ) );
NOR2_X1 _11023_ ( .A1(_03316_ ), .A2(_03090_ ), .ZN(_03339_ ) );
XNOR2_X1 _11024_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [20] ), .ZN(_03340_ ) );
INV_X1 _11025_ ( .A(\ID_EX_typ [7] ), .ZN(_03341_ ) );
AND2_X1 _11026_ ( .A1(\ID_EX_typ [6] ), .A2(\ID_EX_typ [5] ), .ZN(_03342_ ) );
AND3_X1 _11027_ ( .A1(_03340_ ), .A2(_03341_ ), .A3(_03342_ ), .ZN(_03343_ ) );
XNOR2_X1 _11028_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [22] ), .ZN(_03344_ ) );
XNOR2_X1 _11029_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [23] ), .ZN(_03345_ ) );
AND3_X1 _11030_ ( .A1(_03343_ ), .A2(_03344_ ), .A3(_03345_ ), .ZN(_03346_ ) );
XNOR2_X1 _11031_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [24] ), .ZN(_03347_ ) );
XNOR2_X1 _11032_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [21] ), .ZN(_03348_ ) );
NAND3_X1 _11033_ ( .A1(_03346_ ), .A2(_03347_ ), .A3(_03348_ ), .ZN(_03349_ ) );
AOI22_X1 _11034_ ( .A1(\ID_EX_rd [3] ), .A2(_03171_ ), .B1(_03302_ ), .B2(\ID_EX_rd [1] ), .ZN(_03350_ ) );
OR2_X1 _11035_ ( .A1(_03302_ ), .A2(\ID_EX_rd [1] ), .ZN(_03351_ ) );
OAI211_X1 _11036_ ( .A(_03350_ ), .B(_03351_ ), .C1(\ID_EX_rd [3] ), .C2(_03171_ ), .ZN(_03352_ ) );
XNOR2_X1 _11037_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [19] ), .ZN(_03353_ ) );
CLKBUF_X2 _11038_ ( .A(_03342_ ), .Z(_03354_ ) );
NAND3_X1 _11039_ ( .A1(_03353_ ), .A2(_03341_ ), .A3(_03354_ ), .ZN(_03355_ ) );
NOR2_X1 _11040_ ( .A1(_03352_ ), .A2(_03355_ ), .ZN(_03356_ ) );
XNOR2_X1 _11041_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [17] ), .ZN(_03357_ ) );
XNOR2_X1 _11042_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [15] ), .ZN(_03358_ ) );
NAND3_X1 _11043_ ( .A1(_03356_ ), .A2(_03357_ ), .A3(_03358_ ), .ZN(_03359_ ) );
NAND2_X1 _11044_ ( .A1(_03349_ ), .A2(_03359_ ), .ZN(_03360_ ) );
NAND4_X1 _11045_ ( .A1(_03339_ ), .A2(_03313_ ), .A3(_03168_ ), .A4(_03360_ ), .ZN(_03361_ ) );
AND3_X1 _11046_ ( .A1(_03338_ ), .A2(_03062_ ), .A3(_03361_ ), .ZN(_03362_ ) );
AND3_X1 _11047_ ( .A1(_03356_ ), .A2(_03357_ ), .A3(_03358_ ), .ZN(_03363_ ) );
AOI21_X1 _11048_ ( .A(_03363_ ), .B1(_03338_ ), .B2(_03062_ ), .ZN(_03364_ ) );
INV_X1 _11049_ ( .A(IDU_ready_IFU ), .ZN(_03365_ ) );
NOR4_X1 _11050_ ( .A1(_03362_ ), .A2(_03364_ ), .A3(_03365_ ), .A4(_03067_ ), .ZN(_00233_ ) );
AND4_X1 _11051_ ( .A1(_03070_ ), .A2(_03102_ ), .A3(_03073_ ), .A4(_03111_ ), .ZN(_03366_ ) );
NAND2_X1 _11052_ ( .A1(_03366_ ), .A2(_03106_ ), .ZN(_03367_ ) );
AND4_X1 _11053_ ( .A1(_03062_ ), .A2(_03367_ ), .A3(_03339_ ), .A4(_03309_ ), .ZN(_03368_ ) );
NOR2_X1 _11054_ ( .A1(_03130_ ), .A2(_03135_ ), .ZN(_03369_ ) );
NOR2_X1 _11055_ ( .A1(_03369_ ), .A2(_03118_ ), .ZN(_03370_ ) );
INV_X1 _11056_ ( .A(_03370_ ), .ZN(_03371_ ) );
AOI21_X1 _11057_ ( .A(_03071_ ), .B1(_03368_ ), .B2(_03371_ ), .ZN(_00234_ ) );
INV_X1 _11058_ ( .A(_03312_ ), .ZN(_03372_ ) );
NAND3_X1 _11059_ ( .A1(_03106_ ), .A2(_03070_ ), .A3(_03073_ ), .ZN(_03373_ ) );
NOR2_X1 _11060_ ( .A1(_03372_ ), .A2(_03373_ ), .ZN(_03374_ ) );
NOR2_X1 _11061_ ( .A1(_03374_ ), .A2(_03072_ ), .ZN(_03375_ ) );
AND2_X1 _11062_ ( .A1(_03228_ ), .A2(_03265_ ), .ZN(_03376_ ) );
INV_X1 _11063_ ( .A(_03376_ ), .ZN(_03377_ ) );
NAND2_X1 _11064_ ( .A1(_03228_ ), .A2(_03122_ ), .ZN(_03378_ ) );
AND4_X1 _11065_ ( .A1(_03262_ ), .A2(_03377_ ), .A3(_03378_ ), .A4(_03335_ ), .ZN(_03379_ ) );
AOI21_X1 _11066_ ( .A(_03071_ ), .B1(_03375_ ), .B2(_03379_ ), .ZN(_00235_ ) );
NOR3_X1 _11067_ ( .A1(_03276_ ), .A2(_03280_ ), .A3(_03283_ ), .ZN(_03380_ ) );
NAND4_X1 _11068_ ( .A1(_03226_ ), .A2(_03056_ ), .A3(_03237_ ), .A4(_03268_ ), .ZN(_03381_ ) );
AND3_X1 _11069_ ( .A1(_03296_ ), .A2(_03380_ ), .A3(_03381_ ), .ZN(_03382_ ) );
NOR2_X1 _11070_ ( .A1(_03374_ ), .A2(_03314_ ), .ZN(_03383_ ) );
AND3_X1 _11071_ ( .A1(_03236_ ), .A2(_03241_ ), .A3(_03287_ ), .ZN(_03384_ ) );
AND4_X1 _11072_ ( .A1(_03382_ ), .A2(_03383_ ), .A3(_03310_ ), .A4(_03384_ ), .ZN(_03385_ ) );
AOI21_X1 _11073_ ( .A(_03068_ ), .B1(_03385_ ), .B2(_03322_ ), .ZN(_00236_ ) );
AOI211_X1 _11074_ ( .A(_03090_ ), .B(_03247_ ), .C1(_03244_ ), .C2(_03250_ ), .ZN(_03386_ ) );
AOI21_X1 _11075_ ( .A(_03068_ ), .B1(_03322_ ), .B2(_03386_ ), .ZN(_00237_ ) );
NAND2_X1 _11076_ ( .A1(_03236_ ), .A2(_03241_ ), .ZN(_03387_ ) );
NOR3_X1 _11077_ ( .A1(_03316_ ), .A2(_03387_ ), .A3(_03119_ ), .ZN(_03388_ ) );
AOI21_X1 _11078_ ( .A(_03068_ ), .B1(_03388_ ), .B2(_03320_ ), .ZN(_00238_ ) );
AND3_X1 _11079_ ( .A1(_03056_ ), .A2(_03050_ ), .A3(_03051_ ), .ZN(_03389_ ) );
AND2_X1 _11080_ ( .A1(_03389_ ), .A2(_03121_ ), .ZN(_03390_ ) );
OR2_X1 _11081_ ( .A1(_03235_ ), .A2(_03290_ ), .ZN(_03391_ ) );
OAI21_X1 _11082_ ( .A(_03390_ ), .B1(_03391_ ), .B2(_03293_ ), .ZN(_03392_ ) );
AND2_X1 _11083_ ( .A1(_03285_ ), .A2(_03390_ ), .ZN(_03393_ ) );
INV_X1 _11084_ ( .A(_03393_ ), .ZN(_03394_ ) );
NAND2_X1 _11085_ ( .A1(_03392_ ), .A2(_03394_ ), .ZN(_03395_ ) );
AND3_X1 _11086_ ( .A1(_03252_ ), .A2(_03118_ ), .A3(_03121_ ), .ZN(_03396_ ) );
NOR4_X1 _11087_ ( .A1(_03395_ ), .A2(_03167_ ), .A3(_03258_ ), .A4(_03396_ ), .ZN(_03397_ ) );
AND2_X1 _11088_ ( .A1(_03252_ ), .A2(_03121_ ), .ZN(_03398_ ) );
NAND2_X1 _11089_ ( .A1(_03398_ ), .A2(_03285_ ), .ZN(_03399_ ) );
NAND3_X1 _11090_ ( .A1(_03293_ ), .A2(_03121_ ), .A3(_03252_ ), .ZN(_03400_ ) );
NAND4_X1 _11091_ ( .A1(_03252_ ), .A2(_03289_ ), .A3(_03121_ ), .A4(_03231_ ), .ZN(_03401_ ) );
NAND3_X1 _11092_ ( .A1(_03399_ ), .A2(_03400_ ), .A3(_03401_ ), .ZN(_03402_ ) );
AND2_X1 _11093_ ( .A1(_03130_ ), .A2(\IF_ID_inst [14] ), .ZN(_03403_ ) );
AND3_X1 _11094_ ( .A1(_03053_ ), .A2(\IF_ID_inst [13] ), .A3(_03060_ ), .ZN(_03404_ ) );
NOR4_X1 _11095_ ( .A1(_03402_ ), .A2(_03403_ ), .A3(_03119_ ), .A4(_03404_ ), .ZN(_03405_ ) );
AOI21_X1 _11096_ ( .A(_03068_ ), .B1(_03397_ ), .B2(_03405_ ), .ZN(_00239_ ) );
NAND2_X1 _11097_ ( .A1(_03165_ ), .A2(_03282_ ), .ZN(_03406_ ) );
AOI221_X4 _11098_ ( .A(_03059_ ), .B1(_03116_ ), .B2(_03118_ ), .C1(\IF_ID_inst [14] ), .C2(_03135_ ), .ZN(_03407_ ) );
INV_X1 _11099_ ( .A(_03276_ ), .ZN(_03408_ ) );
OAI21_X1 _11100_ ( .A(_03122_ ), .B1(_03260_ ), .B2(_03228_ ), .ZN(_03409_ ) );
AND4_X1 _11101_ ( .A1(_03406_ ), .A2(_03407_ ), .A3(_03408_ ), .A4(_03409_ ), .ZN(_03410_ ) );
AND2_X1 _11102_ ( .A1(_03244_ ), .A2(\IF_ID_inst [14] ), .ZN(_03411_ ) );
INV_X1 _11103_ ( .A(_03411_ ), .ZN(_03412_ ) );
OAI22_X1 _11104_ ( .A1(_03275_ ), .A2(_03285_ ), .B1(_03264_ ), .B2(_03286_ ), .ZN(_03413_ ) );
NOR2_X1 _11105_ ( .A1(_03280_ ), .A2(_03376_ ), .ZN(_03414_ ) );
AND3_X1 _11106_ ( .A1(_03412_ ), .A2(_03413_ ), .A3(_03414_ ), .ZN(_03415_ ) );
AOI21_X1 _11107_ ( .A(_03068_ ), .B1(_03410_ ), .B2(_03415_ ), .ZN(_00240_ ) );
AND2_X1 _11108_ ( .A1(_03285_ ), .A2(_03286_ ), .ZN(_03416_ ) );
AOI211_X1 _11109_ ( .A(_03119_ ), .B(_03416_ ), .C1(_03312_ ), .C2(_03107_ ), .ZN(_03417_ ) );
AND4_X1 _11110_ ( .A1(_03281_ ), .A2(_03268_ ), .A3(_03282_ ), .A4(_03237_ ), .ZN(_03418_ ) );
AND3_X1 _11111_ ( .A1(_03264_ ), .A2(_03237_ ), .A3(_03268_ ), .ZN(_03419_ ) );
AOI211_X1 _11112_ ( .A(_03418_ ), .B(_03419_ ), .C1(_03122_ ), .C2(_03130_ ), .ZN(_03420_ ) );
AND4_X1 _11113_ ( .A1(_03261_ ), .A2(_03417_ ), .A3(_03408_ ), .A4(_03420_ ), .ZN(_03421_ ) );
OAI211_X1 _11114_ ( .A(\IF_ID_inst [14] ), .B(_03117_ ), .C1(_03244_ ), .C2(_03061_ ), .ZN(_03422_ ) );
AND4_X1 _11115_ ( .A1(_03132_ ), .A2(_03421_ ), .A3(_03271_ ), .A4(_03422_ ), .ZN(_03423_ ) );
OAI21_X1 _11116_ ( .A(_03131_ ), .B1(_03135_ ), .B2(_03061_ ), .ZN(_03424_ ) );
NOR3_X1 _11117_ ( .A1(_03054_ ), .A2(_03233_ ), .A3(_03058_ ), .ZN(_03425_ ) );
AOI221_X4 _11118_ ( .A(_03425_ ), .B1(_03285_ ), .B2(_03264_ ), .C1(_03257_ ), .C2(_03265_ ), .ZN(_03426_ ) );
AND2_X1 _11119_ ( .A1(_03226_ ), .A2(_03056_ ), .ZN(_03427_ ) );
AOI22_X1 _11120_ ( .A1(_03427_ ), .A2(_03235_ ), .B1(_03286_ ), .B2(_03279_ ), .ZN(_03428_ ) );
AOI22_X1 _11121_ ( .A1(\IF_ID_inst [14] ), .A2(_03247_ ), .B1(_03228_ ), .B2(_03265_ ), .ZN(_03429_ ) );
AND4_X1 _11122_ ( .A1(_03424_ ), .A2(_03426_ ), .A3(_03428_ ), .A4(_03429_ ), .ZN(_03430_ ) );
AOI21_X1 _11123_ ( .A(_03068_ ), .B1(_03423_ ), .B2(_03430_ ), .ZN(_00241_ ) );
INV_X1 _11124_ ( .A(_03215_ ), .ZN(_03431_ ) );
INV_X2 _11125_ ( .A(fanout_net_41 ), .ZN(_03432_ ) );
BUF_X4 _11126_ ( .A(_03432_ ), .Z(_03433_ ) );
NAND4_X1 _11127_ ( .A1(_03431_ ), .A2(check_quest ), .A3(\myexu.pc_jump [0] ), .A4(_03433_ ), .ZN(_03434_ ) );
NAND2_X1 _11128_ ( .A1(\mtvec [0] ), .A2(fanout_net_41 ), .ZN(_03435_ ) );
AOI21_X1 _11129_ ( .A(fanout_net_2 ), .B1(_03434_ ), .B2(_03435_ ), .ZN(_00245_ ) );
INV_X1 _11130_ ( .A(_03217_ ), .ZN(_03436_ ) );
BUF_X4 _11131_ ( .A(_03436_ ), .Z(_03437_ ) );
AND4_X1 _11132_ ( .A1(\IF_ID_inst [31] ), .A2(_03128_ ), .A3(_03159_ ), .A4(\IF_ID_inst [5] ), .ZN(_03438_ ) );
AND2_X2 _11133_ ( .A1(_03052_ ), .A2(_03438_ ), .ZN(_03439_ ) );
AOI21_X1 _11134_ ( .A(_03439_ ), .B1(_03163_ ), .B2(\IF_ID_inst [31] ), .ZN(_03440_ ) );
AND2_X1 _11135_ ( .A1(_03439_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03441_ ) );
NOR2_X1 _11136_ ( .A1(_03440_ ), .A2(_03441_ ), .ZN(_03442_ ) );
BUF_X4 _11137_ ( .A(_03442_ ), .Z(_03443_ ) );
BUF_X4 _11138_ ( .A(_03443_ ), .Z(_03444_ ) );
XNOR2_X1 _11139_ ( .A(_03444_ ), .B(_01841_ ), .ZN(_03445_ ) );
INV_X1 _11140_ ( .A(_03445_ ), .ZN(_03446_ ) );
AND2_X1 _11141_ ( .A1(_03163_ ), .A2(\IF_ID_inst [19] ), .ZN(_03447_ ) );
INV_X1 _11142_ ( .A(_03439_ ), .ZN(_03448_ ) );
MUX2_X1 _11143_ ( .A(_03267_ ), .B(_03447_ ), .S(_03448_ ), .Z(_03449_ ) );
XOR2_X1 _11144_ ( .A(_03449_ ), .B(\IF_ID_pc [19] ), .Z(_03450_ ) );
XNOR2_X1 _11145_ ( .A(_03442_ ), .B(_01971_ ), .ZN(_03451_ ) );
AND2_X1 _11146_ ( .A1(_03450_ ), .A2(_03451_ ), .ZN(_03452_ ) );
AND2_X1 _11147_ ( .A1(_03163_ ), .A2(\IF_ID_inst [18] ), .ZN(_03453_ ) );
NAND4_X1 _11148_ ( .A1(_03114_ ), .A2(_03159_ ), .A3(_03050_ ), .A4(_03051_ ), .ZN(_03454_ ) );
NOR2_X1 _11149_ ( .A1(_03454_ ), .A2(_03064_ ), .ZN(_03455_ ) );
INV_X1 _11150_ ( .A(_03455_ ), .ZN(_03456_ ) );
MUX2_X1 _11151_ ( .A(_03267_ ), .B(_03453_ ), .S(_03456_ ), .Z(_03457_ ) );
XNOR2_X1 _11152_ ( .A(_03457_ ), .B(_01975_ ), .ZN(_03458_ ) );
AND2_X1 _11153_ ( .A1(_03163_ ), .A2(\IF_ID_inst [17] ), .ZN(_03459_ ) );
MUX2_X1 _11154_ ( .A(_03267_ ), .B(_03459_ ), .S(_03448_ ), .Z(_03460_ ) );
XNOR2_X1 _11155_ ( .A(_03460_ ), .B(_01981_ ), .ZN(_03461_ ) );
AND2_X1 _11156_ ( .A1(_03458_ ), .A2(_03461_ ), .ZN(_03462_ ) );
INV_X1 _11157_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03463_ ) );
NOR3_X1 _11158_ ( .A1(_03454_ ), .A2(_03064_ ), .A3(_03463_ ), .ZN(_03464_ ) );
AOI21_X1 _11159_ ( .A(_03464_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .B2(_03161_ ), .ZN(_03465_ ) );
XOR2_X1 _11160_ ( .A(_03465_ ), .B(\IF_ID_pc [2] ), .Z(_03466_ ) );
INV_X1 _11161_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03467_ ) );
AND3_X1 _11162_ ( .A1(_03052_ ), .A2(_03438_ ), .A3(_03467_ ), .ZN(_03468_ ) );
AOI21_X1 _11163_ ( .A(_03468_ ), .B1(\IF_ID_inst [21] ), .B2(_03161_ ), .ZN(_03469_ ) );
INV_X1 _11164_ ( .A(\IF_ID_pc [1] ), .ZN(_03470_ ) );
NOR2_X1 _11165_ ( .A1(_03469_ ), .A2(_03470_ ), .ZN(_03471_ ) );
AND2_X1 _11166_ ( .A1(_03466_ ), .A2(_03471_ ), .ZN(_03472_ ) );
AND2_X1 _11167_ ( .A1(_03465_ ), .A2(\IF_ID_pc [2] ), .ZN(_03473_ ) );
NOR2_X1 _11168_ ( .A1(_03472_ ), .A2(_03473_ ), .ZN(_03474_ ) );
AOI21_X1 _11169_ ( .A(_03455_ ), .B1(_03161_ ), .B2(\IF_ID_inst [23] ), .ZN(_03475_ ) );
INV_X1 _11170_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03476_ ) );
NOR3_X1 _11171_ ( .A1(_03454_ ), .A2(_03064_ ), .A3(_03476_ ), .ZN(_03477_ ) );
NOR2_X1 _11172_ ( .A1(_03475_ ), .A2(_03477_ ), .ZN(_03478_ ) );
XNOR2_X1 _11173_ ( .A(_03478_ ), .B(fanout_net_7 ), .ZN(_03479_ ) );
OR2_X1 _11174_ ( .A1(_03474_ ), .A2(_03479_ ), .ZN(_03480_ ) );
OR3_X1 _11175_ ( .A1(_03475_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .A3(_03477_ ), .ZN(_03481_ ) );
NAND2_X1 _11176_ ( .A1(_03480_ ), .A2(_03481_ ), .ZN(_03482_ ) );
INV_X1 _11177_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03483_ ) );
NAND3_X1 _11178_ ( .A1(_03052_ ), .A2(_03438_ ), .A3(_03483_ ), .ZN(_03484_ ) );
INV_X1 _11179_ ( .A(_03163_ ), .ZN(_03485_ ) );
OAI21_X1 _11180_ ( .A(_03484_ ), .B1(_03485_ ), .B2(_03080_ ), .ZN(_03486_ ) );
OAI21_X1 _11181_ ( .A(_03482_ ), .B1(fanout_net_11 ), .B2(_03486_ ), .ZN(_03487_ ) );
NAND2_X1 _11182_ ( .A1(_03486_ ), .A2(fanout_net_11 ), .ZN(_03488_ ) );
AND2_X1 _11183_ ( .A1(_03487_ ), .A2(_03488_ ), .ZN(_03489_ ) );
NOR2_X1 _11184_ ( .A1(_03448_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03490_ ) );
AND2_X1 _11185_ ( .A1(_03162_ ), .A2(\IF_ID_inst [25] ), .ZN(_03491_ ) );
NOR2_X1 _11186_ ( .A1(_03490_ ), .A2(_03491_ ), .ZN(_03492_ ) );
INV_X1 _11187_ ( .A(\IF_ID_pc [5] ), .ZN(_03493_ ) );
XNOR2_X1 _11188_ ( .A(_03492_ ), .B(_03493_ ), .ZN(_03494_ ) );
AND2_X1 _11189_ ( .A1(_03162_ ), .A2(\IF_ID_inst [26] ), .ZN(_03495_ ) );
INV_X1 _11190_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03496_ ) );
AOI21_X1 _11191_ ( .A(_03495_ ), .B1(_03496_ ), .B2(_03439_ ), .ZN(_03497_ ) );
XNOR2_X1 _11192_ ( .A(_03497_ ), .B(\IF_ID_pc [6] ), .ZN(_03498_ ) );
INV_X1 _11193_ ( .A(_03498_ ), .ZN(_03499_ ) );
AND2_X1 _11194_ ( .A1(_03161_ ), .A2(\IF_ID_inst [28] ), .ZN(_03500_ ) );
INV_X1 _11195_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03501_ ) );
AOI21_X1 _11196_ ( .A(_03500_ ), .B1(_03501_ ), .B2(_03439_ ), .ZN(_03502_ ) );
XNOR2_X1 _11197_ ( .A(_03502_ ), .B(\IF_ID_pc [8] ), .ZN(_03503_ ) );
NAND2_X1 _11198_ ( .A1(_03162_ ), .A2(\IF_ID_inst [27] ), .ZN(_03504_ ) );
OAI21_X1 _11199_ ( .A(_03504_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_03448_ ), .ZN(_03505_ ) );
XOR2_X1 _11200_ ( .A(_03505_ ), .B(\IF_ID_pc [7] ), .Z(_03506_ ) );
NAND2_X1 _11201_ ( .A1(_03503_ ), .A2(_03506_ ), .ZN(_03507_ ) );
NOR4_X1 _11202_ ( .A1(_03489_ ), .A2(_03494_ ), .A3(_03499_ ), .A4(_03507_ ), .ZN(_03508_ ) );
NAND3_X1 _11203_ ( .A1(_03503_ ), .A2(\IF_ID_pc [7] ), .A3(_03505_ ), .ZN(_03509_ ) );
NOR2_X1 _11204_ ( .A1(_03497_ ), .A2(_01824_ ), .ZN(_03510_ ) );
AND2_X1 _11205_ ( .A1(_03497_ ), .A2(_01824_ ), .ZN(_03511_ ) );
INV_X1 _11206_ ( .A(_03511_ ), .ZN(_03512_ ) );
NOR2_X1 _11207_ ( .A1(_03492_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03513_ ) );
AOI21_X1 _11208_ ( .A(_03510_ ), .B1(_03512_ ), .B2(_03513_ ), .ZN(_03514_ ) );
OAI221_X1 _11209_ ( .A(_03509_ ), .B1(_01886_ ), .B2(_03502_ ), .C1(_03514_ ), .C2(_03507_ ), .ZN(_03515_ ) );
OR2_X1 _11210_ ( .A1(_03508_ ), .A2(_03515_ ), .ZN(_03516_ ) );
AND2_X1 _11211_ ( .A1(_03455_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03517_ ) );
INV_X1 _11212_ ( .A(_03517_ ), .ZN(_03518_ ) );
AND2_X1 _11213_ ( .A1(_03163_ ), .A2(\IF_ID_inst [16] ), .ZN(_03519_ ) );
OAI21_X1 _11214_ ( .A(_03518_ ), .B1(_03519_ ), .B2(_03455_ ), .ZN(_03520_ ) );
XNOR2_X1 _11215_ ( .A(_03520_ ), .B(_01851_ ), .ZN(_03521_ ) );
AND2_X1 _11216_ ( .A1(_03162_ ), .A2(\IF_ID_inst [15] ), .ZN(_03522_ ) );
MUX2_X1 _11217_ ( .A(_03267_ ), .B(_03522_ ), .S(_03448_ ), .Z(_03523_ ) );
AND2_X1 _11218_ ( .A1(_03523_ ), .A2(\IF_ID_pc [15] ), .ZN(_03524_ ) );
NOR2_X1 _11219_ ( .A1(_03523_ ), .A2(\IF_ID_pc [15] ), .ZN(_03525_ ) );
NOR3_X1 _11220_ ( .A1(_03521_ ), .A2(_03524_ ), .A3(_03525_ ), .ZN(_03526_ ) );
AND2_X1 _11221_ ( .A1(_03162_ ), .A2(\IF_ID_inst [13] ), .ZN(_03527_ ) );
MUX2_X1 _11222_ ( .A(_03267_ ), .B(_03527_ ), .S(_03448_ ), .Z(_03528_ ) );
XOR2_X1 _11223_ ( .A(_03528_ ), .B(\IF_ID_pc [13] ), .Z(_03529_ ) );
AND2_X1 _11224_ ( .A1(_03162_ ), .A2(\IF_ID_inst [14] ), .ZN(_03530_ ) );
MUX2_X1 _11225_ ( .A(_03267_ ), .B(_03530_ ), .S(_03448_ ), .Z(_03531_ ) );
XOR2_X1 _11226_ ( .A(_03531_ ), .B(\IF_ID_pc [14] ), .Z(_03532_ ) );
AND2_X1 _11227_ ( .A1(_03529_ ), .A2(_03532_ ), .ZN(_03533_ ) );
NAND2_X1 _11228_ ( .A1(_03162_ ), .A2(\IF_ID_inst [20] ), .ZN(_03534_ ) );
OAI21_X1 _11229_ ( .A(_03534_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_03448_ ), .ZN(_03535_ ) );
XNOR2_X1 _11230_ ( .A(_03535_ ), .B(_01784_ ), .ZN(_03536_ ) );
AOI21_X1 _11231_ ( .A(_03439_ ), .B1(_03163_ ), .B2(\IF_ID_inst [12] ), .ZN(_03537_ ) );
NOR3_X1 _11232_ ( .A1(_03537_ ), .A2(_03517_ ), .A3(_01893_ ), .ZN(_03538_ ) );
INV_X1 _11233_ ( .A(_03538_ ), .ZN(_03539_ ) );
OAI21_X1 _11234_ ( .A(_01893_ ), .B1(_03537_ ), .B2(_03441_ ), .ZN(_03540_ ) );
AND3_X1 _11235_ ( .A1(_03536_ ), .A2(_03539_ ), .A3(_03540_ ), .ZN(_03541_ ) );
AND2_X1 _11236_ ( .A1(_03162_ ), .A2(\IF_ID_inst [29] ), .ZN(_03542_ ) );
INV_X1 _11237_ ( .A(_03542_ ), .ZN(_03543_ ) );
INV_X1 _11238_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03544_ ) );
NAND4_X1 _11239_ ( .A1(_03160_ ), .A2(\IF_ID_inst [31] ), .A3(_03052_ ), .A4(_03544_ ), .ZN(_03545_ ) );
AND3_X1 _11240_ ( .A1(_03543_ ), .A2(_01913_ ), .A3(_03545_ ), .ZN(_03546_ ) );
AOI21_X1 _11241_ ( .A(_01913_ ), .B1(_03543_ ), .B2(_03545_ ), .ZN(_03547_ ) );
NOR2_X1 _11242_ ( .A1(_03546_ ), .A2(_03547_ ), .ZN(_03548_ ) );
AND2_X1 _11243_ ( .A1(_03162_ ), .A2(\IF_ID_inst [30] ), .ZN(_03549_ ) );
INV_X1 _11244_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03550_ ) );
AOI21_X1 _11245_ ( .A(_03549_ ), .B1(_03550_ ), .B2(_03439_ ), .ZN(_03551_ ) );
OR2_X1 _11246_ ( .A1(_03551_ ), .A2(_01900_ ), .ZN(_03552_ ) );
NAND2_X1 _11247_ ( .A1(_03551_ ), .A2(_01900_ ), .ZN(_03553_ ) );
AND3_X1 _11248_ ( .A1(_03548_ ), .A2(_03552_ ), .A3(_03553_ ), .ZN(_03554_ ) );
AND4_X1 _11249_ ( .A1(_03526_ ), .A2(_03533_ ), .A3(_03541_ ), .A4(_03554_ ), .ZN(_03555_ ) );
AND2_X1 _11250_ ( .A1(_03516_ ), .A2(_03555_ ), .ZN(_03556_ ) );
AND3_X1 _11251_ ( .A1(_03552_ ), .A2(_03553_ ), .A3(_03547_ ), .ZN(_03557_ ) );
NOR2_X1 _11252_ ( .A1(_03551_ ), .A2(_01900_ ), .ZN(_03558_ ) );
OAI21_X1 _11253_ ( .A(_03541_ ), .B1(_03557_ ), .B2(_03558_ ), .ZN(_03559_ ) );
NAND4_X1 _11254_ ( .A1(_03539_ ), .A2(\IF_ID_pc [11] ), .A3(_03540_ ), .A4(_03535_ ), .ZN(_03560_ ) );
NAND3_X1 _11255_ ( .A1(_03559_ ), .A2(_03539_ ), .A3(_03560_ ), .ZN(_03561_ ) );
NAND3_X1 _11256_ ( .A1(_03561_ ), .A2(_03526_ ), .A3(_03533_ ), .ZN(_03562_ ) );
OR2_X1 _11257_ ( .A1(_03520_ ), .A2(_01851_ ), .ZN(_03563_ ) );
NOR2_X1 _11258_ ( .A1(_03531_ ), .A2(\IF_ID_pc [14] ), .ZN(_03564_ ) );
AND2_X1 _11259_ ( .A1(_03528_ ), .A2(\IF_ID_pc [13] ), .ZN(_03565_ ) );
INV_X1 _11260_ ( .A(_03565_ ), .ZN(_03566_ ) );
NAND2_X1 _11261_ ( .A1(_03531_ ), .A2(\IF_ID_pc [14] ), .ZN(_03567_ ) );
AOI21_X1 _11262_ ( .A(_03564_ ), .B1(_03566_ ), .B2(_03567_ ), .ZN(_03568_ ) );
NAND2_X1 _11263_ ( .A1(_03568_ ), .A2(_03526_ ), .ZN(_03569_ ) );
INV_X1 _11264_ ( .A(_03524_ ), .ZN(_03570_ ) );
OR2_X1 _11265_ ( .A1(_03570_ ), .A2(_03521_ ), .ZN(_03571_ ) );
NAND4_X1 _11266_ ( .A1(_03562_ ), .A2(_03563_ ), .A3(_03569_ ), .A4(_03571_ ), .ZN(_03572_ ) );
OAI211_X1 _11267_ ( .A(_03452_ ), .B(_03462_ ), .C1(_03556_ ), .C2(_03572_ ), .ZN(_03573_ ) );
OAI211_X1 _11268_ ( .A(_03449_ ), .B(\IF_ID_pc [19] ), .C1(\IF_ID_pc [20] ), .C2(_03442_ ), .ZN(_03574_ ) );
INV_X1 _11269_ ( .A(_03442_ ), .ZN(_03575_ ) );
OAI21_X1 _11270_ ( .A(_03574_ ), .B1(_01971_ ), .B2(_03575_ ), .ZN(_03576_ ) );
AND2_X1 _11271_ ( .A1(_03457_ ), .A2(\IF_ID_pc [18] ), .ZN(_03577_ ) );
AND2_X1 _11272_ ( .A1(_03460_ ), .A2(\IF_ID_pc [17] ), .ZN(_03578_ ) );
AOI21_X1 _11273_ ( .A(_03577_ ), .B1(_03458_ ), .B2(_03578_ ), .ZN(_03579_ ) );
INV_X1 _11274_ ( .A(_03579_ ), .ZN(_03580_ ) );
AOI21_X1 _11275_ ( .A(_03576_ ), .B1(_03580_ ), .B2(_03452_ ), .ZN(_03581_ ) );
AND2_X1 _11276_ ( .A1(_03573_ ), .A2(_03581_ ), .ZN(_03582_ ) );
XNOR2_X1 _11277_ ( .A(_03442_ ), .B(_01817_ ), .ZN(_03583_ ) );
XNOR2_X1 _11278_ ( .A(_03442_ ), .B(_01915_ ), .ZN(_03584_ ) );
NAND2_X1 _11279_ ( .A1(_03583_ ), .A2(_03584_ ), .ZN(_03585_ ) );
XNOR2_X1 _11280_ ( .A(_03443_ ), .B(\IF_ID_pc [22] ), .ZN(_03586_ ) );
XNOR2_X1 _11281_ ( .A(_03443_ ), .B(_01843_ ), .ZN(_03587_ ) );
INV_X1 _11282_ ( .A(_03587_ ), .ZN(_03588_ ) );
NOR4_X1 _11283_ ( .A1(_03582_ ), .A2(_03585_ ), .A3(_03586_ ), .A4(_03588_ ), .ZN(_03589_ ) );
AND2_X1 _11284_ ( .A1(_03583_ ), .A2(_03584_ ), .ZN(_03590_ ) );
AND2_X1 _11285_ ( .A1(_03443_ ), .A2(\IF_ID_pc [22] ), .ZN(_03591_ ) );
AND2_X1 _11286_ ( .A1(_03443_ ), .A2(\IF_ID_pc [21] ), .ZN(_03592_ ) );
OAI21_X1 _11287_ ( .A(_03590_ ), .B1(_03591_ ), .B2(_03592_ ), .ZN(_03593_ ) );
NAND2_X1 _11288_ ( .A1(_03443_ ), .A2(\IF_ID_pc [24] ), .ZN(_03594_ ) );
NAND2_X1 _11289_ ( .A1(_03443_ ), .A2(\IF_ID_pc [23] ), .ZN(_03595_ ) );
NAND3_X1 _11290_ ( .A1(_03593_ ), .A2(_03594_ ), .A3(_03595_ ), .ZN(_03596_ ) );
OR2_X1 _11291_ ( .A1(_03589_ ), .A2(_03596_ ), .ZN(_03597_ ) );
XNOR2_X1 _11292_ ( .A(_03443_ ), .B(_02004_ ), .ZN(_03598_ ) );
XNOR2_X1 _11293_ ( .A(_03443_ ), .B(_01836_ ), .ZN(_03599_ ) );
AND3_X1 _11294_ ( .A1(_03597_ ), .A2(_03598_ ), .A3(_03599_ ), .ZN(_03600_ ) );
XNOR2_X1 _11295_ ( .A(_03444_ ), .B(_01777_ ), .ZN(_03601_ ) );
XNOR2_X1 _11296_ ( .A(_03443_ ), .B(_02001_ ), .ZN(_03602_ ) );
NAND3_X1 _11297_ ( .A1(_03600_ ), .A2(_03601_ ), .A3(_03602_ ), .ZN(_03603_ ) );
OAI21_X1 _11298_ ( .A(_03444_ ), .B1(\IF_ID_pc [26] ), .B2(\IF_ID_pc [25] ), .ZN(_03604_ ) );
INV_X1 _11299_ ( .A(_03604_ ), .ZN(_03605_ ) );
NAND3_X1 _11300_ ( .A1(_03601_ ), .A2(_03602_ ), .A3(_03605_ ), .ZN(_03606_ ) );
NAND2_X1 _11301_ ( .A1(_03444_ ), .A2(\IF_ID_pc [28] ), .ZN(_03607_ ) );
AND2_X1 _11302_ ( .A1(_03444_ ), .A2(\IF_ID_pc [27] ), .ZN(_03608_ ) );
INV_X1 _11303_ ( .A(_03608_ ), .ZN(_03609_ ) );
AND3_X1 _11304_ ( .A1(_03606_ ), .A2(_03607_ ), .A3(_03609_ ), .ZN(_03610_ ) );
AOI21_X1 _11305_ ( .A(_03446_ ), .B1(_03603_ ), .B2(_03610_ ), .ZN(_03611_ ) );
NOR3_X1 _11306_ ( .A1(_03440_ ), .A2(_03517_ ), .A3(_01841_ ), .ZN(_03612_ ) );
OR2_X1 _11307_ ( .A1(_03611_ ), .A2(_03612_ ), .ZN(_03613_ ) );
XNOR2_X1 _11308_ ( .A(_03444_ ), .B(_01770_ ), .ZN(_03614_ ) );
OAI21_X1 _11309_ ( .A(_03437_ ), .B1(_03613_ ), .B2(_03614_ ), .ZN(_03615_ ) );
AOI21_X1 _11310_ ( .A(_03615_ ), .B1(_03613_ ), .B2(_03614_ ), .ZN(_03616_ ) );
BUF_X2 _11311_ ( .A(_03217_ ), .Z(_03617_ ) );
BUF_X4 _11312_ ( .A(_03617_ ), .Z(_03618_ ) );
AOI211_X1 _11313_ ( .A(fanout_net_41 ), .B(_03616_ ), .C1(\myexu.pc_jump [30] ), .C2(_03618_ ), .ZN(_03619_ ) );
BUF_X4 _11314_ ( .A(_03432_ ), .Z(_03620_ ) );
NOR2_X1 _11315_ ( .A1(_03620_ ), .A2(\mtvec [30] ), .ZN(_03621_ ) );
NOR3_X1 _11316_ ( .A1(_03619_ ), .A2(fanout_net_2 ), .A3(_03621_ ), .ZN(_00246_ ) );
BUF_X4 _11317_ ( .A(_03437_ ), .Z(_03622_ ) );
AND3_X1 _11318_ ( .A1(_03573_ ), .A2(_03588_ ), .A3(_03581_ ), .ZN(_03623_ ) );
AOI21_X1 _11319_ ( .A(_03588_ ), .B1(_03573_ ), .B2(_03581_ ), .ZN(_03624_ ) );
OAI21_X1 _11320_ ( .A(_03622_ ), .B1(_03623_ ), .B2(_03624_ ), .ZN(_03625_ ) );
BUF_X4 _11321_ ( .A(_03432_ ), .Z(_03626_ ) );
BUF_X4 _11322_ ( .A(_03437_ ), .Z(_03627_ ) );
OAI211_X1 _11323_ ( .A(_03625_ ), .B(_03626_ ), .C1(\myexu.pc_jump [21] ), .C2(_03627_ ), .ZN(_03628_ ) );
NAND2_X1 _11324_ ( .A1(\mtvec [21] ), .A2(fanout_net_41 ), .ZN(_03629_ ) );
AOI21_X1 _11325_ ( .A(fanout_net_2 ), .B1(_03628_ ), .B2(_03629_ ), .ZN(_00247_ ) );
OAI21_X1 _11326_ ( .A(_03462_ ), .B1(_03556_ ), .B2(_03572_ ), .ZN(_03630_ ) );
NAND2_X1 _11327_ ( .A1(_03630_ ), .A2(_03579_ ), .ZN(_03631_ ) );
AND2_X1 _11328_ ( .A1(_03631_ ), .A2(_03450_ ), .ZN(_03632_ ) );
AOI21_X1 _11329_ ( .A(_03632_ ), .B1(\IF_ID_pc [19] ), .B2(_03449_ ), .ZN(_03633_ ) );
XNOR2_X1 _11330_ ( .A(_03633_ ), .B(_03451_ ), .ZN(_03634_ ) );
MUX2_X1 _11331_ ( .A(\myexu.pc_jump [20] ), .B(_03634_ ), .S(_03436_ ), .Z(_03635_ ) );
MUX2_X1 _11332_ ( .A(\mtvec [20] ), .B(_03635_ ), .S(_03432_ ), .Z(_03636_ ) );
AND2_X1 _11333_ ( .A1(_03636_ ), .A2(_01618_ ), .ZN(_00248_ ) );
OR3_X1 _11334_ ( .A1(_03215_ ), .A2(_03216_ ), .A3(\myexu.pc_jump [19] ), .ZN(_03637_ ) );
XOR2_X1 _11335_ ( .A(_03631_ ), .B(_03450_ ), .Z(_03638_ ) );
OAI211_X1 _11336_ ( .A(_03620_ ), .B(_03637_ ), .C1(_03638_ ), .C2(_03618_ ), .ZN(_03639_ ) );
NAND2_X1 _11337_ ( .A1(\mtvec [19] ), .A2(fanout_net_41 ), .ZN(_03640_ ) );
AOI21_X1 _11338_ ( .A(fanout_net_2 ), .B1(_03639_ ), .B2(_03640_ ), .ZN(_00249_ ) );
OAI21_X1 _11339_ ( .A(_03461_ ), .B1(_03556_ ), .B2(_03572_ ), .ZN(_03641_ ) );
INV_X1 _11340_ ( .A(_03578_ ), .ZN(_03642_ ) );
AND3_X1 _11341_ ( .A1(_03641_ ), .A2(_03642_ ), .A3(_03458_ ), .ZN(_03643_ ) );
AOI21_X1 _11342_ ( .A(_03458_ ), .B1(_03641_ ), .B2(_03642_ ), .ZN(_03644_ ) );
OR3_X1 _11343_ ( .A1(_03643_ ), .A2(_03644_ ), .A3(_03617_ ), .ZN(_03645_ ) );
OAI211_X1 _11344_ ( .A(_03645_ ), .B(_03626_ ), .C1(\myexu.pc_jump [18] ), .C2(_03627_ ), .ZN(_03646_ ) );
NAND2_X1 _11345_ ( .A1(\mtvec [18] ), .A2(fanout_net_41 ), .ZN(_03647_ ) );
AOI21_X1 _11346_ ( .A(fanout_net_2 ), .B1(_03646_ ), .B2(_03647_ ), .ZN(_00250_ ) );
NOR2_X1 _11347_ ( .A1(_03556_ ), .A2(_03572_ ), .ZN(_03648_ ) );
XOR2_X1 _11348_ ( .A(_03648_ ), .B(_03461_ ), .Z(_03649_ ) );
NAND2_X1 _11349_ ( .A1(_03649_ ), .A2(_03622_ ), .ZN(_03650_ ) );
OAI211_X1 _11350_ ( .A(_03650_ ), .B(_03626_ ), .C1(\myexu.pc_jump [17] ), .C2(_03627_ ), .ZN(_03651_ ) );
NAND2_X1 _11351_ ( .A1(\mtvec [17] ), .A2(fanout_net_41 ), .ZN(_03652_ ) );
AOI21_X1 _11352_ ( .A(fanout_net_2 ), .B1(_03651_ ), .B2(_03652_ ), .ZN(_00251_ ) );
INV_X1 _11353_ ( .A(\IF_ID_pc [15] ), .ZN(_03653_ ) );
XNOR2_X1 _11354_ ( .A(_03523_ ), .B(_03653_ ), .ZN(_03654_ ) );
OAI211_X1 _11355_ ( .A(_03541_ ), .B(_03554_ ), .C1(_03508_ ), .C2(_03515_ ), .ZN(_03655_ ) );
AND3_X1 _11356_ ( .A1(_03559_ ), .A2(_03539_ ), .A3(_03560_ ), .ZN(_03656_ ) );
NAND2_X1 _11357_ ( .A1(_03655_ ), .A2(_03656_ ), .ZN(_03657_ ) );
AND2_X1 _11358_ ( .A1(_03657_ ), .A2(_03533_ ), .ZN(_03658_ ) );
OAI21_X1 _11359_ ( .A(_03654_ ), .B1(_03658_ ), .B2(_03568_ ), .ZN(_03659_ ) );
AND3_X1 _11360_ ( .A1(_03659_ ), .A2(_03521_ ), .A3(_03570_ ), .ZN(_03660_ ) );
AOI21_X1 _11361_ ( .A(_03521_ ), .B1(_03659_ ), .B2(_03570_ ), .ZN(_03661_ ) );
OAI21_X1 _11362_ ( .A(_03437_ ), .B1(_03660_ ), .B2(_03661_ ), .ZN(_03662_ ) );
OAI211_X1 _11363_ ( .A(_03662_ ), .B(_03626_ ), .C1(\myexu.pc_jump [16] ), .C2(_03627_ ), .ZN(_03663_ ) );
NAND2_X1 _11364_ ( .A1(\mtvec [16] ), .A2(fanout_net_41 ), .ZN(_03664_ ) );
AOI21_X1 _11365_ ( .A(fanout_net_2 ), .B1(_03663_ ), .B2(_03664_ ), .ZN(_00252_ ) );
NOR2_X1 _11366_ ( .A1(_03433_ ), .A2(\mtvec [15] ), .ZN(_03665_ ) );
OR3_X1 _11367_ ( .A1(_03658_ ), .A2(_03654_ ), .A3(_03568_ ), .ZN(_03666_ ) );
NAND3_X1 _11368_ ( .A1(_03659_ ), .A2(_03627_ ), .A3(_03666_ ), .ZN(_03667_ ) );
AOI21_X1 _11369_ ( .A(fanout_net_41 ), .B1(_03618_ ), .B2(\myexu.pc_jump [15] ), .ZN(_03668_ ) );
AOI211_X1 _11370_ ( .A(fanout_net_2 ), .B(_03665_ ), .C1(_03667_ ), .C2(_03668_ ), .ZN(_00253_ ) );
NAND2_X1 _11371_ ( .A1(_03657_ ), .A2(_03529_ ), .ZN(_03669_ ) );
AND3_X1 _11372_ ( .A1(_03669_ ), .A2(_03566_ ), .A3(_03532_ ), .ZN(_03670_ ) );
AOI21_X1 _11373_ ( .A(_03532_ ), .B1(_03669_ ), .B2(_03566_ ), .ZN(_03671_ ) );
OR3_X1 _11374_ ( .A1(_03670_ ), .A2(_03671_ ), .A3(_03617_ ), .ZN(_03672_ ) );
OAI211_X1 _11375_ ( .A(_03672_ ), .B(_03626_ ), .C1(\myexu.pc_jump [14] ), .C2(_03627_ ), .ZN(_03673_ ) );
NAND2_X1 _11376_ ( .A1(\mtvec [14] ), .A2(fanout_net_41 ), .ZN(_03674_ ) );
AOI21_X1 _11377_ ( .A(fanout_net_2 ), .B1(_03673_ ), .B2(_03674_ ), .ZN(_00254_ ) );
OR3_X1 _11378_ ( .A1(_03215_ ), .A2(_03216_ ), .A3(\myexu.pc_jump [13] ), .ZN(_03675_ ) );
XOR2_X1 _11379_ ( .A(_03657_ ), .B(_03529_ ), .Z(_03676_ ) );
OAI211_X1 _11380_ ( .A(_03626_ ), .B(_03675_ ), .C1(_03676_ ), .C2(_03618_ ), .ZN(_03677_ ) );
NAND2_X1 _11381_ ( .A1(\mtvec [13] ), .A2(fanout_net_41 ), .ZN(_03678_ ) );
AOI21_X1 _11382_ ( .A(fanout_net_2 ), .B1(_03677_ ), .B2(_03678_ ), .ZN(_00255_ ) );
AND2_X1 _11383_ ( .A1(_03516_ ), .A2(_03548_ ), .ZN(_03679_ ) );
NOR2_X1 _11384_ ( .A1(_03679_ ), .A2(_03547_ ), .ZN(_03680_ ) );
NAND2_X1 _11385_ ( .A1(_03680_ ), .A2(_03552_ ), .ZN(_03681_ ) );
NAND3_X1 _11386_ ( .A1(_03681_ ), .A2(_03536_ ), .A3(_03553_ ), .ZN(_03682_ ) );
NAND2_X1 _11387_ ( .A1(_03535_ ), .A2(\IF_ID_pc [11] ), .ZN(_03683_ ) );
AND2_X1 _11388_ ( .A1(_03539_ ), .A2(_03540_ ), .ZN(_03684_ ) );
AND3_X1 _11389_ ( .A1(_03682_ ), .A2(_03683_ ), .A3(_03684_ ), .ZN(_03685_ ) );
AOI21_X1 _11390_ ( .A(_03684_ ), .B1(_03682_ ), .B2(_03683_ ), .ZN(_03686_ ) );
OR3_X1 _11391_ ( .A1(_03685_ ), .A2(_03686_ ), .A3(_03617_ ), .ZN(_03687_ ) );
OAI211_X1 _11392_ ( .A(_03687_ ), .B(_03626_ ), .C1(\myexu.pc_jump [12] ), .C2(_03627_ ), .ZN(_03688_ ) );
NAND2_X1 _11393_ ( .A1(\mtvec [12] ), .A2(fanout_net_41 ), .ZN(_03689_ ) );
AOI21_X1 _11394_ ( .A(fanout_net_2 ), .B1(_03688_ ), .B2(_03689_ ), .ZN(_00256_ ) );
AND2_X1 _11395_ ( .A1(_03603_ ), .A2(_03610_ ), .ZN(_03690_ ) );
OAI21_X1 _11396_ ( .A(_03436_ ), .B1(_03690_ ), .B2(_03446_ ), .ZN(_03691_ ) );
AOI21_X1 _11397_ ( .A(_03691_ ), .B1(_03690_ ), .B2(_03446_ ), .ZN(_03692_ ) );
AOI211_X1 _11398_ ( .A(fanout_net_41 ), .B(_03692_ ), .C1(\myexu.pc_jump [29] ), .C2(_03618_ ), .ZN(_03693_ ) );
NOR2_X1 _11399_ ( .A1(_03620_ ), .A2(\mtvec [29] ), .ZN(_03694_ ) );
NOR3_X1 _11400_ ( .A1(_03693_ ), .A2(fanout_net_2 ), .A3(_03694_ ), .ZN(_00257_ ) );
AND3_X1 _11401_ ( .A1(_03681_ ), .A2(_03536_ ), .A3(_03553_ ), .ZN(_03695_ ) );
AOI21_X1 _11402_ ( .A(_03536_ ), .B1(_03681_ ), .B2(_03553_ ), .ZN(_03696_ ) );
OAI21_X1 _11403_ ( .A(_03437_ ), .B1(_03695_ ), .B2(_03696_ ), .ZN(_03697_ ) );
OAI211_X1 _11404_ ( .A(_03697_ ), .B(_03626_ ), .C1(\myexu.pc_jump [11] ), .C2(_03627_ ), .ZN(_03698_ ) );
NAND2_X1 _11405_ ( .A1(\mtvec [11] ), .A2(fanout_net_41 ), .ZN(_03699_ ) );
AOI21_X1 _11406_ ( .A(fanout_net_2 ), .B1(_03698_ ), .B2(_03699_ ), .ZN(_00258_ ) );
AOI221_X4 _11407_ ( .A(_03547_ ), .B1(_03552_ ), .B2(_03553_ ), .C1(_03516_ ), .C2(_03548_ ), .ZN(_03700_ ) );
NOR2_X1 _11408_ ( .A1(_03700_ ), .A2(_03217_ ), .ZN(_03701_ ) );
OAI211_X1 _11409_ ( .A(_03552_ ), .B(_03553_ ), .C1(_03679_ ), .C2(_03547_ ), .ZN(_03702_ ) );
AOI221_X4 _11410_ ( .A(fanout_net_41 ), .B1(\myexu.pc_jump [10] ), .B2(_03217_ ), .C1(_03701_ ), .C2(_03702_ ), .ZN(_03703_ ) );
NOR2_X1 _11411_ ( .A1(_03620_ ), .A2(\mtvec [10] ), .ZN(_03704_ ) );
NOR3_X1 _11412_ ( .A1(_03703_ ), .A2(fanout_net_2 ), .A3(_03704_ ), .ZN(_00259_ ) );
NOR3_X1 _11413_ ( .A1(_03508_ ), .A2(_03515_ ), .A3(_03548_ ), .ZN(_03705_ ) );
OAI21_X1 _11414_ ( .A(_03437_ ), .B1(_03679_ ), .B2(_03705_ ), .ZN(_03706_ ) );
OAI211_X1 _11415_ ( .A(_03706_ ), .B(_03626_ ), .C1(\myexu.pc_jump [9] ), .C2(_03622_ ), .ZN(_03707_ ) );
NAND2_X1 _11416_ ( .A1(\mtvec [9] ), .A2(fanout_net_41 ), .ZN(_03708_ ) );
AOI21_X1 _11417_ ( .A(fanout_net_2 ), .B1(_03707_ ), .B2(_03708_ ), .ZN(_00260_ ) );
AOI21_X1 _11418_ ( .A(_03494_ ), .B1(_03487_ ), .B2(_03488_ ), .ZN(_03709_ ) );
OR3_X1 _11419_ ( .A1(_03709_ ), .A2(_03510_ ), .A3(_03513_ ), .ZN(_03710_ ) );
NAND3_X1 _11420_ ( .A1(_03710_ ), .A2(_03506_ ), .A3(_03512_ ), .ZN(_03711_ ) );
NAND2_X1 _11421_ ( .A1(_03505_ ), .A2(\IF_ID_pc [7] ), .ZN(_03712_ ) );
NAND2_X1 _11422_ ( .A1(_03711_ ), .A2(_03712_ ), .ZN(_03713_ ) );
XNOR2_X1 _11423_ ( .A(_03713_ ), .B(_03503_ ), .ZN(_03714_ ) );
NOR2_X1 _11424_ ( .A1(_03714_ ), .A2(_03617_ ), .ZN(_03715_ ) );
AOI211_X1 _11425_ ( .A(fanout_net_41 ), .B(_03715_ ), .C1(\myexu.pc_jump [8] ), .C2(_03618_ ), .ZN(_03716_ ) );
NOR2_X1 _11426_ ( .A1(_03620_ ), .A2(\mtvec [8] ), .ZN(_03717_ ) );
NOR3_X1 _11427_ ( .A1(_03716_ ), .A2(fanout_net_2 ), .A3(_03717_ ), .ZN(_00261_ ) );
AND3_X1 _11428_ ( .A1(_03710_ ), .A2(_03506_ ), .A3(_03512_ ), .ZN(_03718_ ) );
AOI21_X1 _11429_ ( .A(_03506_ ), .B1(_03710_ ), .B2(_03512_ ), .ZN(_03719_ ) );
OAI21_X1 _11430_ ( .A(_03437_ ), .B1(_03718_ ), .B2(_03719_ ), .ZN(_03720_ ) );
OAI211_X1 _11431_ ( .A(_03720_ ), .B(_03626_ ), .C1(\myexu.pc_jump [7] ), .C2(_03622_ ), .ZN(_03721_ ) );
NAND2_X1 _11432_ ( .A1(\mtvec [7] ), .A2(fanout_net_41 ), .ZN(_03722_ ) );
AOI21_X1 _11433_ ( .A(fanout_net_2 ), .B1(_03721_ ), .B2(_03722_ ), .ZN(_00262_ ) );
NOR2_X1 _11434_ ( .A1(_03709_ ), .A2(_03513_ ), .ZN(_03723_ ) );
XNOR2_X1 _11435_ ( .A(_03723_ ), .B(_03498_ ), .ZN(_03724_ ) );
MUX2_X1 _11436_ ( .A(\myexu.pc_jump [6] ), .B(_03724_ ), .S(_03436_ ), .Z(_03725_ ) );
MUX2_X1 _11437_ ( .A(\mtvec [6] ), .B(_03725_ ), .S(_03432_ ), .Z(_03726_ ) );
AND2_X1 _11438_ ( .A1(_03726_ ), .A2(_01618_ ), .ZN(_00263_ ) );
AND3_X1 _11439_ ( .A1(_03487_ ), .A2(_03488_ ), .A3(_03494_ ), .ZN(_03727_ ) );
OAI21_X1 _11440_ ( .A(_03437_ ), .B1(_03727_ ), .B2(_03709_ ), .ZN(_03728_ ) );
OAI211_X1 _11441_ ( .A(_03728_ ), .B(_03433_ ), .C1(\myexu.pc_jump [5] ), .C2(_03622_ ), .ZN(_03729_ ) );
NAND2_X1 _11442_ ( .A1(\mtvec [5] ), .A2(fanout_net_41 ), .ZN(_03730_ ) );
AOI21_X1 _11443_ ( .A(fanout_net_2 ), .B1(_03729_ ), .B2(_03730_ ), .ZN(_00264_ ) );
AND2_X1 _11444_ ( .A1(\mtvec [4] ), .A2(fanout_net_41 ), .ZN(_03731_ ) );
XNOR2_X1 _11445_ ( .A(_03486_ ), .B(fanout_net_11 ), .ZN(_03732_ ) );
XNOR2_X1 _11446_ ( .A(_03482_ ), .B(_03732_ ), .ZN(_03733_ ) );
MUX2_X1 _11447_ ( .A(\myexu.pc_jump [4] ), .B(_03733_ ), .S(_03436_ ), .Z(_03734_ ) );
AOI21_X1 _11448_ ( .A(_03731_ ), .B1(_03734_ ), .B2(_03620_ ), .ZN(_03735_ ) );
NOR2_X1 _11449_ ( .A1(_03735_ ), .A2(fanout_net_2 ), .ZN(_00265_ ) );
AND2_X1 _11450_ ( .A1(\mtvec [3] ), .A2(fanout_net_41 ), .ZN(_03736_ ) );
XOR2_X1 _11451_ ( .A(_03474_ ), .B(_03479_ ), .Z(_03737_ ) );
MUX2_X1 _11452_ ( .A(\myexu.pc_jump [3] ), .B(_03737_ ), .S(_03436_ ), .Z(_03738_ ) );
AOI21_X1 _11453_ ( .A(_03736_ ), .B1(_03738_ ), .B2(_03620_ ), .ZN(_03739_ ) );
NOR2_X1 _11454_ ( .A1(_03739_ ), .A2(reset ), .ZN(_00266_ ) );
AND2_X1 _11455_ ( .A1(IDU_ready_IFU ), .A2(\myifu.state [1] ), .ZN(\myifu.pc_$_SDFFE_PP1P__Q_E ) );
INV_X1 _11456_ ( .A(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_03740_ ) );
AOI211_X1 _11457_ ( .A(_03731_ ), .B(_03740_ ), .C1(_03734_ ), .C2(_03432_ ), .ZN(_03741_ ) );
INV_X1 _11458_ ( .A(fanout_net_11 ), .ZN(_03742_ ) );
CLKBUF_X3 _11459_ ( .A(_03742_ ), .Z(_03743_ ) );
CLKBUF_X2 _11460_ ( .A(_03743_ ), .Z(_03744_ ) );
BUF_X2 _11461_ ( .A(_03744_ ), .Z(_03745_ ) );
AOI211_X1 _11462_ ( .A(reset ), .B(_03741_ ), .C1(_03745_ ), .C2(_03740_ ), .ZN(_00267_ ) );
NOR2_X1 _11463_ ( .A1(_03466_ ), .A2(_03471_ ), .ZN(_03746_ ) );
OAI22_X1 _11464_ ( .A1(_03472_ ), .A2(_03746_ ), .B1(_03216_ ), .B2(_03215_ ), .ZN(_03747_ ) );
OAI211_X1 _11465_ ( .A(_03747_ ), .B(_03433_ ), .C1(\myexu.pc_jump [2] ), .C2(_03622_ ), .ZN(_03748_ ) );
NAND2_X1 _11466_ ( .A1(\mtvec [2] ), .A2(fanout_net_41 ), .ZN(_03749_ ) );
AOI21_X1 _11467_ ( .A(reset ), .B1(_03748_ ), .B2(_03749_ ), .ZN(_00268_ ) );
AOI211_X1 _11468_ ( .A(_03736_ ), .B(_03740_ ), .C1(_03738_ ), .C2(_03432_ ), .ZN(_03750_ ) );
INV_X1 _11469_ ( .A(fanout_net_7 ), .ZN(_03751_ ) );
BUF_X4 _11470_ ( .A(_03751_ ), .Z(_03752_ ) );
BUF_X2 _11471_ ( .A(_03752_ ), .Z(_03753_ ) );
AOI211_X1 _11472_ ( .A(reset ), .B(_03750_ ), .C1(_03753_ ), .C2(_03740_ ), .ZN(_00269_ ) );
AND3_X1 _11473_ ( .A1(_03597_ ), .A2(_03598_ ), .A3(_03599_ ), .ZN(_03754_ ) );
OAI21_X1 _11474_ ( .A(_03602_ ), .B1(_03754_ ), .B2(_03605_ ), .ZN(_03755_ ) );
AND3_X1 _11475_ ( .A1(_03755_ ), .A2(_03601_ ), .A3(_03609_ ), .ZN(_03756_ ) );
AOI21_X1 _11476_ ( .A(_03601_ ), .B1(_03755_ ), .B2(_03609_ ), .ZN(_03757_ ) );
OR3_X1 _11477_ ( .A1(_03756_ ), .A2(_03757_ ), .A3(_03617_ ), .ZN(_03758_ ) );
OAI211_X1 _11478_ ( .A(_03758_ ), .B(_03433_ ), .C1(\myexu.pc_jump [28] ), .C2(_03622_ ), .ZN(_03759_ ) );
NAND2_X1 _11479_ ( .A1(\mtvec [28] ), .A2(fanout_net_41 ), .ZN(_03760_ ) );
AOI21_X1 _11480_ ( .A(reset ), .B1(_03759_ ), .B2(_03760_ ), .ZN(_00270_ ) );
XNOR2_X1 _11481_ ( .A(_03469_ ), .B(_03470_ ), .ZN(_03761_ ) );
AOI21_X1 _11482_ ( .A(_03761_ ), .B1(check_quest ), .B2(_03431_ ), .ZN(_03762_ ) );
AOI211_X1 _11483_ ( .A(fanout_net_41 ), .B(_03762_ ), .C1(\myexu.pc_jump [1] ), .C2(_03618_ ), .ZN(_03763_ ) );
NOR2_X1 _11484_ ( .A1(_03620_ ), .A2(\mtvec [1] ), .ZN(_03764_ ) );
NOR3_X1 _11485_ ( .A1(_03763_ ), .A2(reset ), .A3(_03764_ ), .ZN(_00271_ ) );
NAND3_X1 _11486_ ( .A1(_03597_ ), .A2(_03598_ ), .A3(_03599_ ), .ZN(_03765_ ) );
AND3_X1 _11487_ ( .A1(_03765_ ), .A2(_03602_ ), .A3(_03604_ ), .ZN(_03766_ ) );
AOI21_X1 _11488_ ( .A(_03602_ ), .B1(_03765_ ), .B2(_03604_ ), .ZN(_03767_ ) );
OR3_X1 _11489_ ( .A1(_03766_ ), .A2(_03767_ ), .A3(_03617_ ), .ZN(_03768_ ) );
OAI211_X1 _11490_ ( .A(_03768_ ), .B(_03433_ ), .C1(\myexu.pc_jump [27] ), .C2(_03622_ ), .ZN(_03769_ ) );
NAND2_X1 _11491_ ( .A1(\mtvec [27] ), .A2(fanout_net_41 ), .ZN(_03770_ ) );
AOI21_X1 _11492_ ( .A(reset ), .B1(_03769_ ), .B2(_03770_ ), .ZN(_00272_ ) );
NAND2_X1 _11493_ ( .A1(_03597_ ), .A2(_03599_ ), .ZN(_03771_ ) );
NAND2_X1 _11494_ ( .A1(_03444_ ), .A2(\IF_ID_pc [25] ), .ZN(_03772_ ) );
AND3_X1 _11495_ ( .A1(_03771_ ), .A2(_03772_ ), .A3(_03598_ ), .ZN(_03773_ ) );
AOI21_X1 _11496_ ( .A(_03598_ ), .B1(_03771_ ), .B2(_03772_ ), .ZN(_03774_ ) );
OR3_X1 _11497_ ( .A1(_03773_ ), .A2(_03774_ ), .A3(_03217_ ), .ZN(_03775_ ) );
OAI211_X1 _11498_ ( .A(_03775_ ), .B(_03433_ ), .C1(\myexu.pc_jump [26] ), .C2(_03622_ ), .ZN(_03776_ ) );
NAND2_X1 _11499_ ( .A1(\mtvec [26] ), .A2(fanout_net_41 ), .ZN(_03777_ ) );
AOI21_X1 _11500_ ( .A(reset ), .B1(_03776_ ), .B2(_03777_ ), .ZN(_00273_ ) );
NAND3_X1 _11501_ ( .A1(_03431_ ), .A2(check_quest ), .A3(\myexu.pc_jump [25] ), .ZN(_03778_ ) );
XNOR2_X1 _11502_ ( .A(_03597_ ), .B(_03599_ ), .ZN(_03779_ ) );
OAI211_X1 _11503_ ( .A(_03433_ ), .B(_03778_ ), .C1(_03779_ ), .C2(_03617_ ), .ZN(_03780_ ) );
OR2_X1 _11504_ ( .A1(_03432_ ), .A2(\mtvec [25] ), .ZN(_03781_ ) );
AND3_X1 _11505_ ( .A1(_03780_ ), .A2(_01592_ ), .A3(_03781_ ), .ZN(_00274_ ) );
NOR2_X1 _11506_ ( .A1(_03624_ ), .A2(_03592_ ), .ZN(_03782_ ) );
AOI21_X1 _11507_ ( .A(_03782_ ), .B1(_02007_ ), .B2(_03575_ ), .ZN(_03783_ ) );
OAI21_X1 _11508_ ( .A(_03584_ ), .B1(_03783_ ), .B2(_03591_ ), .ZN(_03784_ ) );
AND3_X1 _11509_ ( .A1(_03784_ ), .A2(_03595_ ), .A3(_03583_ ), .ZN(_03785_ ) );
AOI21_X1 _11510_ ( .A(_03583_ ), .B1(_03784_ ), .B2(_03595_ ), .ZN(_03786_ ) );
OR3_X1 _11511_ ( .A1(_03785_ ), .A2(_03786_ ), .A3(_03217_ ), .ZN(_03787_ ) );
OAI211_X1 _11512_ ( .A(_03787_ ), .B(_03433_ ), .C1(\myexu.pc_jump [24] ), .C2(_03622_ ), .ZN(_03788_ ) );
NAND2_X1 _11513_ ( .A1(\mtvec [24] ), .A2(fanout_net_41 ), .ZN(_03789_ ) );
AOI21_X1 _11514_ ( .A(reset ), .B1(_03788_ ), .B2(_03789_ ), .ZN(_00275_ ) );
OR3_X1 _11515_ ( .A1(_03783_ ), .A2(_03584_ ), .A3(_03591_ ), .ZN(_03790_ ) );
AND3_X1 _11516_ ( .A1(_03790_ ), .A2(_03437_ ), .A3(_03784_ ), .ZN(_03791_ ) );
AOI211_X1 _11517_ ( .A(fanout_net_41 ), .B(_03791_ ), .C1(\myexu.pc_jump [23] ), .C2(_03618_ ), .ZN(_03792_ ) );
NOR2_X1 _11518_ ( .A1(_03620_ ), .A2(\mtvec [23] ), .ZN(_03793_ ) );
NOR3_X1 _11519_ ( .A1(_03792_ ), .A2(reset ), .A3(_03793_ ), .ZN(_00276_ ) );
XNOR2_X1 _11520_ ( .A(_03782_ ), .B(_03586_ ), .ZN(_03794_ ) );
NOR2_X1 _11521_ ( .A1(_03794_ ), .A2(_03617_ ), .ZN(_03795_ ) );
AOI211_X1 _11522_ ( .A(fanout_net_41 ), .B(_03795_ ), .C1(\myexu.pc_jump [22] ), .C2(_03617_ ), .ZN(_03796_ ) );
NOR2_X1 _11523_ ( .A1(_03620_ ), .A2(\mtvec [22] ), .ZN(_03797_ ) );
NOR3_X1 _11524_ ( .A1(_03796_ ), .A2(reset ), .A3(_03797_ ), .ZN(_00277_ ) );
NAND2_X1 _11525_ ( .A1(\mtvec [31] ), .A2(\myifu.to_reset ), .ZN(_03798_ ) );
OAI22_X1 _11526_ ( .A1(_03611_ ), .A2(_03612_ ), .B1(\IF_ID_pc [30] ), .B2(_03444_ ), .ZN(_03799_ ) );
NAND2_X1 _11527_ ( .A1(_03444_ ), .A2(\IF_ID_pc [30] ), .ZN(_03800_ ) );
NAND2_X1 _11528_ ( .A1(_03799_ ), .A2(_03800_ ), .ZN(_03801_ ) );
XNOR2_X1 _11529_ ( .A(_03444_ ), .B(\IF_ID_pc [31] ), .ZN(_03802_ ) );
OAI21_X1 _11530_ ( .A(_03437_ ), .B1(_03801_ ), .B2(_03802_ ), .ZN(_03803_ ) );
AOI21_X1 _11531_ ( .A(_03803_ ), .B1(_03801_ ), .B2(_03802_ ), .ZN(_03804_ ) );
OAI21_X1 _11532_ ( .A(_03433_ ), .B1(_03627_ ), .B2(\myexu.pc_jump [31] ), .ZN(_03805_ ) );
OAI211_X1 _11533_ ( .A(_01618_ ), .B(_03798_ ), .C1(_03804_ ), .C2(_03805_ ), .ZN(_00278_ ) );
OR3_X1 _11534_ ( .A1(_01993_ ), .A2(\myclint.state_r_$_NOT__A_Y ), .A3(_02019_ ), .ZN(_03806_ ) );
OAI21_X1 _11535_ ( .A(io_master_rvalid ), .B1(_01993_ ), .B2(_02019_ ), .ZN(_03807_ ) );
AND2_X1 _11536_ ( .A1(_03806_ ), .A2(_03807_ ), .ZN(_03808_ ) );
BUF_X2 _11537_ ( .A(_03808_ ), .Z(_03809_ ) );
AND2_X4 _11538_ ( .A1(_02065_ ), .A2(_02068_ ), .ZN(_03810_ ) );
BUF_X4 _11539_ ( .A(_03810_ ), .Z(_03811_ ) );
BUF_X4 _11540_ ( .A(_03811_ ), .Z(_03812_ ) );
BUF_X2 _11541_ ( .A(_03812_ ), .Z(_03813_ ) );
BUF_X4 _11542_ ( .A(_03813_ ), .Z(_03814_ ) );
NOR2_X1 _11543_ ( .A1(_03814_ ), .A2(io_master_rlast ), .ZN(_03815_ ) );
CLKBUF_X2 _11544_ ( .A(_02020_ ), .Z(_03816_ ) );
NOR2_X1 _11545_ ( .A1(_01993_ ), .A2(_02019_ ), .ZN(_03817_ ) );
INV_X1 _11546_ ( .A(\io_master_rid [1] ), .ZN(_03818_ ) );
NOR2_X1 _11547_ ( .A1(\io_master_rresp [1] ), .A2(\io_master_rresp [0] ), .ZN(_03819_ ) );
NOR2_X1 _11548_ ( .A1(\io_master_rid [3] ), .A2(\io_master_rid [2] ), .ZN(_03820_ ) );
AND4_X1 _11549_ ( .A1(_03818_ ), .A2(_03819_ ), .A3(_03820_ ), .A4(\io_master_rid [0] ), .ZN(_03821_ ) );
OAI21_X1 _11550_ ( .A(_03816_ ), .B1(_03817_ ), .B2(_03821_ ), .ZN(_03822_ ) );
BUF_X2 _11551_ ( .A(_03822_ ), .Z(_03823_ ) );
OR3_X1 _11552_ ( .A1(_03809_ ), .A2(_03815_ ), .A3(_03823_ ), .ZN(_03824_ ) );
INV_X1 _11553_ ( .A(\myifu.tmp_offset [2] ), .ZN(_03825_ ) );
AND3_X1 _11554_ ( .A1(_03824_ ), .A2(_01592_ ), .A3(_03825_ ), .ZN(_00279_ ) );
NOR3_X1 _11555_ ( .A1(reset ), .A2(\myifu.state [1] ), .A3(\myifu.state [2] ), .ZN(_00280_ ) );
AND3_X1 _11556_ ( .A1(_02080_ ), .A2(_03218_ ), .A3(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_03826_ ) );
INV_X1 _11557_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .ZN(_03827_ ) );
MUX2_X1 _11558_ ( .A(_02080_ ), .B(_03827_ ), .S(\myifu.to_reset ), .Z(_03828_ ) );
AOI211_X1 _11559_ ( .A(reset ), .B(_03826_ ), .C1(_03828_ ), .C2(\myifu.state [1] ), .ZN(_00281_ ) );
INV_X1 _11560_ ( .A(_02045_ ), .ZN(_03829_ ) );
NOR2_X1 _11561_ ( .A1(_02055_ ), .A2(_03829_ ), .ZN(_03830_ ) );
INV_X1 _11562_ ( .A(_03830_ ), .ZN(_03831_ ) );
BUF_X2 _11563_ ( .A(_03831_ ), .Z(_03832_ ) );
BUF_X4 _11564_ ( .A(_02092_ ), .Z(_03833_ ) );
BUF_X4 _11565_ ( .A(_03833_ ), .Z(_03834_ ) );
MUX2_X1 _11566_ ( .A(\LS_WB_waddr_csreg [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_03834_ ), .Z(_03835_ ) );
NOR2_X1 _11567_ ( .A1(_02049_ ), .A2(\EX_LS_flag [1] ), .ZN(_03836_ ) );
OR2_X1 _11568_ ( .A1(_03836_ ), .A2(_01989_ ), .ZN(_03837_ ) );
NOR2_X1 _11569_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_03838_ ) );
AND2_X2 _11570_ ( .A1(_03838_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_03839_ ) );
NOR2_X1 _11571_ ( .A1(_03837_ ), .A2(_03839_ ), .ZN(_03840_ ) );
BUF_X4 _11572_ ( .A(_03840_ ), .Z(_03841_ ) );
BUF_X4 _11573_ ( .A(_03841_ ), .Z(_03842_ ) );
BUF_X2 _11574_ ( .A(_03842_ ), .Z(_03843_ ) );
AND3_X1 _11575_ ( .A1(_03832_ ), .A2(_03835_ ), .A3(_03843_ ), .ZN(_00284_ ) );
BUF_X4 _11576_ ( .A(_02023_ ), .Z(_03844_ ) );
NOR2_X1 _11577_ ( .A1(_03830_ ), .A2(_03839_ ), .ZN(_03845_ ) );
INV_X1 _11578_ ( .A(_03845_ ), .ZN(_03846_ ) );
NAND3_X1 _11579_ ( .A1(_02044_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\EX_LS_flag [2] ), .ZN(_03847_ ) );
BUF_X4 _11580_ ( .A(_02049_ ), .Z(_03848_ ) );
NAND2_X1 _11581_ ( .A1(_03848_ ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_03849_ ) );
AOI211_X1 _11582_ ( .A(_03844_ ), .B(_03846_ ), .C1(_03847_ ), .C2(_03849_ ), .ZN(_00285_ ) );
NAND3_X1 _11583_ ( .A1(_02044_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(\EX_LS_flag [2] ), .ZN(_03850_ ) );
NAND2_X1 _11584_ ( .A1(_03848_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_03851_ ) );
AOI211_X1 _11585_ ( .A(_03844_ ), .B(_03846_ ), .C1(_03850_ ), .C2(_03851_ ), .ZN(_00286_ ) );
NAND3_X1 _11586_ ( .A1(_02044_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(\EX_LS_flag [2] ), .ZN(_03852_ ) );
NAND2_X1 _11587_ ( .A1(_03848_ ), .A2(\LS_WB_waddr_csreg [5] ), .ZN(_03853_ ) );
AOI211_X1 _11588_ ( .A(_03844_ ), .B(_03846_ ), .C1(_03852_ ), .C2(_03853_ ), .ZN(_00287_ ) );
NAND3_X1 _11589_ ( .A1(_02044_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\EX_LS_flag [2] ), .ZN(_03854_ ) );
NAND2_X1 _11590_ ( .A1(_03848_ ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_03855_ ) );
AOI211_X1 _11591_ ( .A(_03844_ ), .B(_03846_ ), .C1(_03854_ ), .C2(_03855_ ), .ZN(_00288_ ) );
NAND3_X1 _11592_ ( .A1(_02044_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(\EX_LS_flag [2] ), .ZN(_03856_ ) );
NAND2_X1 _11593_ ( .A1(_03848_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_03857_ ) );
AOI211_X1 _11594_ ( .A(_03844_ ), .B(_03846_ ), .C1(_03856_ ), .C2(_03857_ ), .ZN(_00289_ ) );
NAND3_X1 _11595_ ( .A1(_02044_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\EX_LS_flag [2] ), .ZN(_03858_ ) );
NAND2_X1 _11596_ ( .A1(_03848_ ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_03859_ ) );
AOI211_X1 _11597_ ( .A(_03844_ ), .B(_03846_ ), .C1(_03858_ ), .C2(_03859_ ), .ZN(_00290_ ) );
NAND3_X1 _11598_ ( .A1(_02044_ ), .A2(fanout_net_4 ), .A3(\EX_LS_flag [2] ), .ZN(_03860_ ) );
NAND2_X1 _11599_ ( .A1(_03848_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_03861_ ) );
AOI211_X1 _11600_ ( .A(_03844_ ), .B(_03846_ ), .C1(_03860_ ), .C2(_03861_ ), .ZN(_00291_ ) );
INV_X1 _11601_ ( .A(_02023_ ), .ZN(_03862_ ) );
NOR4_X1 _11602_ ( .A1(_03848_ ), .A2(_02042_ ), .A3(\EX_LS_dest_csreg_mem [9] ), .A4(\EX_LS_flag [0] ), .ZN(_03863_ ) );
NOR2_X1 _11603_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [9] ), .ZN(_03864_ ) );
OAI211_X1 _11604_ ( .A(_03845_ ), .B(_03862_ ), .C1(_03863_ ), .C2(_03864_ ), .ZN(_00292_ ) );
NOR4_X1 _11605_ ( .A1(_03848_ ), .A2(_02042_ ), .A3(\EX_LS_dest_csreg_mem [8] ), .A4(\EX_LS_flag [0] ), .ZN(_03865_ ) );
NOR2_X1 _11606_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_03866_ ) );
OAI211_X1 _11607_ ( .A(_03845_ ), .B(_03862_ ), .C1(_03865_ ), .C2(_03866_ ), .ZN(_00293_ ) );
NOR4_X1 _11608_ ( .A1(_02049_ ), .A2(_02042_ ), .A3(\EX_LS_dest_csreg_mem [6] ), .A4(\EX_LS_flag [0] ), .ZN(_03867_ ) );
NOR2_X1 _11609_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_03868_ ) );
OAI211_X1 _11610_ ( .A(_03845_ ), .B(_03862_ ), .C1(_03867_ ), .C2(_03868_ ), .ZN(_00294_ ) );
NOR4_X1 _11611_ ( .A1(_02049_ ), .A2(_02042_ ), .A3(fanout_net_3 ), .A4(\EX_LS_flag [0] ), .ZN(_03869_ ) );
NOR2_X1 _11612_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [0] ), .ZN(_03870_ ) );
OAI211_X1 _11613_ ( .A(_03845_ ), .B(_03862_ ), .C1(_03869_ ), .C2(_03870_ ), .ZN(_00295_ ) );
INV_X1 _11614_ ( .A(\mysc.state [2] ), .ZN(_03871_ ) );
NOR2_X1 _11615_ ( .A1(_03871_ ), .A2(reset ), .ZN(_00303_ ) );
AND3_X1 _11616_ ( .A1(_01548_ ), .A2(\LS_WB_wen_csreg [6] ), .A3(\LS_WB_wen_csreg [7] ), .ZN(_00093_ ) );
INV_X1 _11617_ ( .A(IDU_valid_EXU ), .ZN(_03872_ ) );
NOR2_X1 _11618_ ( .A1(_03872_ ), .A2(EXU_valid_LSU ), .ZN(\myexu.state_$_ANDNOT__B_Y ) );
INV_X1 _11619_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .ZN(_03873_ ) );
NOR2_X1 _11620_ ( .A1(_03341_ ), .A2(\ID_EX_typ [6] ), .ZN(_03874_ ) );
AND2_X1 _11621_ ( .A1(_03874_ ), .A2(\ID_EX_typ [5] ), .ZN(_03875_ ) );
BUF_X4 _11622_ ( .A(_03875_ ), .Z(_03876_ ) );
INV_X1 _11623_ ( .A(fanout_net_5 ), .ZN(_03877_ ) );
AND2_X1 _11624_ ( .A1(_03876_ ), .A2(_03877_ ), .ZN(_03878_ ) );
INV_X1 _11625_ ( .A(_03878_ ), .ZN(_03879_ ) );
NOR2_X1 _11626_ ( .A1(\ID_EX_typ [5] ), .A2(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03880_ ) );
INV_X1 _11627_ ( .A(\ID_EX_typ [6] ), .ZN(_03881_ ) );
NAND3_X1 _11628_ ( .A1(_03880_ ), .A2(\ID_EX_typ [7] ), .A3(_03881_ ), .ZN(_03882_ ) );
AOI21_X1 _11629_ ( .A(_03873_ ), .B1(_03879_ ), .B2(_03882_ ), .ZN(_03883_ ) );
INV_X1 _11630_ ( .A(\myec.state [1] ), .ZN(_03884_ ) );
NAND2_X1 _11631_ ( .A1(_03884_ ), .A2(\myec.state [0] ), .ZN(_03885_ ) );
AND2_X1 _11632_ ( .A1(_03885_ ), .A2(_03065_ ), .ZN(_03886_ ) );
BUF_X2 _11633_ ( .A(_03886_ ), .Z(_03887_ ) );
AND4_X1 _11634_ ( .A1(\ID_EX_typ [7] ), .A2(_03881_ ), .A3(_01986_ ), .A4(IDU_valid_EXU ), .ZN(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _11635_ ( .A1(_03216_ ), .A2(check_assert ), .ZN(_03888_ ) );
OAI21_X1 _11636_ ( .A(_03887_ ), .B1(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(_03888_ ), .ZN(_03889_ ) );
NOR2_X1 _11637_ ( .A1(_03883_ ), .A2(_03889_ ), .ZN(_00096_ ) );
CLKBUF_X2 _11638_ ( .A(_03885_ ), .Z(_03890_ ) );
CLKBUF_X2 _11639_ ( .A(_03890_ ), .Z(_03891_ ) );
AND3_X1 _11640_ ( .A1(_03891_ ), .A2(\ID_EX_rd [4] ), .A3(_03083_ ), .ZN(_00117_ ) );
AND3_X1 _11641_ ( .A1(_03891_ ), .A2(\ID_EX_rd [3] ), .A3(_03083_ ), .ZN(_00118_ ) );
AND3_X1 _11642_ ( .A1(_03891_ ), .A2(\ID_EX_rd [2] ), .A3(_03083_ ), .ZN(_00119_ ) );
AND3_X1 _11643_ ( .A1(_03891_ ), .A2(\ID_EX_rd [1] ), .A3(_03083_ ), .ZN(_00120_ ) );
AND3_X1 _11644_ ( .A1(_03891_ ), .A2(\ID_EX_rd [0] ), .A3(_03083_ ), .ZN(_00121_ ) );
BUF_X4 _11645_ ( .A(_03876_ ), .Z(_03892_ ) );
AND2_X1 _11646_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_pc [2] ), .ZN(_03893_ ) );
AND2_X1 _11647_ ( .A1(_03893_ ), .A2(\ID_EX_pc [4] ), .ZN(_03894_ ) );
AND2_X1 _11648_ ( .A1(_03894_ ), .A2(\ID_EX_pc [5] ), .ZN(_03895_ ) );
AND2_X1 _11649_ ( .A1(_03895_ ), .A2(\ID_EX_pc [6] ), .ZN(_03896_ ) );
AND2_X1 _11650_ ( .A1(_03896_ ), .A2(\ID_EX_pc [7] ), .ZN(_03897_ ) );
AND2_X1 _11651_ ( .A1(_03897_ ), .A2(\ID_EX_pc [8] ), .ZN(_03898_ ) );
AND2_X1 _11652_ ( .A1(_03898_ ), .A2(\ID_EX_pc [9] ), .ZN(_03899_ ) );
AND2_X1 _11653_ ( .A1(_03899_ ), .A2(\ID_EX_pc [10] ), .ZN(_03900_ ) );
AND2_X1 _11654_ ( .A1(_03900_ ), .A2(\ID_EX_pc [11] ), .ZN(_03901_ ) );
AND3_X1 _11655_ ( .A1(_03901_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_03902_ ) );
AND3_X1 _11656_ ( .A1(_03902_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_03903_ ) );
AND3_X1 _11657_ ( .A1(_03903_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_pc [16] ), .ZN(_03904_ ) );
AND3_X1 _11658_ ( .A1(_03904_ ), .A2(\ID_EX_pc [19] ), .A3(\ID_EX_pc [18] ), .ZN(_03905_ ) );
AND3_X1 _11659_ ( .A1(_03905_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_03906_ ) );
AND3_X1 _11660_ ( .A1(_03906_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_03907_ ) );
AND3_X1 _11661_ ( .A1(_03907_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_pc [24] ), .ZN(_03908_ ) );
AND3_X1 _11662_ ( .A1(_03908_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_03909_ ) );
NAND3_X1 _11663_ ( .A1(_03909_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_03910_ ) );
INV_X1 _11664_ ( .A(\ID_EX_pc [30] ), .ZN(_03911_ ) );
XNOR2_X1 _11665_ ( .A(_03910_ ), .B(_03911_ ), .ZN(_03912_ ) );
NOR2_X1 _11666_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_5 ), .ZN(_03913_ ) );
AND2_X1 _11667_ ( .A1(_03913_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_03914_ ) );
INV_X1 _11668_ ( .A(_03914_ ), .ZN(_03915_ ) );
INV_X1 _11669_ ( .A(_02765_ ), .ZN(_03916_ ) );
XOR2_X2 _11670_ ( .A(\EX_LS_dest_reg [4] ), .B(\ID_EX_rs2 [4] ), .Z(_03917_ ) );
INV_X2 _11671_ ( .A(_03917_ ), .ZN(_03918_ ) );
XNOR2_X1 _11672_ ( .A(\EX_LS_dest_reg [3] ), .B(\ID_EX_rs2 [3] ), .ZN(_03919_ ) );
XNOR2_X1 _11673_ ( .A(\EX_LS_dest_reg [1] ), .B(\ID_EX_rs2 [1] ), .ZN(_03920_ ) );
XNOR2_X1 _11674_ ( .A(\EX_LS_dest_reg [0] ), .B(\ID_EX_rs2 [0] ), .ZN(_03921_ ) );
XNOR2_X1 _11675_ ( .A(\EX_LS_dest_reg [2] ), .B(\ID_EX_rs2 [2] ), .ZN(_03922_ ) );
AND4_X1 _11676_ ( .A1(_03919_ ), .A2(_03920_ ), .A3(_03921_ ), .A4(_03922_ ), .ZN(_03923_ ) );
NAND4_X4 _11677_ ( .A1(_02094_ ), .A2(_02099_ ), .A3(_03918_ ), .A4(_03923_ ), .ZN(_03924_ ) );
BUF_X2 _11678_ ( .A(_03924_ ), .Z(_03925_ ) );
INV_X1 _11679_ ( .A(\EX_LS_result_reg [11] ), .ZN(_03926_ ) );
INV_X1 _11680_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .ZN(_03927_ ) );
OR3_X1 _11681_ ( .A1(_03925_ ), .A2(_03926_ ), .A3(_03927_ ), .ZN(_03928_ ) );
INV_X1 _11682_ ( .A(fanout_net_39 ), .ZN(_03929_ ) );
BUF_X4 _11683_ ( .A(_03929_ ), .Z(_03930_ ) );
OR2_X1 _11684_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[0][11] ), .ZN(_03931_ ) );
INV_X1 _11685_ ( .A(fanout_net_36 ), .ZN(_03932_ ) );
BUF_X4 _11686_ ( .A(_03932_ ), .Z(_03933_ ) );
BUF_X4 _11687_ ( .A(_03933_ ), .Z(_03934_ ) );
INV_X1 _11688_ ( .A(fanout_net_28 ), .ZN(_03935_ ) );
BUF_X4 _11689_ ( .A(_03935_ ), .Z(_03936_ ) );
BUF_X4 _11690_ ( .A(_03936_ ), .Z(_03937_ ) );
OAI211_X1 _11691_ ( .A(_03931_ ), .B(_03934_ ), .C1(_03937_ ), .C2(\myreg.Reg[1][11] ), .ZN(_03938_ ) );
OR2_X1 _11692_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[2][11] ), .ZN(_03939_ ) );
BUF_X4 _11693_ ( .A(_03936_ ), .Z(_03940_ ) );
OAI211_X1 _11694_ ( .A(_03939_ ), .B(fanout_net_36 ), .C1(_03940_ ), .C2(\myreg.Reg[3][11] ), .ZN(_03941_ ) );
INV_X1 _11695_ ( .A(fanout_net_38 ), .ZN(_03942_ ) );
BUF_X4 _11696_ ( .A(_03942_ ), .Z(_03943_ ) );
NAND3_X1 _11697_ ( .A1(_03938_ ), .A2(_03941_ ), .A3(_03943_ ), .ZN(_03944_ ) );
MUX2_X1 _11698_ ( .A(\myreg.Reg[6][11] ), .B(\myreg.Reg[7][11] ), .S(fanout_net_28 ), .Z(_03945_ ) );
MUX2_X1 _11699_ ( .A(\myreg.Reg[4][11] ), .B(\myreg.Reg[5][11] ), .S(fanout_net_28 ), .Z(_03946_ ) );
BUF_X4 _11700_ ( .A(_03932_ ), .Z(_03947_ ) );
MUX2_X1 _11701_ ( .A(_03945_ ), .B(_03946_ ), .S(_03947_ ), .Z(_03948_ ) );
BUF_X4 _11702_ ( .A(_03942_ ), .Z(_03949_ ) );
BUF_X4 _11703_ ( .A(_03949_ ), .Z(_03950_ ) );
OAI211_X1 _11704_ ( .A(_03930_ ), .B(_03944_ ), .C1(_03948_ ), .C2(_03950_ ), .ZN(_03951_ ) );
OR2_X1 _11705_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[14][11] ), .ZN(_03952_ ) );
OAI211_X1 _11706_ ( .A(_03952_ ), .B(fanout_net_36 ), .C1(_03937_ ), .C2(\myreg.Reg[15][11] ), .ZN(_03953_ ) );
OR2_X1 _11707_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[12][11] ), .ZN(_03954_ ) );
OAI211_X1 _11708_ ( .A(_03954_ ), .B(_03934_ ), .C1(_03940_ ), .C2(\myreg.Reg[13][11] ), .ZN(_03955_ ) );
NAND3_X1 _11709_ ( .A1(_03953_ ), .A2(_03955_ ), .A3(fanout_net_38 ), .ZN(_03956_ ) );
MUX2_X1 _11710_ ( .A(\myreg.Reg[8][11] ), .B(\myreg.Reg[9][11] ), .S(fanout_net_28 ), .Z(_03957_ ) );
MUX2_X1 _11711_ ( .A(\myreg.Reg[10][11] ), .B(\myreg.Reg[11][11] ), .S(fanout_net_28 ), .Z(_03958_ ) );
MUX2_X1 _11712_ ( .A(_03957_ ), .B(_03958_ ), .S(fanout_net_36 ), .Z(_03959_ ) );
OAI211_X1 _11713_ ( .A(fanout_net_39 ), .B(_03956_ ), .C1(_03959_ ), .C2(fanout_net_38 ), .ZN(_03960_ ) );
NAND2_X1 _11714_ ( .A1(_03951_ ), .A2(_03960_ ), .ZN(_03961_ ) );
BUF_X2 _11715_ ( .A(_03927_ ), .Z(_03962_ ) );
OAI21_X1 _11716_ ( .A(_03961_ ), .B1(_03925_ ), .B2(_03962_ ), .ZN(_03963_ ) );
AND2_X1 _11717_ ( .A1(_03928_ ), .A2(_03963_ ), .ZN(_03964_ ) );
XNOR2_X2 _11718_ ( .A(_03916_ ), .B(_03964_ ), .ZN(_03965_ ) );
BUF_X4 _11719_ ( .A(_03935_ ), .Z(_03966_ ) );
NOR2_X1 _11720_ ( .A1(_03966_ ), .A2(\myreg.Reg[11][10] ), .ZN(_03967_ ) );
OAI21_X1 _11721_ ( .A(fanout_net_36 ), .B1(fanout_net_28 ), .B2(\myreg.Reg[10][10] ), .ZN(_03968_ ) );
NOR2_X1 _11722_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[8][10] ), .ZN(_03969_ ) );
OAI21_X1 _11723_ ( .A(_03947_ ), .B1(_03966_ ), .B2(\myreg.Reg[9][10] ), .ZN(_03970_ ) );
OAI221_X1 _11724_ ( .A(_03943_ ), .B1(_03967_ ), .B2(_03968_ ), .C1(_03969_ ), .C2(_03970_ ), .ZN(_03971_ ) );
MUX2_X1 _11725_ ( .A(\myreg.Reg[12][10] ), .B(\myreg.Reg[13][10] ), .S(fanout_net_28 ), .Z(_03972_ ) );
MUX2_X1 _11726_ ( .A(\myreg.Reg[14][10] ), .B(\myreg.Reg[15][10] ), .S(fanout_net_28 ), .Z(_03973_ ) );
MUX2_X1 _11727_ ( .A(_03972_ ), .B(_03973_ ), .S(fanout_net_36 ), .Z(_03974_ ) );
OAI211_X1 _11728_ ( .A(fanout_net_39 ), .B(_03971_ ), .C1(_03974_ ), .C2(_03950_ ), .ZN(_03975_ ) );
OR2_X1 _11729_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[4][10] ), .ZN(_03976_ ) );
OAI211_X1 _11730_ ( .A(_03976_ ), .B(_03947_ ), .C1(_03940_ ), .C2(\myreg.Reg[5][10] ), .ZN(_03977_ ) );
OR2_X1 _11731_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[6][10] ), .ZN(_03978_ ) );
OAI211_X1 _11732_ ( .A(_03978_ ), .B(fanout_net_36 ), .C1(_03940_ ), .C2(\myreg.Reg[7][10] ), .ZN(_03979_ ) );
NAND3_X1 _11733_ ( .A1(_03977_ ), .A2(_03979_ ), .A3(fanout_net_38 ), .ZN(_03980_ ) );
MUX2_X1 _11734_ ( .A(\myreg.Reg[2][10] ), .B(\myreg.Reg[3][10] ), .S(fanout_net_28 ), .Z(_03981_ ) );
MUX2_X1 _11735_ ( .A(\myreg.Reg[0][10] ), .B(\myreg.Reg[1][10] ), .S(fanout_net_28 ), .Z(_03982_ ) );
MUX2_X1 _11736_ ( .A(_03981_ ), .B(_03982_ ), .S(_03947_ ), .Z(_03983_ ) );
OAI211_X1 _11737_ ( .A(_03930_ ), .B(_03980_ ), .C1(_03983_ ), .C2(fanout_net_38 ), .ZN(_03984_ ) );
NAND2_X1 _11738_ ( .A1(_03975_ ), .A2(_03984_ ), .ZN(_03985_ ) );
OAI21_X1 _11739_ ( .A(_03985_ ), .B1(_03925_ ), .B2(_03962_ ), .ZN(_03986_ ) );
OAI21_X1 _11740_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .B1(_02100_ ), .B2(\ID_EX_rs2 [1] ), .ZN(_03987_ ) );
AOI211_X1 _11741_ ( .A(_03987_ ), .B(_02098_ ), .C1(_02100_ ), .C2(\ID_EX_rs2 [1] ), .ZN(_03988_ ) );
AND4_X2 _11742_ ( .A1(_03919_ ), .A2(_03918_ ), .A3(_03921_ ), .A4(_03922_ ), .ZN(_03989_ ) );
NAND4_X1 _11743_ ( .A1(_02094_ ), .A2(\EX_LS_result_reg [10] ), .A3(_03988_ ), .A4(_03989_ ), .ZN(_03990_ ) );
AND2_X1 _11744_ ( .A1(_03986_ ), .A2(_03990_ ), .ZN(_03991_ ) );
XOR2_X1 _11745_ ( .A(_02741_ ), .B(_03991_ ), .Z(_03992_ ) );
AND2_X1 _11746_ ( .A1(_03965_ ), .A2(_03992_ ), .ZN(_03993_ ) );
NOR2_X4 _11747_ ( .A1(_03924_ ), .A2(_03927_ ), .ZN(_03994_ ) );
OR2_X1 _11748_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[4][8] ), .ZN(_03995_ ) );
BUF_X4 _11749_ ( .A(_03947_ ), .Z(_03996_ ) );
BUF_X4 _11750_ ( .A(_03966_ ), .Z(_03997_ ) );
OAI211_X1 _11751_ ( .A(_03995_ ), .B(_03996_ ), .C1(_03997_ ), .C2(\myreg.Reg[5][8] ), .ZN(_03998_ ) );
OR2_X1 _11752_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[6][8] ), .ZN(_03999_ ) );
BUF_X4 _11753_ ( .A(_03966_ ), .Z(_04000_ ) );
OAI211_X1 _11754_ ( .A(_03999_ ), .B(fanout_net_36 ), .C1(_04000_ ), .C2(\myreg.Reg[7][8] ), .ZN(_04001_ ) );
NAND3_X1 _11755_ ( .A1(_03998_ ), .A2(_04001_ ), .A3(fanout_net_38 ), .ZN(_04002_ ) );
MUX2_X1 _11756_ ( .A(\myreg.Reg[2][8] ), .B(\myreg.Reg[3][8] ), .S(fanout_net_28 ), .Z(_04003_ ) );
MUX2_X1 _11757_ ( .A(\myreg.Reg[0][8] ), .B(\myreg.Reg[1][8] ), .S(fanout_net_28 ), .Z(_04004_ ) );
BUF_X4 _11758_ ( .A(_03933_ ), .Z(_04005_ ) );
MUX2_X1 _11759_ ( .A(_04003_ ), .B(_04004_ ), .S(_04005_ ), .Z(_04006_ ) );
OAI211_X1 _11760_ ( .A(_03930_ ), .B(_04002_ ), .C1(_04006_ ), .C2(fanout_net_38 ), .ZN(_04007_ ) );
NOR2_X1 _11761_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[8][8] ), .ZN(_04008_ ) );
OAI21_X1 _11762_ ( .A(_03934_ ), .B1(_03940_ ), .B2(\myreg.Reg[9][8] ), .ZN(_04009_ ) );
AND2_X1 _11763_ ( .A1(_03966_ ), .A2(\myreg.Reg[10][8] ), .ZN(_04010_ ) );
AOI21_X1 _11764_ ( .A(_04010_ ), .B1(fanout_net_28 ), .B2(\myreg.Reg[11][8] ), .ZN(_04011_ ) );
BUF_X4 _11765_ ( .A(_03934_ ), .Z(_04012_ ) );
OAI221_X1 _11766_ ( .A(_03943_ ), .B1(_04008_ ), .B2(_04009_ ), .C1(_04011_ ), .C2(_04012_ ), .ZN(_04013_ ) );
BUF_X4 _11767_ ( .A(_03943_ ), .Z(_04014_ ) );
MUX2_X1 _11768_ ( .A(\myreg.Reg[12][8] ), .B(\myreg.Reg[13][8] ), .S(fanout_net_28 ), .Z(_04015_ ) );
MUX2_X1 _11769_ ( .A(\myreg.Reg[14][8] ), .B(\myreg.Reg[15][8] ), .S(fanout_net_28 ), .Z(_04016_ ) );
MUX2_X1 _11770_ ( .A(_04015_ ), .B(_04016_ ), .S(fanout_net_36 ), .Z(_04017_ ) );
OAI211_X1 _11771_ ( .A(_04013_ ), .B(fanout_net_39 ), .C1(_04014_ ), .C2(_04017_ ), .ZN(_04018_ ) );
AOI21_X1 _11772_ ( .A(_03994_ ), .B1(_04007_ ), .B2(_04018_ ), .ZN(_04019_ ) );
AND4_X1 _11773_ ( .A1(\EX_LS_result_reg [8] ), .A2(_02094_ ), .A3(_03989_ ), .A4(_03988_ ), .ZN(_04020_ ) );
NOR2_X1 _11774_ ( .A1(_04019_ ), .A2(_04020_ ), .ZN(_04021_ ) );
INV_X1 _11775_ ( .A(_02789_ ), .ZN(_04022_ ) );
XNOR2_X1 _11776_ ( .A(_04021_ ), .B(_04022_ ), .ZN(_04023_ ) );
INV_X1 _11777_ ( .A(_02812_ ), .ZN(_04024_ ) );
INV_X1 _11778_ ( .A(\EX_LS_result_reg [9] ), .ZN(_04025_ ) );
OR3_X1 _11779_ ( .A1(_03924_ ), .A2(_04025_ ), .A3(_03927_ ), .ZN(_04026_ ) );
OR2_X1 _11780_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[0][9] ), .ZN(_04027_ ) );
OAI211_X1 _11781_ ( .A(_04027_ ), .B(_03932_ ), .C1(_03936_ ), .C2(\myreg.Reg[1][9] ), .ZN(_04028_ ) );
OR2_X1 _11782_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[2][9] ), .ZN(_04029_ ) );
OAI211_X1 _11783_ ( .A(_04029_ ), .B(fanout_net_36 ), .C1(_03935_ ), .C2(\myreg.Reg[3][9] ), .ZN(_04030_ ) );
NAND3_X1 _11784_ ( .A1(_04028_ ), .A2(_04030_ ), .A3(_03942_ ), .ZN(_04031_ ) );
MUX2_X1 _11785_ ( .A(\myreg.Reg[6][9] ), .B(\myreg.Reg[7][9] ), .S(fanout_net_28 ), .Z(_04032_ ) );
MUX2_X1 _11786_ ( .A(\myreg.Reg[4][9] ), .B(\myreg.Reg[5][9] ), .S(fanout_net_28 ), .Z(_04033_ ) );
MUX2_X1 _11787_ ( .A(_04032_ ), .B(_04033_ ), .S(_03932_ ), .Z(_04034_ ) );
OAI211_X1 _11788_ ( .A(_03929_ ), .B(_04031_ ), .C1(_04034_ ), .C2(_03949_ ), .ZN(_04035_ ) );
OR2_X1 _11789_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[14][9] ), .ZN(_04036_ ) );
OAI211_X1 _11790_ ( .A(_04036_ ), .B(fanout_net_36 ), .C1(_03935_ ), .C2(\myreg.Reg[15][9] ), .ZN(_04037_ ) );
OR2_X1 _11791_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[12][9] ), .ZN(_04038_ ) );
OAI211_X1 _11792_ ( .A(_04038_ ), .B(_03932_ ), .C1(_03935_ ), .C2(\myreg.Reg[13][9] ), .ZN(_04039_ ) );
NAND3_X1 _11793_ ( .A1(_04037_ ), .A2(_04039_ ), .A3(fanout_net_38 ), .ZN(_04040_ ) );
MUX2_X1 _11794_ ( .A(\myreg.Reg[8][9] ), .B(\myreg.Reg[9][9] ), .S(fanout_net_29 ), .Z(_04041_ ) );
MUX2_X1 _11795_ ( .A(\myreg.Reg[10][9] ), .B(\myreg.Reg[11][9] ), .S(fanout_net_29 ), .Z(_04042_ ) );
MUX2_X1 _11796_ ( .A(_04041_ ), .B(_04042_ ), .S(fanout_net_36 ), .Z(_04043_ ) );
OAI211_X1 _11797_ ( .A(fanout_net_39 ), .B(_04040_ ), .C1(_04043_ ), .C2(fanout_net_38 ), .ZN(_04044_ ) );
NAND2_X1 _11798_ ( .A1(_04035_ ), .A2(_04044_ ), .ZN(_04045_ ) );
OAI21_X1 _11799_ ( .A(_04045_ ), .B1(_03924_ ), .B2(_03927_ ), .ZN(_04046_ ) );
AND2_X2 _11800_ ( .A1(_04026_ ), .A2(_04046_ ), .ZN(_04047_ ) );
XNOR2_X1 _11801_ ( .A(_04024_ ), .B(_04047_ ), .ZN(_04048_ ) );
AND3_X1 _11802_ ( .A1(_03993_ ), .A2(_04023_ ), .A3(_04048_ ), .ZN(_04049_ ) );
INV_X1 _11803_ ( .A(_04049_ ), .ZN(_04050_ ) );
INV_X1 _11804_ ( .A(\EX_LS_result_reg [13] ), .ZN(_04051_ ) );
OR3_X1 _11805_ ( .A1(_03925_ ), .A2(_04051_ ), .A3(_03962_ ), .ZN(_04052_ ) );
OR2_X1 _11806_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[0][13] ), .ZN(_04053_ ) );
OAI211_X1 _11807_ ( .A(_04053_ ), .B(_03996_ ), .C1(_03997_ ), .C2(\myreg.Reg[1][13] ), .ZN(_04054_ ) );
OR2_X1 _11808_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[2][13] ), .ZN(_04055_ ) );
OAI211_X1 _11809_ ( .A(_04055_ ), .B(fanout_net_36 ), .C1(_04000_ ), .C2(\myreg.Reg[3][13] ), .ZN(_04056_ ) );
NAND3_X1 _11810_ ( .A1(_04054_ ), .A2(_04056_ ), .A3(_03950_ ), .ZN(_04057_ ) );
MUX2_X1 _11811_ ( .A(\myreg.Reg[6][13] ), .B(\myreg.Reg[7][13] ), .S(fanout_net_29 ), .Z(_04058_ ) );
MUX2_X1 _11812_ ( .A(\myreg.Reg[4][13] ), .B(\myreg.Reg[5][13] ), .S(fanout_net_29 ), .Z(_04059_ ) );
MUX2_X1 _11813_ ( .A(_04058_ ), .B(_04059_ ), .S(_04005_ ), .Z(_04060_ ) );
OAI211_X1 _11814_ ( .A(_03930_ ), .B(_04057_ ), .C1(_04060_ ), .C2(_04014_ ), .ZN(_04061_ ) );
OR2_X1 _11815_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[14][13] ), .ZN(_04062_ ) );
OAI211_X1 _11816_ ( .A(_04062_ ), .B(fanout_net_36 ), .C1(_04000_ ), .C2(\myreg.Reg[15][13] ), .ZN(_04063_ ) );
OR2_X1 _11817_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[12][13] ), .ZN(_04064_ ) );
OAI211_X1 _11818_ ( .A(_04064_ ), .B(_04005_ ), .C1(_04000_ ), .C2(\myreg.Reg[13][13] ), .ZN(_04065_ ) );
NAND3_X1 _11819_ ( .A1(_04063_ ), .A2(_04065_ ), .A3(fanout_net_38 ), .ZN(_04066_ ) );
MUX2_X1 _11820_ ( .A(\myreg.Reg[8][13] ), .B(\myreg.Reg[9][13] ), .S(fanout_net_29 ), .Z(_04067_ ) );
MUX2_X1 _11821_ ( .A(\myreg.Reg[10][13] ), .B(\myreg.Reg[11][13] ), .S(fanout_net_29 ), .Z(_04068_ ) );
MUX2_X1 _11822_ ( .A(_04067_ ), .B(_04068_ ), .S(fanout_net_36 ), .Z(_04069_ ) );
OAI211_X1 _11823_ ( .A(fanout_net_39 ), .B(_04066_ ), .C1(_04069_ ), .C2(fanout_net_38 ), .ZN(_04070_ ) );
NAND2_X1 _11824_ ( .A1(_04061_ ), .A2(_04070_ ), .ZN(_04071_ ) );
BUF_X2 _11825_ ( .A(_03962_ ), .Z(_04072_ ) );
OAI21_X1 _11826_ ( .A(_04071_ ), .B1(_03925_ ), .B2(_04072_ ), .ZN(_04073_ ) );
AND2_X1 _11827_ ( .A1(_04052_ ), .A2(_04073_ ), .ZN(_04074_ ) );
NAND2_X1 _11828_ ( .A1(_02667_ ), .A2(_02668_ ), .ZN(_04075_ ) );
AND2_X1 _11829_ ( .A1(_04074_ ), .A2(_04075_ ), .ZN(_04076_ ) );
NOR2_X1 _11830_ ( .A1(_04074_ ), .A2(_04075_ ), .ZN(_04077_ ) );
NOR2_X1 _11831_ ( .A1(_04076_ ), .A2(_04077_ ), .ZN(_04078_ ) );
INV_X1 _11832_ ( .A(_02647_ ), .ZN(_04079_ ) );
INV_X1 _11833_ ( .A(\EX_LS_result_reg [12] ), .ZN(_04080_ ) );
OR3_X1 _11834_ ( .A1(_03925_ ), .A2(_04080_ ), .A3(_03962_ ), .ZN(_04081_ ) );
BUF_X4 _11835_ ( .A(_03930_ ), .Z(_04082_ ) );
OR2_X1 _11836_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[0][12] ), .ZN(_04083_ ) );
BUF_X4 _11837_ ( .A(_03937_ ), .Z(_04084_ ) );
OAI211_X1 _11838_ ( .A(_04083_ ), .B(_04012_ ), .C1(_04084_ ), .C2(\myreg.Reg[1][12] ), .ZN(_04085_ ) );
OR2_X1 _11839_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[2][12] ), .ZN(_04086_ ) );
OAI211_X1 _11840_ ( .A(_04086_ ), .B(fanout_net_36 ), .C1(_03997_ ), .C2(\myreg.Reg[3][12] ), .ZN(_04087_ ) );
NAND3_X1 _11841_ ( .A1(_04085_ ), .A2(_04087_ ), .A3(_03950_ ), .ZN(_04088_ ) );
MUX2_X1 _11842_ ( .A(\myreg.Reg[6][12] ), .B(\myreg.Reg[7][12] ), .S(fanout_net_29 ), .Z(_04089_ ) );
MUX2_X1 _11843_ ( .A(\myreg.Reg[4][12] ), .B(\myreg.Reg[5][12] ), .S(fanout_net_29 ), .Z(_04090_ ) );
MUX2_X1 _11844_ ( .A(_04089_ ), .B(_04090_ ), .S(_03996_ ), .Z(_04091_ ) );
BUF_X4 _11845_ ( .A(_03950_ ), .Z(_04092_ ) );
OAI211_X1 _11846_ ( .A(_04082_ ), .B(_04088_ ), .C1(_04091_ ), .C2(_04092_ ), .ZN(_04093_ ) );
OR2_X1 _11847_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[14][12] ), .ZN(_04094_ ) );
OAI211_X1 _11848_ ( .A(_04094_ ), .B(fanout_net_36 ), .C1(_03997_ ), .C2(\myreg.Reg[15][12] ), .ZN(_04095_ ) );
OR2_X1 _11849_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[12][12] ), .ZN(_04096_ ) );
OAI211_X1 _11850_ ( .A(_04096_ ), .B(_03996_ ), .C1(_03997_ ), .C2(\myreg.Reg[13][12] ), .ZN(_04097_ ) );
NAND3_X1 _11851_ ( .A1(_04095_ ), .A2(_04097_ ), .A3(fanout_net_38 ), .ZN(_04098_ ) );
MUX2_X1 _11852_ ( .A(\myreg.Reg[8][12] ), .B(\myreg.Reg[9][12] ), .S(fanout_net_29 ), .Z(_04099_ ) );
MUX2_X1 _11853_ ( .A(\myreg.Reg[10][12] ), .B(\myreg.Reg[11][12] ), .S(fanout_net_29 ), .Z(_04100_ ) );
MUX2_X1 _11854_ ( .A(_04099_ ), .B(_04100_ ), .S(fanout_net_36 ), .Z(_04101_ ) );
OAI211_X1 _11855_ ( .A(fanout_net_39 ), .B(_04098_ ), .C1(_04101_ ), .C2(fanout_net_38 ), .ZN(_04102_ ) );
NAND2_X1 _11856_ ( .A1(_04093_ ), .A2(_04102_ ), .ZN(_04103_ ) );
BUF_X2 _11857_ ( .A(_03924_ ), .Z(_04104_ ) );
OAI21_X1 _11858_ ( .A(_04103_ ), .B1(_04104_ ), .B2(_04072_ ), .ZN(_04105_ ) );
AND2_X1 _11859_ ( .A1(_04081_ ), .A2(_04105_ ), .ZN(_04106_ ) );
XNOR2_X2 _11860_ ( .A(_04079_ ), .B(_04106_ ), .ZN(_04107_ ) );
AND2_X1 _11861_ ( .A1(_04078_ ), .A2(_04107_ ), .ZN(_04108_ ) );
INV_X1 _11862_ ( .A(_02694_ ), .ZN(_04109_ ) );
INV_X1 _11863_ ( .A(\EX_LS_result_reg [15] ), .ZN(_04110_ ) );
OR3_X1 _11864_ ( .A1(_03925_ ), .A2(_04110_ ), .A3(_03962_ ), .ZN(_04111_ ) );
OR2_X1 _11865_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[0][15] ), .ZN(_04112_ ) );
OAI211_X1 _11866_ ( .A(_04112_ ), .B(_04005_ ), .C1(_03937_ ), .C2(\myreg.Reg[1][15] ), .ZN(_04113_ ) );
OR2_X1 _11867_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[2][15] ), .ZN(_04114_ ) );
OAI211_X1 _11868_ ( .A(_04114_ ), .B(fanout_net_36 ), .C1(_03937_ ), .C2(\myreg.Reg[3][15] ), .ZN(_04115_ ) );
NAND3_X1 _11869_ ( .A1(_04113_ ), .A2(_04115_ ), .A3(_03943_ ), .ZN(_04116_ ) );
MUX2_X1 _11870_ ( .A(\myreg.Reg[6][15] ), .B(\myreg.Reg[7][15] ), .S(fanout_net_29 ), .Z(_04117_ ) );
MUX2_X1 _11871_ ( .A(\myreg.Reg[4][15] ), .B(\myreg.Reg[5][15] ), .S(fanout_net_29 ), .Z(_04118_ ) );
MUX2_X1 _11872_ ( .A(_04117_ ), .B(_04118_ ), .S(_03934_ ), .Z(_04119_ ) );
OAI211_X1 _11873_ ( .A(_03930_ ), .B(_04116_ ), .C1(_04119_ ), .C2(_03950_ ), .ZN(_04120_ ) );
OR2_X1 _11874_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[14][15] ), .ZN(_04121_ ) );
OAI211_X1 _11875_ ( .A(_04121_ ), .B(fanout_net_36 ), .C1(_03937_ ), .C2(\myreg.Reg[15][15] ), .ZN(_04122_ ) );
OR2_X1 _11876_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[12][15] ), .ZN(_04123_ ) );
OAI211_X1 _11877_ ( .A(_04123_ ), .B(_03934_ ), .C1(_03937_ ), .C2(\myreg.Reg[13][15] ), .ZN(_04124_ ) );
NAND3_X1 _11878_ ( .A1(_04122_ ), .A2(_04124_ ), .A3(fanout_net_38 ), .ZN(_04125_ ) );
MUX2_X1 _11879_ ( .A(\myreg.Reg[8][15] ), .B(\myreg.Reg[9][15] ), .S(fanout_net_29 ), .Z(_04126_ ) );
MUX2_X1 _11880_ ( .A(\myreg.Reg[10][15] ), .B(\myreg.Reg[11][15] ), .S(fanout_net_29 ), .Z(_04127_ ) );
MUX2_X1 _11881_ ( .A(_04126_ ), .B(_04127_ ), .S(fanout_net_36 ), .Z(_04128_ ) );
OAI211_X1 _11882_ ( .A(fanout_net_39 ), .B(_04125_ ), .C1(_04128_ ), .C2(fanout_net_38 ), .ZN(_04129_ ) );
NAND2_X1 _11883_ ( .A1(_04120_ ), .A2(_04129_ ), .ZN(_04130_ ) );
OAI21_X1 _11884_ ( .A(_04130_ ), .B1(_03925_ ), .B2(_03962_ ), .ZN(_04131_ ) );
AND2_X1 _11885_ ( .A1(_04111_ ), .A2(_04131_ ), .ZN(_04132_ ) );
XNOR2_X1 _11886_ ( .A(_04109_ ), .B(_04132_ ), .ZN(_04133_ ) );
INV_X1 _11887_ ( .A(_02717_ ), .ZN(_04134_ ) );
AOI22_X1 _11888_ ( .A1(_02110_ ), .A2(\ID_EX_rs2 [3] ), .B1(_03331_ ), .B2(\EX_LS_dest_reg [1] ), .ZN(_04135_ ) );
NAND3_X1 _11889_ ( .A1(_03918_ ), .A2(_03922_ ), .A3(_04135_ ), .ZN(_04136_ ) );
AOI211_X2 _11890_ ( .A(_03927_ ), .B(_04136_ ), .C1(\EX_LS_dest_reg [3] ), .C2(_03327_ ), .ZN(_04137_ ) );
NAND2_X1 _11891_ ( .A1(_04137_ ), .A2(_02094_ ), .ZN(_04138_ ) );
CLKBUF_X2 _11892_ ( .A(_04138_ ), .Z(_04139_ ) );
OAI221_X1 _11893_ ( .A(_03921_ ), .B1(\EX_LS_dest_reg [1] ), .B2(_03331_ ), .C1(_02096_ ), .C2(_02097_ ), .ZN(_04140_ ) );
CLKBUF_X2 _11894_ ( .A(_04140_ ), .Z(_04141_ ) );
OR3_X1 _11895_ ( .A1(_04139_ ), .A2(\EX_LS_result_reg [14] ), .A3(_04141_ ), .ZN(_04142_ ) );
OR2_X1 _11896_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[4][14] ), .ZN(_04143_ ) );
BUF_X4 _11897_ ( .A(_04005_ ), .Z(_04144_ ) );
BUF_X4 _11898_ ( .A(_04000_ ), .Z(_04145_ ) );
OAI211_X1 _11899_ ( .A(_04143_ ), .B(_04144_ ), .C1(_04145_ ), .C2(\myreg.Reg[5][14] ), .ZN(_04146_ ) );
OR2_X1 _11900_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[6][14] ), .ZN(_04147_ ) );
OAI211_X1 _11901_ ( .A(_04147_ ), .B(fanout_net_36 ), .C1(_04084_ ), .C2(\myreg.Reg[7][14] ), .ZN(_04148_ ) );
NAND3_X1 _11902_ ( .A1(_04146_ ), .A2(_04148_ ), .A3(fanout_net_38 ), .ZN(_04149_ ) );
MUX2_X1 _11903_ ( .A(\myreg.Reg[2][14] ), .B(\myreg.Reg[3][14] ), .S(fanout_net_29 ), .Z(_04150_ ) );
MUX2_X1 _11904_ ( .A(\myreg.Reg[0][14] ), .B(\myreg.Reg[1][14] ), .S(fanout_net_30 ), .Z(_04151_ ) );
MUX2_X1 _11905_ ( .A(_04150_ ), .B(_04151_ ), .S(_04012_ ), .Z(_04152_ ) );
OAI211_X1 _11906_ ( .A(_04082_ ), .B(_04149_ ), .C1(_04152_ ), .C2(fanout_net_38 ), .ZN(_04153_ ) );
NOR2_X1 _11907_ ( .A1(_03997_ ), .A2(\myreg.Reg[11][14] ), .ZN(_04154_ ) );
OAI21_X1 _11908_ ( .A(fanout_net_36 ), .B1(fanout_net_30 ), .B2(\myreg.Reg[10][14] ), .ZN(_04155_ ) );
NOR2_X1 _11909_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[8][14] ), .ZN(_04156_ ) );
OAI21_X1 _11910_ ( .A(_04012_ ), .B1(_04084_ ), .B2(\myreg.Reg[9][14] ), .ZN(_04157_ ) );
OAI221_X1 _11911_ ( .A(_04014_ ), .B1(_04154_ ), .B2(_04155_ ), .C1(_04156_ ), .C2(_04157_ ), .ZN(_04158_ ) );
MUX2_X1 _11912_ ( .A(\myreg.Reg[12][14] ), .B(\myreg.Reg[13][14] ), .S(fanout_net_30 ), .Z(_04159_ ) );
MUX2_X1 _11913_ ( .A(\myreg.Reg[14][14] ), .B(\myreg.Reg[15][14] ), .S(fanout_net_30 ), .Z(_04160_ ) );
MUX2_X1 _11914_ ( .A(_04159_ ), .B(_04160_ ), .S(fanout_net_36 ), .Z(_04161_ ) );
OAI211_X1 _11915_ ( .A(fanout_net_39 ), .B(_04158_ ), .C1(_04161_ ), .C2(_04092_ ), .ZN(_04162_ ) );
OAI211_X1 _11916_ ( .A(_04153_ ), .B(_04162_ ), .C1(_04139_ ), .C2(_04141_ ), .ZN(_04163_ ) );
NAND2_X1 _11917_ ( .A1(_04142_ ), .A2(_04163_ ), .ZN(_04164_ ) );
XNOR2_X1 _11918_ ( .A(_04134_ ), .B(_04164_ ), .ZN(_04165_ ) );
NAND3_X1 _11919_ ( .A1(_04108_ ), .A2(_04133_ ), .A3(_04165_ ), .ZN(_04166_ ) );
NOR2_X1 _11920_ ( .A1(_04050_ ), .A2(_04166_ ), .ZN(_04167_ ) );
OR2_X1 _11921_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[4][6] ), .ZN(_04168_ ) );
OAI211_X1 _11922_ ( .A(_04168_ ), .B(_04005_ ), .C1(_04000_ ), .C2(\myreg.Reg[5][6] ), .ZN(_04169_ ) );
OR2_X1 _11923_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[6][6] ), .ZN(_04170_ ) );
OAI211_X1 _11924_ ( .A(_04170_ ), .B(fanout_net_36 ), .C1(_03937_ ), .C2(\myreg.Reg[7][6] ), .ZN(_04171_ ) );
NAND3_X1 _11925_ ( .A1(_04169_ ), .A2(_04171_ ), .A3(fanout_net_38 ), .ZN(_04172_ ) );
MUX2_X1 _11926_ ( .A(\myreg.Reg[2][6] ), .B(\myreg.Reg[3][6] ), .S(fanout_net_30 ), .Z(_04173_ ) );
MUX2_X1 _11927_ ( .A(\myreg.Reg[0][6] ), .B(\myreg.Reg[1][6] ), .S(fanout_net_30 ), .Z(_04174_ ) );
MUX2_X1 _11928_ ( .A(_04173_ ), .B(_04174_ ), .S(_03934_ ), .Z(_04175_ ) );
OAI211_X1 _11929_ ( .A(_03930_ ), .B(_04172_ ), .C1(_04175_ ), .C2(fanout_net_38 ), .ZN(_04176_ ) );
NOR2_X1 _11930_ ( .A1(_03940_ ), .A2(\myreg.Reg[11][6] ), .ZN(_04177_ ) );
OAI21_X1 _11931_ ( .A(fanout_net_36 ), .B1(fanout_net_30 ), .B2(\myreg.Reg[10][6] ), .ZN(_04178_ ) );
NOR2_X1 _11932_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[8][6] ), .ZN(_04179_ ) );
OAI21_X1 _11933_ ( .A(_03934_ ), .B1(_03940_ ), .B2(\myreg.Reg[9][6] ), .ZN(_04180_ ) );
OAI221_X1 _11934_ ( .A(_03943_ ), .B1(_04177_ ), .B2(_04178_ ), .C1(_04179_ ), .C2(_04180_ ), .ZN(_04181_ ) );
MUX2_X1 _11935_ ( .A(\myreg.Reg[12][6] ), .B(\myreg.Reg[13][6] ), .S(fanout_net_30 ), .Z(_04182_ ) );
MUX2_X1 _11936_ ( .A(\myreg.Reg[14][6] ), .B(\myreg.Reg[15][6] ), .S(fanout_net_30 ), .Z(_04183_ ) );
MUX2_X1 _11937_ ( .A(_04182_ ), .B(_04183_ ), .S(fanout_net_36 ), .Z(_04184_ ) );
OAI211_X1 _11938_ ( .A(fanout_net_39 ), .B(_04181_ ), .C1(_04184_ ), .C2(_03950_ ), .ZN(_04185_ ) );
AOI21_X1 _11939_ ( .A(_03994_ ), .B1(_04176_ ), .B2(_04185_ ), .ZN(_04186_ ) );
AND4_X1 _11940_ ( .A1(\EX_LS_result_reg [6] ), .A2(_02094_ ), .A3(_03989_ ), .A4(_03988_ ), .ZN(_04187_ ) );
NOR2_X1 _11941_ ( .A1(_04186_ ), .A2(_04187_ ), .ZN(_04188_ ) );
INV_X1 _11942_ ( .A(_02565_ ), .ZN(_04189_ ) );
XNOR2_X1 _11943_ ( .A(_04188_ ), .B(_04189_ ), .ZN(_04190_ ) );
NOR2_X1 _11944_ ( .A1(_03966_ ), .A2(\myreg.Reg[11][7] ), .ZN(_04191_ ) );
OAI21_X1 _11945_ ( .A(fanout_net_36 ), .B1(fanout_net_30 ), .B2(\myreg.Reg[10][7] ), .ZN(_04192_ ) );
NOR2_X1 _11946_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[8][7] ), .ZN(_04193_ ) );
OAI21_X1 _11947_ ( .A(_03947_ ), .B1(_03966_ ), .B2(\myreg.Reg[9][7] ), .ZN(_04194_ ) );
OAI221_X1 _11948_ ( .A(_03949_ ), .B1(_04191_ ), .B2(_04192_ ), .C1(_04193_ ), .C2(_04194_ ), .ZN(_04195_ ) );
MUX2_X1 _11949_ ( .A(\myreg.Reg[12][7] ), .B(\myreg.Reg[13][7] ), .S(fanout_net_30 ), .Z(_04196_ ) );
MUX2_X1 _11950_ ( .A(\myreg.Reg[14][7] ), .B(\myreg.Reg[15][7] ), .S(fanout_net_30 ), .Z(_04197_ ) );
MUX2_X1 _11951_ ( .A(_04196_ ), .B(_04197_ ), .S(fanout_net_36 ), .Z(_04198_ ) );
OAI211_X1 _11952_ ( .A(fanout_net_39 ), .B(_04195_ ), .C1(_04198_ ), .C2(_03943_ ), .ZN(_04199_ ) );
OR2_X1 _11953_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[4][7] ), .ZN(_04200_ ) );
OAI211_X1 _11954_ ( .A(_04200_ ), .B(_03947_ ), .C1(_03940_ ), .C2(\myreg.Reg[5][7] ), .ZN(_04201_ ) );
OR2_X1 _11955_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[6][7] ), .ZN(_04202_ ) );
OAI211_X1 _11956_ ( .A(_04202_ ), .B(fanout_net_36 ), .C1(_03966_ ), .C2(\myreg.Reg[7][7] ), .ZN(_04203_ ) );
NAND3_X1 _11957_ ( .A1(_04201_ ), .A2(_04203_ ), .A3(fanout_net_38 ), .ZN(_04204_ ) );
MUX2_X1 _11958_ ( .A(\myreg.Reg[2][7] ), .B(\myreg.Reg[3][7] ), .S(fanout_net_30 ), .Z(_04205_ ) );
MUX2_X1 _11959_ ( .A(\myreg.Reg[0][7] ), .B(\myreg.Reg[1][7] ), .S(fanout_net_30 ), .Z(_04206_ ) );
MUX2_X1 _11960_ ( .A(_04205_ ), .B(_04206_ ), .S(_03947_ ), .Z(_04207_ ) );
OAI211_X1 _11961_ ( .A(_03930_ ), .B(_04204_ ), .C1(_04207_ ), .C2(fanout_net_38 ), .ZN(_04208_ ) );
NAND2_X1 _11962_ ( .A1(_04199_ ), .A2(_04208_ ), .ZN(_04209_ ) );
OAI21_X1 _11963_ ( .A(_04209_ ), .B1(_03925_ ), .B2(_03962_ ), .ZN(_04210_ ) );
NAND4_X1 _11964_ ( .A1(_02094_ ), .A2(\EX_LS_result_reg [7] ), .A3(_03988_ ), .A4(_03989_ ), .ZN(_04211_ ) );
AND2_X1 _11965_ ( .A1(_04210_ ), .A2(_04211_ ), .ZN(_04212_ ) );
XOR2_X1 _11966_ ( .A(_02543_ ), .B(_04212_ ), .Z(_04213_ ) );
AND2_X1 _11967_ ( .A1(_04190_ ), .A2(_04213_ ), .ZN(_04214_ ) );
OR3_X1 _11968_ ( .A1(_04138_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_04140_ ), .ZN(_04215_ ) );
OR2_X1 _11969_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04216_ ) );
OAI211_X1 _11970_ ( .A(_04216_ ), .B(_03947_ ), .C1(_03966_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04217_ ) );
OR2_X1 _11971_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04218_ ) );
OAI211_X1 _11972_ ( .A(_04218_ ), .B(fanout_net_37 ), .C1(_03966_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04219_ ) );
NAND3_X1 _11973_ ( .A1(_04217_ ), .A2(_04219_ ), .A3(fanout_net_38 ), .ZN(_04220_ ) );
MUX2_X1 _11974_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04221_ ) );
MUX2_X1 _11975_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04222_ ) );
MUX2_X1 _11976_ ( .A(_04221_ ), .B(_04222_ ), .S(_03933_ ), .Z(_04223_ ) );
OAI211_X1 _11977_ ( .A(_03929_ ), .B(_04220_ ), .C1(_04223_ ), .C2(fanout_net_38 ), .ZN(_04224_ ) );
NOR2_X1 _11978_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04225_ ) );
OAI21_X1 _11979_ ( .A(_03933_ ), .B1(_03936_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04226_ ) );
MUX2_X1 _11980_ ( .A(_02571_ ), .B(_02572_ ), .S(fanout_net_30 ), .Z(_04227_ ) );
OAI221_X1 _11981_ ( .A(_03949_ ), .B1(_04225_ ), .B2(_04226_ ), .C1(_04227_ ), .C2(_03947_ ), .ZN(_04228_ ) );
MUX2_X1 _11982_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04229_ ) );
MUX2_X1 _11983_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04230_ ) );
MUX2_X1 _11984_ ( .A(_04229_ ), .B(_04230_ ), .S(fanout_net_37 ), .Z(_04231_ ) );
OAI211_X1 _11985_ ( .A(fanout_net_39 ), .B(_04228_ ), .C1(_04231_ ), .C2(_03943_ ), .ZN(_04232_ ) );
OAI211_X1 _11986_ ( .A(_04224_ ), .B(_04232_ ), .C1(_04138_ ), .C2(_04140_ ), .ZN(_04233_ ) );
NAND2_X1 _11987_ ( .A1(_04215_ ), .A2(_04233_ ), .ZN(_04234_ ) );
XNOR2_X2 _11988_ ( .A(_04234_ ), .B(_02589_ ), .ZN(_04235_ ) );
INV_X1 _11989_ ( .A(_02464_ ), .ZN(_04236_ ) );
OR2_X1 _11990_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[8][1] ), .ZN(_04237_ ) );
OAI211_X1 _11991_ ( .A(_04237_ ), .B(_03933_ ), .C1(_03936_ ), .C2(\myreg.Reg[9][1] ), .ZN(_04238_ ) );
OR2_X1 _11992_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[10][1] ), .ZN(_04239_ ) );
OAI211_X1 _11993_ ( .A(_04239_ ), .B(fanout_net_37 ), .C1(_03936_ ), .C2(\myreg.Reg[11][1] ), .ZN(_04240_ ) );
NAND3_X1 _11994_ ( .A1(_04238_ ), .A2(_04240_ ), .A3(_03942_ ), .ZN(_04241_ ) );
MUX2_X1 _11995_ ( .A(\myreg.Reg[14][1] ), .B(\myreg.Reg[15][1] ), .S(fanout_net_31 ), .Z(_04242_ ) );
MUX2_X1 _11996_ ( .A(\myreg.Reg[12][1] ), .B(\myreg.Reg[13][1] ), .S(fanout_net_31 ), .Z(_04243_ ) );
MUX2_X1 _11997_ ( .A(_04242_ ), .B(_04243_ ), .S(_03933_ ), .Z(_04244_ ) );
OAI211_X1 _11998_ ( .A(fanout_net_39 ), .B(_04241_ ), .C1(_04244_ ), .C2(_03949_ ), .ZN(_04245_ ) );
MUX2_X1 _11999_ ( .A(\myreg.Reg[0][1] ), .B(\myreg.Reg[1][1] ), .S(fanout_net_31 ), .Z(_04246_ ) );
AND2_X1 _12000_ ( .A1(_04246_ ), .A2(_03932_ ), .ZN(_04247_ ) );
MUX2_X1 _12001_ ( .A(\myreg.Reg[2][1] ), .B(\myreg.Reg[3][1] ), .S(fanout_net_31 ), .Z(_04248_ ) );
AOI211_X1 _12002_ ( .A(fanout_net_38 ), .B(_04247_ ), .C1(fanout_net_37 ), .C2(_04248_ ), .ZN(_04249_ ) );
MUX2_X1 _12003_ ( .A(\myreg.Reg[6][1] ), .B(\myreg.Reg[7][1] ), .S(fanout_net_31 ), .Z(_04250_ ) );
MUX2_X1 _12004_ ( .A(\myreg.Reg[4][1] ), .B(\myreg.Reg[5][1] ), .S(fanout_net_31 ), .Z(_04251_ ) );
MUX2_X1 _12005_ ( .A(_04250_ ), .B(_04251_ ), .S(_03932_ ), .Z(_04252_ ) );
OAI21_X1 _12006_ ( .A(_03929_ ), .B1(_04252_ ), .B2(_03949_ ), .ZN(_04253_ ) );
OAI221_X1 _12007_ ( .A(_04245_ ), .B1(_04249_ ), .B2(_04253_ ), .C1(_04138_ ), .C2(_04140_ ), .ZN(_04254_ ) );
OR3_X2 _12008_ ( .A1(_04138_ ), .A2(\EX_LS_result_reg [1] ), .A3(_04140_ ), .ZN(_04255_ ) );
NAND2_X2 _12009_ ( .A1(_04254_ ), .A2(_04255_ ), .ZN(_04256_ ) );
XNOR2_X2 _12010_ ( .A(_04236_ ), .B(_04256_ ), .ZN(_04257_ ) );
INV_X1 _12011_ ( .A(_02611_ ), .ZN(_04258_ ) );
NAND2_X1 _12012_ ( .A1(_03994_ ), .A2(\EX_LS_result_reg [4] ), .ZN(_04259_ ) );
OR2_X1 _12013_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[0][4] ), .ZN(_04260_ ) );
OAI211_X1 _12014_ ( .A(_04260_ ), .B(_04012_ ), .C1(_04084_ ), .C2(\myreg.Reg[1][4] ), .ZN(_04261_ ) );
OR2_X1 _12015_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[2][4] ), .ZN(_04262_ ) );
OAI211_X1 _12016_ ( .A(_04262_ ), .B(fanout_net_37 ), .C1(_03997_ ), .C2(\myreg.Reg[3][4] ), .ZN(_04263_ ) );
NAND3_X1 _12017_ ( .A1(_04261_ ), .A2(_04263_ ), .A3(_03950_ ), .ZN(_04264_ ) );
MUX2_X1 _12018_ ( .A(\myreg.Reg[6][4] ), .B(\myreg.Reg[7][4] ), .S(fanout_net_31 ), .Z(_04265_ ) );
MUX2_X1 _12019_ ( .A(\myreg.Reg[4][4] ), .B(\myreg.Reg[5][4] ), .S(fanout_net_31 ), .Z(_04266_ ) );
MUX2_X1 _12020_ ( .A(_04265_ ), .B(_04266_ ), .S(_03996_ ), .Z(_04267_ ) );
OAI211_X1 _12021_ ( .A(_04082_ ), .B(_04264_ ), .C1(_04267_ ), .C2(_04092_ ), .ZN(_04268_ ) );
OR2_X1 _12022_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[14][4] ), .ZN(_04269_ ) );
OAI211_X1 _12023_ ( .A(_04269_ ), .B(fanout_net_37 ), .C1(_03997_ ), .C2(\myreg.Reg[15][4] ), .ZN(_04270_ ) );
OR2_X1 _12024_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[12][4] ), .ZN(_04271_ ) );
OAI211_X1 _12025_ ( .A(_04271_ ), .B(_04012_ ), .C1(_03997_ ), .C2(\myreg.Reg[13][4] ), .ZN(_04272_ ) );
NAND3_X1 _12026_ ( .A1(_04270_ ), .A2(_04272_ ), .A3(fanout_net_38 ), .ZN(_04273_ ) );
MUX2_X1 _12027_ ( .A(\myreg.Reg[8][4] ), .B(\myreg.Reg[9][4] ), .S(fanout_net_31 ), .Z(_04274_ ) );
MUX2_X1 _12028_ ( .A(\myreg.Reg[10][4] ), .B(\myreg.Reg[11][4] ), .S(fanout_net_31 ), .Z(_04275_ ) );
MUX2_X1 _12029_ ( .A(_04274_ ), .B(_04275_ ), .S(fanout_net_37 ), .Z(_04276_ ) );
OAI211_X1 _12030_ ( .A(fanout_net_39 ), .B(_04273_ ), .C1(_04276_ ), .C2(fanout_net_38 ), .ZN(_04277_ ) );
NAND2_X1 _12031_ ( .A1(_04268_ ), .A2(_04277_ ), .ZN(_04278_ ) );
OAI21_X1 _12032_ ( .A(_04278_ ), .B1(_04104_ ), .B2(_04072_ ), .ZN(_04279_ ) );
AND2_X1 _12033_ ( .A1(_04259_ ), .A2(_04279_ ), .ZN(_04280_ ) );
XNOR2_X1 _12034_ ( .A(_04258_ ), .B(_04280_ ), .ZN(_04281_ ) );
OR2_X1 _12035_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[0][2] ), .ZN(_04282_ ) );
OAI211_X1 _12036_ ( .A(_04282_ ), .B(_04005_ ), .C1(_03937_ ), .C2(\myreg.Reg[1][2] ), .ZN(_04283_ ) );
OR2_X1 _12037_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[2][2] ), .ZN(_04284_ ) );
OAI211_X1 _12038_ ( .A(_04284_ ), .B(fanout_net_37 ), .C1(_03940_ ), .C2(\myreg.Reg[3][2] ), .ZN(_04285_ ) );
NAND3_X1 _12039_ ( .A1(_04283_ ), .A2(_04285_ ), .A3(_03943_ ), .ZN(_04286_ ) );
MUX2_X1 _12040_ ( .A(\myreg.Reg[6][2] ), .B(\myreg.Reg[7][2] ), .S(fanout_net_31 ), .Z(_04287_ ) );
MUX2_X1 _12041_ ( .A(\myreg.Reg[4][2] ), .B(\myreg.Reg[5][2] ), .S(fanout_net_31 ), .Z(_04288_ ) );
MUX2_X1 _12042_ ( .A(_04287_ ), .B(_04288_ ), .S(_03934_ ), .Z(_04289_ ) );
OAI211_X1 _12043_ ( .A(_03930_ ), .B(_04286_ ), .C1(_04289_ ), .C2(_03950_ ), .ZN(_04290_ ) );
OR2_X1 _12044_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[14][2] ), .ZN(_04291_ ) );
OAI211_X1 _12045_ ( .A(_04291_ ), .B(fanout_net_37 ), .C1(_03937_ ), .C2(\myreg.Reg[15][2] ), .ZN(_04292_ ) );
OR2_X1 _12046_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[12][2] ), .ZN(_04293_ ) );
OAI211_X1 _12047_ ( .A(_04293_ ), .B(_03934_ ), .C1(_03940_ ), .C2(\myreg.Reg[13][2] ), .ZN(_04294_ ) );
NAND3_X1 _12048_ ( .A1(_04292_ ), .A2(_04294_ ), .A3(fanout_net_38 ), .ZN(_04295_ ) );
MUX2_X1 _12049_ ( .A(\myreg.Reg[8][2] ), .B(\myreg.Reg[9][2] ), .S(fanout_net_31 ), .Z(_04296_ ) );
MUX2_X1 _12050_ ( .A(\myreg.Reg[10][2] ), .B(\myreg.Reg[11][2] ), .S(fanout_net_31 ), .Z(_04297_ ) );
MUX2_X1 _12051_ ( .A(_04296_ ), .B(_04297_ ), .S(fanout_net_37 ), .Z(_04298_ ) );
OAI211_X1 _12052_ ( .A(fanout_net_39 ), .B(_04295_ ), .C1(_04298_ ), .C2(fanout_net_38 ), .ZN(_04299_ ) );
NAND2_X1 _12053_ ( .A1(_04290_ ), .A2(_04299_ ), .ZN(_04300_ ) );
OAI21_X1 _12054_ ( .A(_04300_ ), .B1(_03925_ ), .B2(_03962_ ), .ZN(_04301_ ) );
INV_X1 _12055_ ( .A(\EX_LS_result_reg [2] ), .ZN(_04302_ ) );
OR3_X1 _12056_ ( .A1(_03924_ ), .A2(_04302_ ), .A3(_03927_ ), .ZN(_04303_ ) );
AND3_X1 _12057_ ( .A1(_02441_ ), .A2(_04301_ ), .A3(_04303_ ), .ZN(_04304_ ) );
AOI21_X1 _12058_ ( .A(_02441_ ), .B1(_04301_ ), .B2(_04303_ ), .ZN(_04305_ ) );
NOR2_X4 _12059_ ( .A1(_04304_ ), .A2(_04305_ ), .ZN(_04306_ ) );
NAND3_X1 _12060_ ( .A1(_04257_ ), .A2(_04281_ ), .A3(_04306_ ), .ZN(_04307_ ) );
OR3_X1 _12061_ ( .A1(_04139_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_04141_ ), .ZN(_04308_ ) );
OR2_X1 _12062_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04309_ ) );
OAI211_X1 _12063_ ( .A(_04309_ ), .B(_04012_ ), .C1(_04084_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04310_ ) );
OR2_X1 _12064_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04311_ ) );
OAI211_X1 _12065_ ( .A(_04311_ ), .B(fanout_net_37 ), .C1(_04084_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04312_ ) );
NAND3_X1 _12066_ ( .A1(_04310_ ), .A2(_04312_ ), .A3(_04014_ ), .ZN(_04313_ ) );
MUX2_X1 _12067_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04314_ ) );
MUX2_X1 _12068_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04315_ ) );
MUX2_X1 _12069_ ( .A(_04314_ ), .B(_04315_ ), .S(_03996_ ), .Z(_04316_ ) );
OAI211_X1 _12070_ ( .A(fanout_net_39 ), .B(_04313_ ), .C1(_04316_ ), .C2(_04092_ ), .ZN(_04317_ ) );
OR2_X1 _12071_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04318_ ) );
OAI211_X1 _12072_ ( .A(_04318_ ), .B(_04012_ ), .C1(_04084_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04319_ ) );
OR2_X1 _12073_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04320_ ) );
OAI211_X1 _12074_ ( .A(_04320_ ), .B(fanout_net_37 ), .C1(_03997_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04321_ ) );
NAND3_X1 _12075_ ( .A1(_04319_ ), .A2(_04321_ ), .A3(_04014_ ), .ZN(_04322_ ) );
MUX2_X1 _12076_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04323_ ) );
MUX2_X1 _12077_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04324_ ) );
MUX2_X1 _12078_ ( .A(_04323_ ), .B(_04324_ ), .S(_03996_ ), .Z(_04325_ ) );
OAI211_X1 _12079_ ( .A(_04082_ ), .B(_04322_ ), .C1(_04325_ ), .C2(_04092_ ), .ZN(_04326_ ) );
OAI211_X1 _12080_ ( .A(_04317_ ), .B(_04326_ ), .C1(_04139_ ), .C2(_04141_ ), .ZN(_04327_ ) );
NAND2_X1 _12081_ ( .A1(_04308_ ), .A2(_04327_ ), .ZN(_04328_ ) );
XNOR2_X1 _12082_ ( .A(_04328_ ), .B(_02516_ ), .ZN(_04329_ ) );
INV_X1 _12083_ ( .A(_04329_ ), .ZN(_04330_ ) );
AND2_X2 _12084_ ( .A1(_02468_ ), .A2(_02488_ ), .ZN(_04331_ ) );
OR2_X1 _12085_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[0][0] ), .ZN(_04332_ ) );
OAI211_X1 _12086_ ( .A(_04332_ ), .B(_03933_ ), .C1(_03936_ ), .C2(\myreg.Reg[1][0] ), .ZN(_04333_ ) );
NOR2_X1 _12087_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[2][0] ), .ZN(_04334_ ) );
OAI21_X1 _12088_ ( .A(fanout_net_37 ), .B1(_03936_ ), .B2(\myreg.Reg[3][0] ), .ZN(_04335_ ) );
OAI211_X1 _12089_ ( .A(_04333_ ), .B(_03949_ ), .C1(_04334_ ), .C2(_04335_ ), .ZN(_04336_ ) );
MUX2_X1 _12090_ ( .A(\myreg.Reg[6][0] ), .B(\myreg.Reg[7][0] ), .S(fanout_net_32 ), .Z(_04337_ ) );
MUX2_X1 _12091_ ( .A(\myreg.Reg[4][0] ), .B(\myreg.Reg[5][0] ), .S(fanout_net_32 ), .Z(_04338_ ) );
MUX2_X1 _12092_ ( .A(_04337_ ), .B(_04338_ ), .S(_03933_ ), .Z(_04339_ ) );
OAI211_X1 _12093_ ( .A(_03929_ ), .B(_04336_ ), .C1(_04339_ ), .C2(_03949_ ), .ZN(_04340_ ) );
OR2_X1 _12094_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[8][0] ), .ZN(_04341_ ) );
OAI211_X1 _12095_ ( .A(_04341_ ), .B(_03933_ ), .C1(_03936_ ), .C2(\myreg.Reg[9][0] ), .ZN(_04342_ ) );
OR2_X1 _12096_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[10][0] ), .ZN(_04343_ ) );
OAI211_X1 _12097_ ( .A(_04343_ ), .B(fanout_net_37 ), .C1(_03936_ ), .C2(\myreg.Reg[11][0] ), .ZN(_04344_ ) );
NAND3_X1 _12098_ ( .A1(_04342_ ), .A2(_04344_ ), .A3(_03949_ ), .ZN(_04345_ ) );
MUX2_X1 _12099_ ( .A(\myreg.Reg[14][0] ), .B(\myreg.Reg[15][0] ), .S(fanout_net_32 ), .Z(_04346_ ) );
MUX2_X1 _12100_ ( .A(\myreg.Reg[12][0] ), .B(\myreg.Reg[13][0] ), .S(fanout_net_32 ), .Z(_04347_ ) );
MUX2_X1 _12101_ ( .A(_04346_ ), .B(_04347_ ), .S(_03933_ ), .Z(_04348_ ) );
OAI211_X1 _12102_ ( .A(fanout_net_39 ), .B(_04345_ ), .C1(_04348_ ), .C2(_03949_ ), .ZN(_04349_ ) );
NAND2_X1 _12103_ ( .A1(_04340_ ), .A2(_04349_ ), .ZN(_04350_ ) );
OAI21_X1 _12104_ ( .A(_04350_ ), .B1(_03924_ ), .B2(_03927_ ), .ZN(_04351_ ) );
NAND4_X1 _12105_ ( .A1(_02094_ ), .A2(\EX_LS_result_reg [0] ), .A3(_03988_ ), .A4(_03989_ ), .ZN(_04352_ ) );
AND2_X1 _12106_ ( .A1(_04351_ ), .A2(_04352_ ), .ZN(_04353_ ) );
XNOR2_X1 _12107_ ( .A(_04331_ ), .B(_04353_ ), .ZN(_04354_ ) );
NOR3_X1 _12108_ ( .A1(_04307_ ), .A2(_04330_ ), .A3(_04354_ ), .ZN(_04355_ ) );
AND4_X1 _12109_ ( .A1(_04167_ ), .A2(_04214_ ), .A3(_04235_ ), .A4(_04355_ ), .ZN(_04356_ ) );
INV_X1 _12110_ ( .A(_02346_ ), .ZN(_04357_ ) );
OR3_X1 _12111_ ( .A1(_04139_ ), .A2(\EX_LS_result_reg [18] ), .A3(_04141_ ), .ZN(_04358_ ) );
OR2_X1 _12112_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[0][18] ), .ZN(_04359_ ) );
BUF_X4 _12113_ ( .A(_04144_ ), .Z(_04360_ ) );
BUF_X4 _12114_ ( .A(_04145_ ), .Z(_04361_ ) );
OAI211_X1 _12115_ ( .A(_04359_ ), .B(_04360_ ), .C1(_04361_ ), .C2(\myreg.Reg[1][18] ), .ZN(_04362_ ) );
OR2_X1 _12116_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[2][18] ), .ZN(_04363_ ) );
OAI211_X1 _12117_ ( .A(_04363_ ), .B(fanout_net_37 ), .C1(_04145_ ), .C2(\myreg.Reg[3][18] ), .ZN(_04364_ ) );
NAND3_X1 _12118_ ( .A1(_04362_ ), .A2(_04364_ ), .A3(_04092_ ), .ZN(_04365_ ) );
MUX2_X1 _12119_ ( .A(\myreg.Reg[6][18] ), .B(\myreg.Reg[7][18] ), .S(fanout_net_32 ), .Z(_04366_ ) );
MUX2_X1 _12120_ ( .A(\myreg.Reg[4][18] ), .B(\myreg.Reg[5][18] ), .S(fanout_net_32 ), .Z(_04367_ ) );
MUX2_X1 _12121_ ( .A(_04366_ ), .B(_04367_ ), .S(_04144_ ), .Z(_04368_ ) );
BUF_X4 _12122_ ( .A(_04014_ ), .Z(_04369_ ) );
OAI211_X1 _12123_ ( .A(_04082_ ), .B(_04365_ ), .C1(_04368_ ), .C2(_04369_ ), .ZN(_04370_ ) );
OR2_X1 _12124_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[14][18] ), .ZN(_04371_ ) );
OAI211_X1 _12125_ ( .A(_04371_ ), .B(fanout_net_37 ), .C1(_04361_ ), .C2(\myreg.Reg[15][18] ), .ZN(_04372_ ) );
OR2_X1 _12126_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[12][18] ), .ZN(_04373_ ) );
OAI211_X1 _12127_ ( .A(_04373_ ), .B(_04144_ ), .C1(_04145_ ), .C2(\myreg.Reg[13][18] ), .ZN(_04374_ ) );
NAND3_X1 _12128_ ( .A1(_04372_ ), .A2(_04374_ ), .A3(fanout_net_38 ), .ZN(_04375_ ) );
MUX2_X1 _12129_ ( .A(\myreg.Reg[8][18] ), .B(\myreg.Reg[9][18] ), .S(fanout_net_32 ), .Z(_04376_ ) );
MUX2_X1 _12130_ ( .A(\myreg.Reg[10][18] ), .B(\myreg.Reg[11][18] ), .S(fanout_net_32 ), .Z(_04377_ ) );
MUX2_X1 _12131_ ( .A(_04376_ ), .B(_04377_ ), .S(fanout_net_37 ), .Z(_04378_ ) );
OAI211_X1 _12132_ ( .A(fanout_net_39 ), .B(_04375_ ), .C1(_04378_ ), .C2(fanout_net_38 ), .ZN(_04379_ ) );
OAI211_X1 _12133_ ( .A(_04370_ ), .B(_04379_ ), .C1(_04139_ ), .C2(_04141_ ), .ZN(_04380_ ) );
NAND2_X1 _12134_ ( .A1(_04358_ ), .A2(_04380_ ), .ZN(_04381_ ) );
XNOR2_X1 _12135_ ( .A(_04357_ ), .B(_04381_ ), .ZN(_04382_ ) );
INV_X2 _12136_ ( .A(_02370_ ), .ZN(_04383_ ) );
INV_X1 _12137_ ( .A(\EX_LS_result_reg [19] ), .ZN(_04384_ ) );
OR3_X1 _12138_ ( .A1(_04104_ ), .A2(_04384_ ), .A3(_03962_ ), .ZN(_04385_ ) );
OR2_X1 _12139_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[8][19] ), .ZN(_04386_ ) );
OAI211_X1 _12140_ ( .A(_04386_ ), .B(_04012_ ), .C1(_04084_ ), .C2(\myreg.Reg[9][19] ), .ZN(_04387_ ) );
OR2_X1 _12141_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[10][19] ), .ZN(_04388_ ) );
OAI211_X1 _12142_ ( .A(_04388_ ), .B(fanout_net_37 ), .C1(_04084_ ), .C2(\myreg.Reg[11][19] ), .ZN(_04389_ ) );
NAND3_X1 _12143_ ( .A1(_04387_ ), .A2(_04389_ ), .A3(_04014_ ), .ZN(_04390_ ) );
MUX2_X1 _12144_ ( .A(\myreg.Reg[14][19] ), .B(\myreg.Reg[15][19] ), .S(fanout_net_32 ), .Z(_04391_ ) );
MUX2_X1 _12145_ ( .A(\myreg.Reg[12][19] ), .B(\myreg.Reg[13][19] ), .S(fanout_net_32 ), .Z(_04392_ ) );
MUX2_X1 _12146_ ( .A(_04391_ ), .B(_04392_ ), .S(_03996_ ), .Z(_04393_ ) );
OAI211_X1 _12147_ ( .A(fanout_net_39 ), .B(_04390_ ), .C1(_04393_ ), .C2(_04092_ ), .ZN(_04394_ ) );
MUX2_X1 _12148_ ( .A(\myreg.Reg[0][19] ), .B(\myreg.Reg[1][19] ), .S(fanout_net_32 ), .Z(_04395_ ) );
AND2_X1 _12149_ ( .A1(_04395_ ), .A2(_04012_ ), .ZN(_04396_ ) );
MUX2_X1 _12150_ ( .A(\myreg.Reg[2][19] ), .B(\myreg.Reg[3][19] ), .S(fanout_net_32 ), .Z(_04397_ ) );
AOI211_X1 _12151_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_04396_ ), .C1(fanout_net_37 ), .C2(_04397_ ), .ZN(_04398_ ) );
MUX2_X1 _12152_ ( .A(\myreg.Reg[6][19] ), .B(\myreg.Reg[7][19] ), .S(fanout_net_32 ), .Z(_04399_ ) );
MUX2_X1 _12153_ ( .A(\myreg.Reg[4][19] ), .B(\myreg.Reg[5][19] ), .S(fanout_net_32 ), .Z(_04400_ ) );
MUX2_X1 _12154_ ( .A(_04399_ ), .B(_04400_ ), .S(_03996_ ), .Z(_04401_ ) );
OAI21_X1 _12155_ ( .A(_04082_ ), .B1(_04401_ ), .B2(_04092_ ), .ZN(_04402_ ) );
OAI21_X1 _12156_ ( .A(_04394_ ), .B1(_04398_ ), .B2(_04402_ ), .ZN(_04403_ ) );
OAI21_X1 _12157_ ( .A(_04403_ ), .B1(_04072_ ), .B2(_04104_ ), .ZN(_04404_ ) );
AND2_X1 _12158_ ( .A1(_04385_ ), .A2(_04404_ ), .ZN(_04405_ ) );
XNOR2_X1 _12159_ ( .A(_04383_ ), .B(_04405_ ), .ZN(_04406_ ) );
AND2_X1 _12160_ ( .A1(_04382_ ), .A2(_04406_ ), .ZN(_04407_ ) );
OR2_X1 _12161_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[0][17] ), .ZN(_04408_ ) );
OAI211_X1 _12162_ ( .A(_04408_ ), .B(_04360_ ), .C1(_04361_ ), .C2(\myreg.Reg[1][17] ), .ZN(_04409_ ) );
OR2_X1 _12163_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[2][17] ), .ZN(_04410_ ) );
OAI211_X1 _12164_ ( .A(_04410_ ), .B(fanout_net_37 ), .C1(_04361_ ), .C2(\myreg.Reg[3][17] ), .ZN(_04411_ ) );
NAND3_X1 _12165_ ( .A1(_04409_ ), .A2(_04411_ ), .A3(_04092_ ), .ZN(_04412_ ) );
MUX2_X1 _12166_ ( .A(\myreg.Reg[6][17] ), .B(\myreg.Reg[7][17] ), .S(fanout_net_32 ), .Z(_04413_ ) );
MUX2_X1 _12167_ ( .A(\myreg.Reg[4][17] ), .B(\myreg.Reg[5][17] ), .S(fanout_net_32 ), .Z(_04414_ ) );
MUX2_X1 _12168_ ( .A(_04413_ ), .B(_04414_ ), .S(_04144_ ), .Z(_04415_ ) );
OAI211_X1 _12169_ ( .A(_04082_ ), .B(_04412_ ), .C1(_04415_ ), .C2(_04369_ ), .ZN(_04416_ ) );
OR2_X1 _12170_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[14][17] ), .ZN(_04417_ ) );
OAI211_X1 _12171_ ( .A(_04417_ ), .B(fanout_net_37 ), .C1(_04361_ ), .C2(\myreg.Reg[15][17] ), .ZN(_04418_ ) );
OR2_X1 _12172_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[12][17] ), .ZN(_04419_ ) );
OAI211_X1 _12173_ ( .A(_04419_ ), .B(_04144_ ), .C1(_04145_ ), .C2(\myreg.Reg[13][17] ), .ZN(_04420_ ) );
NAND3_X1 _12174_ ( .A1(_04418_ ), .A2(_04420_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04421_ ) );
MUX2_X1 _12175_ ( .A(\myreg.Reg[8][17] ), .B(\myreg.Reg[9][17] ), .S(fanout_net_33 ), .Z(_04422_ ) );
MUX2_X1 _12176_ ( .A(\myreg.Reg[10][17] ), .B(\myreg.Reg[11][17] ), .S(fanout_net_33 ), .Z(_04423_ ) );
MUX2_X1 _12177_ ( .A(_04422_ ), .B(_04423_ ), .S(fanout_net_37 ), .Z(_04424_ ) );
OAI211_X1 _12178_ ( .A(fanout_net_39 ), .B(_04421_ ), .C1(_04424_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04425_ ) );
AOI21_X1 _12179_ ( .A(_03994_ ), .B1(_04416_ ), .B2(_04425_ ), .ZN(_04426_ ) );
INV_X1 _12180_ ( .A(\EX_LS_result_reg [17] ), .ZN(_04427_ ) );
NOR3_X1 _12181_ ( .A1(_04104_ ), .A2(_04427_ ), .A3(_04072_ ), .ZN(_04428_ ) );
NOR2_X1 _12182_ ( .A1(_04426_ ), .A2(_04428_ ), .ZN(_04429_ ) );
INV_X4 _12183_ ( .A(_02394_ ), .ZN(_04430_ ) );
XNOR2_X2 _12184_ ( .A(_04429_ ), .B(_04430_ ), .ZN(_04431_ ) );
INV_X1 _12185_ ( .A(_02417_ ), .ZN(_04432_ ) );
OR3_X1 _12186_ ( .A1(_04139_ ), .A2(\EX_LS_result_reg [16] ), .A3(_04141_ ), .ZN(_04433_ ) );
BUF_X4 _12187_ ( .A(_04082_ ), .Z(_04434_ ) );
OR2_X1 _12188_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[0][16] ), .ZN(_04435_ ) );
BUF_X4 _12189_ ( .A(_04144_ ), .Z(_04436_ ) );
BUF_X4 _12190_ ( .A(_04145_ ), .Z(_04437_ ) );
OAI211_X1 _12191_ ( .A(_04435_ ), .B(_04436_ ), .C1(_04437_ ), .C2(\myreg.Reg[1][16] ), .ZN(_04438_ ) );
OR2_X1 _12192_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[2][16] ), .ZN(_04439_ ) );
OAI211_X1 _12193_ ( .A(_04439_ ), .B(fanout_net_37 ), .C1(_04437_ ), .C2(\myreg.Reg[3][16] ), .ZN(_04440_ ) );
NAND3_X1 _12194_ ( .A1(_04438_ ), .A2(_04440_ ), .A3(_04369_ ), .ZN(_04441_ ) );
MUX2_X1 _12195_ ( .A(\myreg.Reg[6][16] ), .B(\myreg.Reg[7][16] ), .S(fanout_net_33 ), .Z(_04442_ ) );
MUX2_X1 _12196_ ( .A(\myreg.Reg[4][16] ), .B(\myreg.Reg[5][16] ), .S(fanout_net_33 ), .Z(_04443_ ) );
MUX2_X1 _12197_ ( .A(_04442_ ), .B(_04443_ ), .S(_04360_ ), .Z(_04444_ ) );
BUF_X4 _12198_ ( .A(_04369_ ), .Z(_04445_ ) );
OAI211_X1 _12199_ ( .A(_04434_ ), .B(_04441_ ), .C1(_04444_ ), .C2(_04445_ ), .ZN(_04446_ ) );
OR2_X1 _12200_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[14][16] ), .ZN(_04447_ ) );
OAI211_X1 _12201_ ( .A(_04447_ ), .B(fanout_net_37 ), .C1(_04437_ ), .C2(\myreg.Reg[15][16] ), .ZN(_04448_ ) );
OR2_X1 _12202_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[12][16] ), .ZN(_04449_ ) );
OAI211_X1 _12203_ ( .A(_04449_ ), .B(_04360_ ), .C1(_04437_ ), .C2(\myreg.Reg[13][16] ), .ZN(_04450_ ) );
NAND3_X1 _12204_ ( .A1(_04448_ ), .A2(_04450_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04451_ ) );
MUX2_X1 _12205_ ( .A(\myreg.Reg[8][16] ), .B(\myreg.Reg[9][16] ), .S(fanout_net_33 ), .Z(_04452_ ) );
MUX2_X1 _12206_ ( .A(\myreg.Reg[10][16] ), .B(\myreg.Reg[11][16] ), .S(fanout_net_33 ), .Z(_04453_ ) );
MUX2_X1 _12207_ ( .A(_04452_ ), .B(_04453_ ), .S(fanout_net_37 ), .Z(_04454_ ) );
OAI211_X1 _12208_ ( .A(fanout_net_39 ), .B(_04451_ ), .C1(_04454_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04455_ ) );
CLKBUF_X2 _12209_ ( .A(_04139_ ), .Z(_04456_ ) );
BUF_X2 _12210_ ( .A(_04141_ ), .Z(_04457_ ) );
OAI211_X1 _12211_ ( .A(_04446_ ), .B(_04455_ ), .C1(_04456_ ), .C2(_04457_ ), .ZN(_04458_ ) );
NAND2_X1 _12212_ ( .A1(_04433_ ), .A2(_04458_ ), .ZN(_04459_ ) );
XNOR2_X1 _12213_ ( .A(_04432_ ), .B(_04459_ ), .ZN(_04460_ ) );
AND3_X1 _12214_ ( .A1(_04407_ ), .A2(_04431_ ), .A3(_04460_ ), .ZN(_04461_ ) );
INV_X1 _12215_ ( .A(_04461_ ), .ZN(_04462_ ) );
OR3_X1 _12216_ ( .A1(_04456_ ), .A2(\EX_LS_result_reg [20] ), .A3(_04141_ ), .ZN(_04463_ ) );
OR2_X1 _12217_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[0][20] ), .ZN(_04464_ ) );
BUF_X4 _12218_ ( .A(_04360_ ), .Z(_04465_ ) );
BUF_X4 _12219_ ( .A(_04361_ ), .Z(_04466_ ) );
OAI211_X1 _12220_ ( .A(_04464_ ), .B(_04465_ ), .C1(_04466_ ), .C2(\myreg.Reg[1][20] ), .ZN(_04467_ ) );
OR2_X1 _12221_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[2][20] ), .ZN(_04468_ ) );
BUF_X4 _12222_ ( .A(_04145_ ), .Z(_04469_ ) );
OAI211_X1 _12223_ ( .A(_04468_ ), .B(fanout_net_37 ), .C1(_04469_ ), .C2(\myreg.Reg[3][20] ), .ZN(_04470_ ) );
NAND3_X1 _12224_ ( .A1(_04467_ ), .A2(_04470_ ), .A3(_04445_ ), .ZN(_04471_ ) );
MUX2_X1 _12225_ ( .A(\myreg.Reg[6][20] ), .B(\myreg.Reg[7][20] ), .S(fanout_net_33 ), .Z(_04472_ ) );
MUX2_X1 _12226_ ( .A(\myreg.Reg[4][20] ), .B(\myreg.Reg[5][20] ), .S(fanout_net_33 ), .Z(_04473_ ) );
MUX2_X1 _12227_ ( .A(_04472_ ), .B(_04473_ ), .S(_04436_ ), .Z(_04474_ ) );
BUF_X4 _12228_ ( .A(_04369_ ), .Z(_04475_ ) );
OAI211_X1 _12229_ ( .A(_04434_ ), .B(_04471_ ), .C1(_04474_ ), .C2(_04475_ ), .ZN(_04476_ ) );
OR2_X1 _12230_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[14][20] ), .ZN(_04477_ ) );
OAI211_X1 _12231_ ( .A(_04477_ ), .B(fanout_net_37 ), .C1(_04469_ ), .C2(\myreg.Reg[15][20] ), .ZN(_04478_ ) );
OR2_X1 _12232_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[12][20] ), .ZN(_04479_ ) );
OAI211_X1 _12233_ ( .A(_04479_ ), .B(_04436_ ), .C1(_04469_ ), .C2(\myreg.Reg[13][20] ), .ZN(_04480_ ) );
NAND3_X1 _12234_ ( .A1(_04478_ ), .A2(_04480_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04481_ ) );
MUX2_X1 _12235_ ( .A(\myreg.Reg[8][20] ), .B(\myreg.Reg[9][20] ), .S(fanout_net_33 ), .Z(_04482_ ) );
MUX2_X1 _12236_ ( .A(\myreg.Reg[10][20] ), .B(\myreg.Reg[11][20] ), .S(fanout_net_33 ), .Z(_04483_ ) );
MUX2_X1 _12237_ ( .A(_04482_ ), .B(_04483_ ), .S(fanout_net_37 ), .Z(_04484_ ) );
OAI211_X1 _12238_ ( .A(fanout_net_39 ), .B(_04481_ ), .C1(_04484_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04485_ ) );
OAI211_X1 _12239_ ( .A(_04476_ ), .B(_04485_ ), .C1(_04456_ ), .C2(_04457_ ), .ZN(_04486_ ) );
NAND2_X1 _12240_ ( .A1(_04463_ ), .A2(_04486_ ), .ZN(_04487_ ) );
XNOR2_X2 _12241_ ( .A(_04487_ ), .B(_02294_ ), .ZN(_04488_ ) );
OR2_X1 _12242_ ( .A1(\myreg.Reg[0][21] ), .A2(fanout_net_33 ), .ZN(_04489_ ) );
OAI211_X1 _12243_ ( .A(_04489_ ), .B(_04465_ ), .C1(\myreg.Reg[1][21] ), .C2(_04469_ ), .ZN(_04490_ ) );
OR2_X1 _12244_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[2][21] ), .ZN(_04491_ ) );
OAI211_X1 _12245_ ( .A(_04491_ ), .B(fanout_net_37 ), .C1(_04469_ ), .C2(\myreg.Reg[3][21] ), .ZN(_04492_ ) );
NAND3_X1 _12246_ ( .A1(_04490_ ), .A2(_04492_ ), .A3(_04445_ ), .ZN(_04493_ ) );
MUX2_X1 _12247_ ( .A(\myreg.Reg[6][21] ), .B(\myreg.Reg[7][21] ), .S(fanout_net_33 ), .Z(_04494_ ) );
MUX2_X1 _12248_ ( .A(\myreg.Reg[4][21] ), .B(\myreg.Reg[5][21] ), .S(fanout_net_33 ), .Z(_04495_ ) );
MUX2_X1 _12249_ ( .A(_04494_ ), .B(_04495_ ), .S(_04436_ ), .Z(_04496_ ) );
OAI211_X1 _12250_ ( .A(_04434_ ), .B(_04493_ ), .C1(_04496_ ), .C2(_04475_ ), .ZN(_04497_ ) );
OR2_X1 _12251_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[14][21] ), .ZN(_04498_ ) );
OAI211_X1 _12252_ ( .A(_04498_ ), .B(fanout_net_37 ), .C1(_04469_ ), .C2(\myreg.Reg[15][21] ), .ZN(_04499_ ) );
OR2_X1 _12253_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[12][21] ), .ZN(_04500_ ) );
OAI211_X1 _12254_ ( .A(_04500_ ), .B(_04465_ ), .C1(_04469_ ), .C2(\myreg.Reg[13][21] ), .ZN(_04501_ ) );
NAND3_X1 _12255_ ( .A1(_04499_ ), .A2(_04501_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04502_ ) );
MUX2_X1 _12256_ ( .A(\myreg.Reg[8][21] ), .B(\myreg.Reg[9][21] ), .S(fanout_net_33 ), .Z(_04503_ ) );
MUX2_X1 _12257_ ( .A(\myreg.Reg[10][21] ), .B(\myreg.Reg[11][21] ), .S(fanout_net_33 ), .Z(_04504_ ) );
MUX2_X1 _12258_ ( .A(_04503_ ), .B(_04504_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04505_ ) );
OAI211_X1 _12259_ ( .A(fanout_net_39 ), .B(_04502_ ), .C1(_04505_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04506_ ) );
AOI21_X1 _12260_ ( .A(_03994_ ), .B1(_04497_ ), .B2(_04506_ ), .ZN(_04507_ ) );
INV_X1 _12261_ ( .A(\EX_LS_result_reg [21] ), .ZN(_04508_ ) );
NOR3_X1 _12262_ ( .A1(_04104_ ), .A2(_04508_ ), .A3(_04072_ ), .ZN(_04509_ ) );
NOR2_X1 _12263_ ( .A1(_04507_ ), .A2(_04509_ ), .ZN(_04510_ ) );
NAND2_X4 _12264_ ( .A1(_02297_ ), .A2(_02317_ ), .ZN(_04511_ ) );
AND2_X1 _12265_ ( .A1(_04510_ ), .A2(_04511_ ), .ZN(_04512_ ) );
NOR2_X1 _12266_ ( .A1(_04510_ ), .A2(_04511_ ), .ZN(_04513_ ) );
NOR3_X1 _12267_ ( .A1(_04488_ ), .A2(_04512_ ), .A3(_04513_ ), .ZN(_04514_ ) );
OR2_X1 _12268_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[0][23] ), .ZN(_04515_ ) );
OAI211_X1 _12269_ ( .A(_04515_ ), .B(_04005_ ), .C1(_04000_ ), .C2(\myreg.Reg[1][23] ), .ZN(_04516_ ) );
NOR2_X1 _12270_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[2][23] ), .ZN(_04517_ ) );
OAI21_X1 _12271_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(_04000_ ), .B2(\myreg.Reg[3][23] ), .ZN(_04518_ ) );
OAI211_X1 _12272_ ( .A(_04516_ ), .B(_03943_ ), .C1(_04517_ ), .C2(_04518_ ), .ZN(_04519_ ) );
MUX2_X1 _12273_ ( .A(\myreg.Reg[6][23] ), .B(\myreg.Reg[7][23] ), .S(fanout_net_33 ), .Z(_04520_ ) );
MUX2_X1 _12274_ ( .A(\myreg.Reg[4][23] ), .B(\myreg.Reg[5][23] ), .S(fanout_net_34 ), .Z(_04521_ ) );
MUX2_X1 _12275_ ( .A(_04520_ ), .B(_04521_ ), .S(_04005_ ), .Z(_04522_ ) );
OAI211_X1 _12276_ ( .A(_03930_ ), .B(_04519_ ), .C1(_04522_ ), .C2(_04014_ ), .ZN(_04523_ ) );
OR2_X1 _12277_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[8][23] ), .ZN(_04524_ ) );
OAI211_X1 _12278_ ( .A(_04524_ ), .B(_03996_ ), .C1(_04000_ ), .C2(\myreg.Reg[9][23] ), .ZN(_04525_ ) );
OR2_X1 _12279_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[10][23] ), .ZN(_04526_ ) );
OAI211_X1 _12280_ ( .A(_04526_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04000_ ), .C2(\myreg.Reg[11][23] ), .ZN(_04527_ ) );
NAND3_X1 _12281_ ( .A1(_04525_ ), .A2(_04527_ ), .A3(_03950_ ), .ZN(_04528_ ) );
MUX2_X1 _12282_ ( .A(\myreg.Reg[14][23] ), .B(\myreg.Reg[15][23] ), .S(fanout_net_34 ), .Z(_04529_ ) );
MUX2_X1 _12283_ ( .A(\myreg.Reg[12][23] ), .B(\myreg.Reg[13][23] ), .S(fanout_net_34 ), .Z(_04530_ ) );
MUX2_X1 _12284_ ( .A(_04529_ ), .B(_04530_ ), .S(_04005_ ), .Z(_04531_ ) );
OAI211_X1 _12285_ ( .A(fanout_net_39 ), .B(_04528_ ), .C1(_04531_ ), .C2(_04014_ ), .ZN(_04532_ ) );
NAND2_X1 _12286_ ( .A1(_04523_ ), .A2(_04532_ ), .ZN(_04533_ ) );
OAI21_X1 _12287_ ( .A(_04533_ ), .B1(_04104_ ), .B2(_04072_ ), .ZN(_04534_ ) );
NAND4_X1 _12288_ ( .A1(_02094_ ), .A2(\EX_LS_result_reg [23] ), .A3(_03988_ ), .A4(_03989_ ), .ZN(_04535_ ) );
AND2_X1 _12289_ ( .A1(_04534_ ), .A2(_04535_ ), .ZN(_04536_ ) );
XOR2_X1 _12290_ ( .A(_02247_ ), .B(_04536_ ), .Z(_04537_ ) );
INV_X1 _12291_ ( .A(_02270_ ), .ZN(_04538_ ) );
INV_X1 _12292_ ( .A(\EX_LS_result_reg [22] ), .ZN(_04539_ ) );
OR3_X1 _12293_ ( .A1(_04104_ ), .A2(_04539_ ), .A3(_04072_ ), .ZN(_04540_ ) );
OR2_X1 _12294_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[0][22] ), .ZN(_04541_ ) );
OAI211_X1 _12295_ ( .A(_04541_ ), .B(_04144_ ), .C1(_04145_ ), .C2(\myreg.Reg[1][22] ), .ZN(_04542_ ) );
OR2_X1 _12296_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[2][22] ), .ZN(_04543_ ) );
OAI211_X1 _12297_ ( .A(_04543_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04145_ ), .C2(\myreg.Reg[3][22] ), .ZN(_04544_ ) );
NAND3_X1 _12298_ ( .A1(_04542_ ), .A2(_04544_ ), .A3(_04014_ ), .ZN(_04545_ ) );
MUX2_X1 _12299_ ( .A(\myreg.Reg[6][22] ), .B(\myreg.Reg[7][22] ), .S(fanout_net_34 ), .Z(_04546_ ) );
MUX2_X1 _12300_ ( .A(\myreg.Reg[4][22] ), .B(\myreg.Reg[5][22] ), .S(fanout_net_34 ), .Z(_04547_ ) );
MUX2_X1 _12301_ ( .A(_04546_ ), .B(_04547_ ), .S(_04144_ ), .Z(_04548_ ) );
OAI211_X1 _12302_ ( .A(_04082_ ), .B(_04545_ ), .C1(_04548_ ), .C2(_04092_ ), .ZN(_04549_ ) );
OR2_X1 _12303_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[14][22] ), .ZN(_04550_ ) );
OAI211_X1 _12304_ ( .A(_04550_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04145_ ), .C2(\myreg.Reg[15][22] ), .ZN(_04551_ ) );
OR2_X1 _12305_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[12][22] ), .ZN(_04552_ ) );
OAI211_X1 _12306_ ( .A(_04552_ ), .B(_04144_ ), .C1(_04084_ ), .C2(\myreg.Reg[13][22] ), .ZN(_04553_ ) );
NAND3_X1 _12307_ ( .A1(_04551_ ), .A2(_04553_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04554_ ) );
MUX2_X1 _12308_ ( .A(\myreg.Reg[8][22] ), .B(\myreg.Reg[9][22] ), .S(fanout_net_34 ), .Z(_04555_ ) );
MUX2_X1 _12309_ ( .A(\myreg.Reg[10][22] ), .B(\myreg.Reg[11][22] ), .S(fanout_net_34 ), .Z(_04556_ ) );
MUX2_X1 _12310_ ( .A(_04555_ ), .B(_04556_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04557_ ) );
OAI211_X1 _12311_ ( .A(fanout_net_39 ), .B(_04554_ ), .C1(_04557_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04558_ ) );
NAND2_X1 _12312_ ( .A1(_04549_ ), .A2(_04558_ ), .ZN(_04559_ ) );
OAI21_X1 _12313_ ( .A(_04559_ ), .B1(_04104_ ), .B2(_04072_ ), .ZN(_04560_ ) );
AND2_X1 _12314_ ( .A1(_04540_ ), .A2(_04560_ ), .ZN(_04561_ ) );
XNOR2_X1 _12315_ ( .A(_04538_ ), .B(_04561_ ), .ZN(_04562_ ) );
NAND3_X1 _12316_ ( .A1(_04514_ ), .A2(_04537_ ), .A3(_04562_ ), .ZN(_04563_ ) );
NOR2_X1 _12317_ ( .A1(_04462_ ), .A2(_04563_ ), .ZN(_04564_ ) );
OR2_X1 _12318_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04565_ ) );
OAI211_X1 _12319_ ( .A(_04565_ ), .B(_04436_ ), .C1(_04437_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04566_ ) );
OR2_X1 _12320_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04567_ ) );
OAI211_X1 _12321_ ( .A(_04567_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04437_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04568_ ) );
NAND3_X1 _12322_ ( .A1(_04566_ ), .A2(_04568_ ), .A3(_04369_ ), .ZN(_04569_ ) );
MUX2_X1 _12323_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04570_ ) );
MUX2_X1 _12324_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04571_ ) );
MUX2_X1 _12325_ ( .A(_04570_ ), .B(_04571_ ), .S(_04360_ ), .Z(_04572_ ) );
OAI211_X1 _12326_ ( .A(_04434_ ), .B(_04569_ ), .C1(_04572_ ), .C2(_04445_ ), .ZN(_04573_ ) );
OR2_X1 _12327_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04574_ ) );
OAI211_X1 _12328_ ( .A(_04574_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04437_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04575_ ) );
OR2_X1 _12329_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04576_ ) );
OAI211_X1 _12330_ ( .A(_04576_ ), .B(_04360_ ), .C1(_04437_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04577_ ) );
NAND3_X1 _12331_ ( .A1(_04575_ ), .A2(_04577_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04578_ ) );
MUX2_X1 _12332_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04579_ ) );
MUX2_X1 _12333_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04580_ ) );
MUX2_X1 _12334_ ( .A(_04579_ ), .B(_04580_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04581_ ) );
OAI211_X1 _12335_ ( .A(fanout_net_39 ), .B(_04578_ ), .C1(_04581_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04582_ ) );
AOI21_X1 _12336_ ( .A(_03994_ ), .B1(_04573_ ), .B2(_04582_ ), .ZN(_04583_ ) );
AND2_X1 _12337_ ( .A1(_03994_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04584_ ) );
NOR2_X1 _12338_ ( .A1(_04583_ ), .A2(_04584_ ), .ZN(_04585_ ) );
NOR2_X1 _12339_ ( .A1(_04585_ ), .A2(_02940_ ), .ZN(_04586_ ) );
NOR3_X1 _12340_ ( .A1(_02934_ ), .A2(_04583_ ), .A3(_04584_ ), .ZN(_04587_ ) );
NOR2_X1 _12341_ ( .A1(_04586_ ), .A2(_04587_ ), .ZN(_04588_ ) );
OR3_X1 _12342_ ( .A1(_04139_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_04141_ ), .ZN(_04589_ ) );
OR2_X1 _12343_ ( .A1(fanout_net_34 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04590_ ) );
OAI211_X1 _12344_ ( .A(_04590_ ), .B(_04436_ ), .C1(_04469_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04591_ ) );
OR2_X1 _12345_ ( .A1(fanout_net_34 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04592_ ) );
OAI211_X1 _12346_ ( .A(_04592_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04469_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04593_ ) );
NAND3_X1 _12347_ ( .A1(_04591_ ), .A2(_04593_ ), .A3(_04369_ ), .ZN(_04594_ ) );
MUX2_X1 _12348_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04595_ ) );
MUX2_X1 _12349_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04596_ ) );
MUX2_X1 _12350_ ( .A(_04595_ ), .B(_04596_ ), .S(_04436_ ), .Z(_04597_ ) );
OAI211_X1 _12351_ ( .A(fanout_net_39 ), .B(_04594_ ), .C1(_04597_ ), .C2(_04445_ ), .ZN(_04598_ ) );
OR2_X1 _12352_ ( .A1(fanout_net_34 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04599_ ) );
OAI211_X1 _12353_ ( .A(_04599_ ), .B(_04436_ ), .C1(_04469_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04600_ ) );
OR2_X1 _12354_ ( .A1(fanout_net_34 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04601_ ) );
OAI211_X1 _12355_ ( .A(_04601_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04437_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04602_ ) );
NAND3_X1 _12356_ ( .A1(_04600_ ), .A2(_04602_ ), .A3(_04369_ ), .ZN(_04603_ ) );
MUX2_X1 _12357_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04604_ ) );
MUX2_X1 _12358_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04605_ ) );
MUX2_X1 _12359_ ( .A(_04604_ ), .B(_04605_ ), .S(_04436_ ), .Z(_04606_ ) );
OAI211_X1 _12360_ ( .A(_04434_ ), .B(_04603_ ), .C1(_04606_ ), .C2(_04445_ ), .ZN(_04607_ ) );
OAI211_X1 _12361_ ( .A(_04598_ ), .B(_04607_ ), .C1(_04456_ ), .C2(_04457_ ), .ZN(_04608_ ) );
NAND2_X1 _12362_ ( .A1(_04589_ ), .A2(_04608_ ), .ZN(_04609_ ) );
XNOR2_X1 _12363_ ( .A(_04609_ ), .B(_02167_ ), .ZN(_04610_ ) );
AND2_X1 _12364_ ( .A1(_04588_ ), .A2(_04610_ ), .ZN(_04611_ ) );
OR3_X1 _12365_ ( .A1(_04456_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_04457_ ), .ZN(_04612_ ) );
OR2_X1 _12366_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04613_ ) );
BUF_X4 _12367_ ( .A(_04436_ ), .Z(_04614_ ) );
OAI211_X1 _12368_ ( .A(_04613_ ), .B(_04614_ ), .C1(_04466_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04615_ ) );
OR2_X1 _12369_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04616_ ) );
OAI211_X1 _12370_ ( .A(_04616_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04466_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04617_ ) );
NAND3_X1 _12371_ ( .A1(_04615_ ), .A2(_04617_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04618_ ) );
MUX2_X1 _12372_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04619_ ) );
MUX2_X1 _12373_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04620_ ) );
MUX2_X1 _12374_ ( .A(_04619_ ), .B(_04620_ ), .S(_04465_ ), .Z(_04621_ ) );
OAI211_X1 _12375_ ( .A(_04434_ ), .B(_04618_ ), .C1(_04621_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04622_ ) );
NOR2_X1 _12376_ ( .A1(_04466_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04623_ ) );
OAI21_X1 _12377_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_35 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04624_ ) );
NOR2_X1 _12378_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04625_ ) );
OAI21_X1 _12379_ ( .A(_04465_ ), .B1(_04466_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04626_ ) );
OAI221_X1 _12380_ ( .A(_04445_ ), .B1(_04623_ ), .B2(_04624_ ), .C1(_04625_ ), .C2(_04626_ ), .ZN(_04627_ ) );
MUX2_X1 _12381_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04628_ ) );
MUX2_X1 _12382_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04629_ ) );
MUX2_X1 _12383_ ( .A(_04628_ ), .B(_04629_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04630_ ) );
OAI211_X1 _12384_ ( .A(fanout_net_39 ), .B(_04627_ ), .C1(_04630_ ), .C2(_04475_ ), .ZN(_04631_ ) );
OAI211_X1 _12385_ ( .A(_04622_ ), .B(_04631_ ), .C1(_04456_ ), .C2(_04457_ ), .ZN(_04632_ ) );
NAND2_X1 _12386_ ( .A1(_04612_ ), .A2(_04632_ ), .ZN(_04633_ ) );
XNOR2_X1 _12387_ ( .A(_04633_ ), .B(_02990_ ), .ZN(_04634_ ) );
NAND2_X1 _12388_ ( .A1(_03994_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .ZN(_04635_ ) );
OR2_X1 _12389_ ( .A1(fanout_net_35 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04636_ ) );
OAI211_X1 _12390_ ( .A(_04636_ ), .B(_04360_ ), .C1(_04361_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04637_ ) );
OR2_X1 _12391_ ( .A1(fanout_net_35 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04638_ ) );
OAI211_X1 _12392_ ( .A(_04638_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04361_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04639_ ) );
NAND3_X1 _12393_ ( .A1(_04637_ ), .A2(_04639_ ), .A3(_04369_ ), .ZN(_04640_ ) );
MUX2_X1 _12394_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04641_ ) );
MUX2_X1 _12395_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04642_ ) );
MUX2_X1 _12396_ ( .A(_04641_ ), .B(_04642_ ), .S(_04360_ ), .Z(_04643_ ) );
OAI211_X1 _12397_ ( .A(_04082_ ), .B(_04640_ ), .C1(_04643_ ), .C2(_04369_ ), .ZN(_04644_ ) );
OR2_X1 _12398_ ( .A1(fanout_net_35 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04645_ ) );
OAI211_X1 _12399_ ( .A(_04645_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04361_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04646_ ) );
OR2_X1 _12400_ ( .A1(fanout_net_35 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04647_ ) );
OAI211_X1 _12401_ ( .A(_04647_ ), .B(_04360_ ), .C1(_04361_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04648_ ) );
NAND3_X1 _12402_ ( .A1(_04646_ ), .A2(_04648_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04649_ ) );
MUX2_X1 _12403_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04650_ ) );
MUX2_X1 _12404_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04651_ ) );
MUX2_X1 _12405_ ( .A(_04650_ ), .B(_04651_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04652_ ) );
OAI211_X1 _12406_ ( .A(fanout_net_39 ), .B(_04649_ ), .C1(_04652_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04653_ ) );
NAND2_X1 _12407_ ( .A1(_04644_ ), .A2(_04653_ ), .ZN(_04654_ ) );
OAI21_X1 _12408_ ( .A(_04654_ ), .B1(_04104_ ), .B2(_04072_ ), .ZN(_04655_ ) );
AND2_X1 _12409_ ( .A1(_04635_ ), .A2(_04655_ ), .ZN(_04656_ ) );
INV_X1 _12410_ ( .A(_04656_ ), .ZN(_04657_ ) );
XNOR2_X2 _12411_ ( .A(_02963_ ), .B(_04657_ ), .ZN(_04658_ ) );
AND3_X1 _12412_ ( .A1(_04611_ ), .A2(_04634_ ), .A3(_04658_ ), .ZN(_04659_ ) );
NOR2_X1 _12413_ ( .A1(_04139_ ), .A2(_04457_ ), .ZN(_04660_ ) );
INV_X1 _12414_ ( .A(_04660_ ), .ZN(_04661_ ) );
OR2_X1 _12415_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04662_ ) );
BUF_X4 _12416_ ( .A(_04437_ ), .Z(_04663_ ) );
OAI211_X1 _12417_ ( .A(_04662_ ), .B(_04614_ ), .C1(_04663_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04664_ ) );
OR2_X1 _12418_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04665_ ) );
OAI211_X1 _12419_ ( .A(_04665_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04663_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04666_ ) );
NAND3_X1 _12420_ ( .A1(_04664_ ), .A2(_04666_ ), .A3(_04475_ ), .ZN(_04667_ ) );
MUX2_X1 _12421_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04668_ ) );
MUX2_X1 _12422_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04669_ ) );
MUX2_X1 _12423_ ( .A(_04668_ ), .B(_04669_ ), .S(_04614_ ), .Z(_04670_ ) );
OAI211_X1 _12424_ ( .A(fanout_net_39 ), .B(_04667_ ), .C1(_04670_ ), .C2(_04475_ ), .ZN(_04671_ ) );
OR2_X1 _12425_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04672_ ) );
OAI211_X1 _12426_ ( .A(_04672_ ), .B(_04465_ ), .C1(_04466_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04673_ ) );
NOR2_X1 _12427_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04674_ ) );
OAI21_X1 _12428_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(_04466_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04675_ ) );
OAI211_X1 _12429_ ( .A(_04673_ ), .B(_04445_ ), .C1(_04674_ ), .C2(_04675_ ), .ZN(_04676_ ) );
MUX2_X1 _12430_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04677_ ) );
MUX2_X1 _12431_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04678_ ) );
MUX2_X1 _12432_ ( .A(_04677_ ), .B(_04678_ ), .S(_04465_ ), .Z(_04679_ ) );
OAI211_X1 _12433_ ( .A(_04434_ ), .B(_04676_ ), .C1(_04679_ ), .C2(_04475_ ), .ZN(_04680_ ) );
NAND3_X1 _12434_ ( .A1(_04661_ ), .A2(_04671_ ), .A3(_04680_ ), .ZN(_04681_ ) );
INV_X1 _12435_ ( .A(\EX_LS_result_reg [26] ), .ZN(_04682_ ) );
OR3_X1 _12436_ ( .A1(_04456_ ), .A2(_04682_ ), .A3(_04457_ ), .ZN(_04683_ ) );
NAND2_X1 _12437_ ( .A1(_04681_ ), .A2(_04683_ ), .ZN(_04684_ ) );
XNOR2_X1 _12438_ ( .A(_04684_ ), .B(_02196_ ), .ZN(_04685_ ) );
OR2_X1 _12439_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04686_ ) );
OAI211_X1 _12440_ ( .A(_04686_ ), .B(_04614_ ), .C1(_04663_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04687_ ) );
OR2_X1 _12441_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04688_ ) );
OAI211_X1 _12442_ ( .A(_04688_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04663_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04689_ ) );
NAND3_X1 _12443_ ( .A1(_04687_ ), .A2(_04689_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04690_ ) );
MUX2_X1 _12444_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04691_ ) );
MUX2_X1 _12445_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04692_ ) );
MUX2_X1 _12446_ ( .A(_04691_ ), .B(_04692_ ), .S(_04614_ ), .Z(_04693_ ) );
OAI211_X1 _12447_ ( .A(_04434_ ), .B(_04690_ ), .C1(_04693_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04694_ ) );
NOR2_X1 _12448_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04695_ ) );
OAI21_X1 _12449_ ( .A(_04465_ ), .B1(_04466_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04696_ ) );
MUX2_X1 _12450_ ( .A(_02212_ ), .B(_02213_ ), .S(fanout_net_35 ), .Z(_04697_ ) );
OAI221_X1 _12451_ ( .A(_04445_ ), .B1(_04695_ ), .B2(_04696_ ), .C1(_04697_ ), .C2(_04614_ ), .ZN(_04698_ ) );
MUX2_X1 _12452_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04699_ ) );
MUX2_X1 _12453_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04700_ ) );
MUX2_X1 _12454_ ( .A(_04699_ ), .B(_04700_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04701_ ) );
OAI211_X1 _12455_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04698_ ), .C1(_04701_ ), .C2(_04475_ ), .ZN(_04702_ ) );
NAND3_X1 _12456_ ( .A1(_04661_ ), .A2(_04694_ ), .A3(_04702_ ), .ZN(_04703_ ) );
INV_X1 _12457_ ( .A(\EX_LS_result_reg [27] ), .ZN(_04704_ ) );
OR3_X1 _12458_ ( .A1(_04456_ ), .A2(_04704_ ), .A3(_04457_ ), .ZN(_04705_ ) );
NAND2_X1 _12459_ ( .A1(_04703_ ), .A2(_04705_ ), .ZN(_04706_ ) );
NAND2_X1 _12460_ ( .A1(_02199_ ), .A2(_02220_ ), .ZN(_04707_ ) );
INV_X1 _12461_ ( .A(_04707_ ), .ZN(_04708_ ) );
OR2_X1 _12462_ ( .A1(_04706_ ), .A2(_04708_ ), .ZN(_04709_ ) );
NAND2_X1 _12463_ ( .A1(_04706_ ), .A2(_04708_ ), .ZN(_04710_ ) );
AND3_X1 _12464_ ( .A1(_04685_ ), .A2(_04709_ ), .A3(_04710_ ), .ZN(_04711_ ) );
OR2_X1 _12465_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04712_ ) );
OAI211_X1 _12466_ ( .A(_04712_ ), .B(_04614_ ), .C1(_04663_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04713_ ) );
OR2_X1 _12467_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04714_ ) );
OAI211_X1 _12468_ ( .A(_04714_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04663_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04715_ ) );
NAND3_X1 _12469_ ( .A1(_04713_ ), .A2(_04715_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04716_ ) );
MUX2_X1 _12470_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04717_ ) );
MUX2_X1 _12471_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04718_ ) );
MUX2_X1 _12472_ ( .A(_04717_ ), .B(_04718_ ), .S(_04614_ ), .Z(_04719_ ) );
OAI211_X1 _12473_ ( .A(_04434_ ), .B(_04716_ ), .C1(_04719_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04720_ ) );
NOR2_X1 _12474_ ( .A1(_04663_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04721_ ) );
OAI21_X1 _12475_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04722_ ) );
NOR2_X1 _12476_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04723_ ) );
OAI21_X1 _12477_ ( .A(_04614_ ), .B1(_04663_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04724_ ) );
OAI221_X1 _12478_ ( .A(_04475_ ), .B1(_04721_ ), .B2(_04722_ ), .C1(_04723_ ), .C2(_04724_ ), .ZN(_04725_ ) );
MUX2_X1 _12479_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04726_ ) );
MUX2_X1 _12480_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04727_ ) );
MUX2_X1 _12481_ ( .A(_04726_ ), .B(_04727_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04728_ ) );
OAI211_X1 _12482_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04725_ ), .C1(_04728_ ), .C2(_04475_ ), .ZN(_04729_ ) );
NAND3_X1 _12483_ ( .A1(_04661_ ), .A2(_04720_ ), .A3(_04729_ ), .ZN(_04730_ ) );
INV_X1 _12484_ ( .A(\EX_LS_result_reg [24] ), .ZN(_04731_ ) );
OR3_X1 _12485_ ( .A1(_04456_ ), .A2(_04731_ ), .A3(_04457_ ), .ZN(_04732_ ) );
NAND2_X1 _12486_ ( .A1(_04730_ ), .A2(_04732_ ), .ZN(_04733_ ) );
XNOR2_X1 _12487_ ( .A(_04733_ ), .B(_02876_ ), .ZN(_04734_ ) );
OR2_X1 _12488_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04735_ ) );
OAI211_X1 _12489_ ( .A(_04735_ ), .B(_04614_ ), .C1(_04663_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04736_ ) );
OR2_X1 _12490_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04737_ ) );
OAI211_X1 _12491_ ( .A(_04737_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04663_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04738_ ) );
NAND3_X1 _12492_ ( .A1(_04736_ ), .A2(_04738_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04739_ ) );
MUX2_X1 _12493_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04740_ ) );
MUX2_X1 _12494_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04741_ ) );
MUX2_X1 _12495_ ( .A(_04740_ ), .B(_04741_ ), .S(_04465_ ), .Z(_04742_ ) );
OAI211_X1 _12496_ ( .A(_04434_ ), .B(_04739_ ), .C1(_04742_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04743_ ) );
NOR2_X1 _12497_ ( .A1(_04466_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04744_ ) );
OAI21_X1 _12498_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04745_ ) );
NOR2_X1 _12499_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04746_ ) );
OAI21_X1 _12500_ ( .A(_04465_ ), .B1(_04466_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04747_ ) );
OAI221_X1 _12501_ ( .A(_04445_ ), .B1(_04744_ ), .B2(_04745_ ), .C1(_04746_ ), .C2(_04747_ ), .ZN(_04748_ ) );
MUX2_X1 _12502_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04749_ ) );
MUX2_X1 _12503_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04750_ ) );
MUX2_X1 _12504_ ( .A(_04749_ ), .B(_04750_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04751_ ) );
OAI211_X1 _12505_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04748_ ), .C1(_04751_ ), .C2(_04475_ ), .ZN(_04752_ ) );
NAND3_X1 _12506_ ( .A1(_04661_ ), .A2(_04743_ ), .A3(_04752_ ), .ZN(_04753_ ) );
INV_X1 _12507_ ( .A(\EX_LS_result_reg [25] ), .ZN(_04754_ ) );
OR3_X1 _12508_ ( .A1(_04456_ ), .A2(_04754_ ), .A3(_04457_ ), .ZN(_04755_ ) );
NAND2_X1 _12509_ ( .A1(_04753_ ), .A2(_04755_ ), .ZN(_04756_ ) );
NAND2_X1 _12510_ ( .A1(_04756_ ), .A2(_02907_ ), .ZN(_04757_ ) );
NAND3_X1 _12511_ ( .A1(_04753_ ), .A2(_02899_ ), .A3(_04755_ ), .ZN(_04758_ ) );
AND2_X2 _12512_ ( .A1(_04757_ ), .A2(_04758_ ), .ZN(_04759_ ) );
AND2_X1 _12513_ ( .A1(_04734_ ), .A2(_04759_ ), .ZN(_04760_ ) );
AND3_X2 _12514_ ( .A1(_04659_ ), .A2(_04711_ ), .A3(_04760_ ), .ZN(_04761_ ) );
AND2_X1 _12515_ ( .A1(_04564_ ), .A2(_04761_ ), .ZN(_04762_ ) );
AND2_X1 _12516_ ( .A1(_04356_ ), .A2(_04762_ ), .ZN(_04763_ ) );
NOR2_X1 _12517_ ( .A1(_03877_ ), .A2(\ID_EX_typ [1] ), .ZN(_04764_ ) );
AND2_X1 _12518_ ( .A1(_04764_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04765_ ) );
INV_X1 _12519_ ( .A(_04765_ ), .ZN(_04766_ ) );
INV_X1 _12520_ ( .A(\ID_EX_typ [1] ), .ZN(_04767_ ) );
NOR2_X1 _12521_ ( .A1(_04767_ ), .A2(fanout_net_5 ), .ZN(_04768_ ) );
INV_X2 _12522_ ( .A(\ID_EX_typ [2] ), .ZN(_04769_ ) );
AND2_X2 _12523_ ( .A1(_04768_ ), .A2(_04769_ ), .ZN(_04770_ ) );
INV_X1 _12524_ ( .A(_04770_ ), .ZN(_04771_ ) );
INV_X1 _12525_ ( .A(fanout_net_6 ), .ZN(_04772_ ) );
BUF_X4 _12526_ ( .A(_04772_ ), .Z(_04773_ ) );
BUF_X4 _12527_ ( .A(_04773_ ), .Z(_04774_ ) );
NAND3_X1 _12528_ ( .A1(_04589_ ), .A2(_04774_ ), .A3(_04608_ ), .ZN(_04775_ ) );
NAND2_X1 _12529_ ( .A1(fanout_net_6 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04776_ ) );
AND2_X2 _12530_ ( .A1(_04775_ ), .A2(_04776_ ), .ZN(_04777_ ) );
INV_X1 _12531_ ( .A(_02167_ ), .ZN(_04778_ ) );
XNOR2_X1 _12532_ ( .A(_04777_ ), .B(_04778_ ), .ZN(_04779_ ) );
INV_X1 _12533_ ( .A(_04779_ ), .ZN(_04780_ ) );
OAI21_X1 _12534_ ( .A(_04774_ ), .B1(_04583_ ), .B2(_04584_ ), .ZN(_04781_ ) );
NAND2_X1 _12535_ ( .A1(fanout_net_6 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04782_ ) );
AND2_X2 _12536_ ( .A1(_04781_ ), .A2(_04782_ ), .ZN(_04783_ ) );
AND2_X1 _12537_ ( .A1(_04783_ ), .A2(_02934_ ), .ZN(_04784_ ) );
AOI21_X1 _12538_ ( .A(_02934_ ), .B1(_04781_ ), .B2(_04782_ ), .ZN(_04785_ ) );
OAI21_X1 _12539_ ( .A(_04780_ ), .B1(_04784_ ), .B2(_04785_ ), .ZN(_04786_ ) );
BUF_X2 _12540_ ( .A(_04774_ ), .Z(_04787_ ) );
NAND3_X1 _12541_ ( .A1(_04681_ ), .A2(_04787_ ), .A3(_04683_ ), .ZN(_04788_ ) );
NAND2_X1 _12542_ ( .A1(_02197_ ), .A2(fanout_net_6 ), .ZN(_04789_ ) );
NAND2_X1 _12543_ ( .A1(_04788_ ), .A2(_04789_ ), .ZN(_04790_ ) );
INV_X1 _12544_ ( .A(_02196_ ), .ZN(_04791_ ) );
NOR2_X1 _12545_ ( .A1(_04790_ ), .A2(_04791_ ), .ZN(_04792_ ) );
AOI21_X1 _12546_ ( .A(_02196_ ), .B1(_04788_ ), .B2(_04789_ ), .ZN(_04793_ ) );
NOR2_X1 _12547_ ( .A1(_04792_ ), .A2(_04793_ ), .ZN(_04794_ ) );
INV_X1 _12548_ ( .A(_04794_ ), .ZN(_04795_ ) );
NAND3_X1 _12549_ ( .A1(_04703_ ), .A2(_04774_ ), .A3(_04705_ ), .ZN(_04796_ ) );
NAND2_X1 _12550_ ( .A1(_02200_ ), .A2(fanout_net_6 ), .ZN(_04797_ ) );
NAND2_X1 _12551_ ( .A1(_04796_ ), .A2(_04797_ ), .ZN(_04798_ ) );
NOR2_X1 _12552_ ( .A1(_04798_ ), .A2(_04708_ ), .ZN(_04799_ ) );
AOI21_X1 _12553_ ( .A(_04707_ ), .B1(_04796_ ), .B2(_04797_ ), .ZN(_04800_ ) );
NOR2_X1 _12554_ ( .A1(_04799_ ), .A2(_04800_ ), .ZN(_04801_ ) );
INV_X1 _12555_ ( .A(_04801_ ), .ZN(_04802_ ) );
NAND2_X1 _12556_ ( .A1(_04795_ ), .A2(_04802_ ), .ZN(_04803_ ) );
NAND3_X1 _12557_ ( .A1(_04730_ ), .A2(_04787_ ), .A3(_04732_ ), .ZN(_04804_ ) );
NAND2_X1 _12558_ ( .A1(_02877_ ), .A2(fanout_net_6 ), .ZN(_04805_ ) );
NAND2_X1 _12559_ ( .A1(_04804_ ), .A2(_04805_ ), .ZN(_04806_ ) );
INV_X1 _12560_ ( .A(_02876_ ), .ZN(_04807_ ) );
NOR2_X1 _12561_ ( .A1(_04806_ ), .A2(_04807_ ), .ZN(_04808_ ) );
AOI21_X1 _12562_ ( .A(_02876_ ), .B1(_04804_ ), .B2(_04805_ ), .ZN(_04809_ ) );
NOR2_X1 _12563_ ( .A1(_04808_ ), .A2(_04809_ ), .ZN(_04810_ ) );
NAND3_X1 _12564_ ( .A1(_04753_ ), .A2(_04787_ ), .A3(_04755_ ), .ZN(_04811_ ) );
NAND2_X1 _12565_ ( .A1(_02900_ ), .A2(fanout_net_6 ), .ZN(_04812_ ) );
NAND2_X1 _12566_ ( .A1(_04811_ ), .A2(_04812_ ), .ZN(_04813_ ) );
NOR2_X1 _12567_ ( .A1(_04813_ ), .A2(_02907_ ), .ZN(_04814_ ) );
AOI21_X1 _12568_ ( .A(_02899_ ), .B1(_04811_ ), .B2(_04812_ ), .ZN(_04815_ ) );
NOR2_X1 _12569_ ( .A1(_04814_ ), .A2(_04815_ ), .ZN(_04816_ ) );
NOR3_X1 _12570_ ( .A1(_04803_ ), .A2(_04810_ ), .A3(_04816_ ), .ZN(_04817_ ) );
AOI21_X1 _12571_ ( .A(fanout_net_6 ), .B1(_04111_ ), .B2(_04131_ ), .ZN(_04818_ ) );
AND2_X1 _12572_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [15] ), .ZN(_04819_ ) );
NOR2_X4 _12573_ ( .A1(_04818_ ), .A2(_04819_ ), .ZN(_04820_ ) );
XNOR2_X1 _12574_ ( .A(_04820_ ), .B(_02694_ ), .ZN(_04821_ ) );
NAND3_X1 _12575_ ( .A1(_04142_ ), .A2(_04773_ ), .A3(_04163_ ), .ZN(_04822_ ) );
NAND2_X1 _12576_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [14] ), .ZN(_04823_ ) );
AND2_X1 _12577_ ( .A1(_04822_ ), .A2(_04823_ ), .ZN(_04824_ ) );
NOR2_X1 _12578_ ( .A1(_04824_ ), .A2(_04134_ ), .ZN(_04825_ ) );
INV_X1 _12579_ ( .A(_04825_ ), .ZN(_04826_ ) );
NAND3_X1 _12580_ ( .A1(_04822_ ), .A2(_04134_ ), .A3(_04823_ ), .ZN(_04827_ ) );
AOI21_X1 _12581_ ( .A(_04821_ ), .B1(_04826_ ), .B2(_04827_ ), .ZN(_04828_ ) );
NAND3_X1 _12582_ ( .A1(_04052_ ), .A2(_04773_ ), .A3(_04073_ ), .ZN(_04829_ ) );
NAND2_X1 _12583_ ( .A1(_02669_ ), .A2(fanout_net_6 ), .ZN(_04830_ ) );
NAND2_X1 _12584_ ( .A1(_04829_ ), .A2(_04830_ ), .ZN(_04831_ ) );
XNOR2_X1 _12585_ ( .A(_04831_ ), .B(_04075_ ), .ZN(_04832_ ) );
INV_X1 _12586_ ( .A(_04832_ ), .ZN(_04833_ ) );
NAND3_X1 _12587_ ( .A1(_04081_ ), .A2(_04773_ ), .A3(_04105_ ), .ZN(_04834_ ) );
NAND2_X1 _12588_ ( .A1(_02648_ ), .A2(fanout_net_6 ), .ZN(_04835_ ) );
NAND2_X1 _12589_ ( .A1(_04834_ ), .A2(_04835_ ), .ZN(_04836_ ) );
XNOR2_X1 _12590_ ( .A(_04836_ ), .B(_02647_ ), .ZN(_04837_ ) );
INV_X1 _12591_ ( .A(_04837_ ), .ZN(_04838_ ) );
AND3_X1 _12592_ ( .A1(_04828_ ), .A2(_04833_ ), .A3(_04838_ ), .ZN(_04839_ ) );
OR2_X1 _12593_ ( .A1(_04047_ ), .A2(fanout_net_6 ), .ZN(_04840_ ) );
NAND2_X1 _12594_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [9] ), .ZN(_04841_ ) );
AND2_X1 _12595_ ( .A1(_04840_ ), .A2(_04841_ ), .ZN(_04842_ ) );
XNOR2_X1 _12596_ ( .A(_04842_ ), .B(_02812_ ), .ZN(_04843_ ) );
INV_X1 _12597_ ( .A(_04843_ ), .ZN(_04844_ ) );
OR3_X1 _12598_ ( .A1(_04019_ ), .A2(fanout_net_6 ), .A3(_04020_ ), .ZN(_04845_ ) );
NAND2_X1 _12599_ ( .A1(_02790_ ), .A2(fanout_net_6 ), .ZN(_04846_ ) );
NAND2_X1 _12600_ ( .A1(_04845_ ), .A2(_04846_ ), .ZN(_04847_ ) );
XNOR2_X1 _12601_ ( .A(_04847_ ), .B(_02789_ ), .ZN(_04848_ ) );
INV_X1 _12602_ ( .A(_04848_ ), .ZN(_04849_ ) );
NAND3_X1 _12603_ ( .A1(_03928_ ), .A2(_04773_ ), .A3(_03963_ ), .ZN(_04850_ ) );
NAND2_X1 _12604_ ( .A1(_02766_ ), .A2(fanout_net_6 ), .ZN(_04851_ ) );
NAND2_X1 _12605_ ( .A1(_04850_ ), .A2(_04851_ ), .ZN(_04852_ ) );
XNOR2_X1 _12606_ ( .A(_04852_ ), .B(_02765_ ), .ZN(_04853_ ) );
AOI21_X1 _12607_ ( .A(fanout_net_6 ), .B1(_03986_ ), .B2(_03990_ ), .ZN(_04854_ ) );
AND2_X1 _12608_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [10] ), .ZN(_04855_ ) );
NOR2_X1 _12609_ ( .A1(_04854_ ), .A2(_04855_ ), .ZN(_04856_ ) );
XNOR2_X1 _12610_ ( .A(_04856_ ), .B(_02742_ ), .ZN(_04857_ ) );
NOR2_X1 _12611_ ( .A1(_04853_ ), .A2(_04857_ ), .ZN(_04858_ ) );
NAND4_X1 _12612_ ( .A1(_04839_ ), .A2(_04844_ ), .A3(_04849_ ), .A4(_04858_ ), .ZN(_04859_ ) );
NAND2_X2 _12613_ ( .A1(_04256_ ), .A2(_04772_ ), .ZN(_04860_ ) );
BUF_X4 _12614_ ( .A(_04860_ ), .Z(_04861_ ) );
NAND2_X1 _12615_ ( .A1(_02465_ ), .A2(fanout_net_6 ), .ZN(_04862_ ) );
BUF_X4 _12616_ ( .A(_04862_ ), .Z(_04863_ ) );
AND3_X4 _12617_ ( .A1(_04861_ ), .A2(_02464_ ), .A3(_04863_ ), .ZN(_04864_ ) );
AOI21_X1 _12618_ ( .A(_02464_ ), .B1(_04861_ ), .B2(_04863_ ), .ZN(_04865_ ) );
NOR2_X2 _12619_ ( .A1(_04864_ ), .A2(_04865_ ), .ZN(_04866_ ) );
NAND3_X1 _12620_ ( .A1(_04351_ ), .A2(_04772_ ), .A3(_04352_ ), .ZN(_04867_ ) );
OR2_X1 _12621_ ( .A1(_04772_ ), .A2(\ID_EX_imm [0] ), .ZN(_04868_ ) );
NAND2_X2 _12622_ ( .A1(_04867_ ), .A2(_04868_ ), .ZN(_04869_ ) );
NOR2_X1 _12623_ ( .A1(_04331_ ), .A2(_04869_ ), .ZN(_04870_ ) );
NOR2_X1 _12624_ ( .A1(_04866_ ), .A2(_04870_ ), .ZN(_04871_ ) );
NAND2_X4 _12625_ ( .A1(_04860_ ), .A2(_04862_ ), .ZN(_04872_ ) );
AOI21_X1 _12626_ ( .A(_04871_ ), .B1(_02464_ ), .B2(_04872_ ), .ZN(_04873_ ) );
NAND3_X1 _12627_ ( .A1(_04308_ ), .A2(_04773_ ), .A3(_04327_ ), .ZN(_04874_ ) );
NAND2_X1 _12628_ ( .A1(fanout_net_6 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_04875_ ) );
AND2_X2 _12629_ ( .A1(_04874_ ), .A2(_04875_ ), .ZN(_04876_ ) );
XNOR2_X1 _12630_ ( .A(_04876_ ), .B(_02520_ ), .ZN(_04877_ ) );
NAND3_X1 _12631_ ( .A1(_04303_ ), .A2(_04773_ ), .A3(_04301_ ), .ZN(_04878_ ) );
NAND2_X1 _12632_ ( .A1(_02442_ ), .A2(fanout_net_6 ), .ZN(_04879_ ) );
NAND2_X2 _12633_ ( .A1(_04878_ ), .A2(_04879_ ), .ZN(_04880_ ) );
XNOR2_X1 _12634_ ( .A(_04880_ ), .B(_02441_ ), .ZN(_04881_ ) );
OR3_X2 _12635_ ( .A1(_04873_ ), .A2(_04877_ ), .A3(_04881_ ), .ZN(_04882_ ) );
OR2_X1 _12636_ ( .A1(_04876_ ), .A2(_02520_ ), .ZN(_04883_ ) );
AND2_X1 _12637_ ( .A1(_04876_ ), .A2(_02516_ ), .ZN(_04884_ ) );
NOR2_X1 _12638_ ( .A1(_04876_ ), .A2(_02516_ ), .ZN(_04885_ ) );
OAI211_X1 _12639_ ( .A(_02441_ ), .B(_04880_ ), .C1(_04884_ ), .C2(_04885_ ), .ZN(_04886_ ) );
NAND3_X1 _12640_ ( .A1(_04882_ ), .A2(_04883_ ), .A3(_04886_ ), .ZN(_04887_ ) );
NAND3_X1 _12641_ ( .A1(_04210_ ), .A2(_04773_ ), .A3(_04211_ ), .ZN(_04888_ ) );
OR2_X1 _12642_ ( .A1(_04772_ ), .A2(\ID_EX_imm [7] ), .ZN(_04889_ ) );
NAND2_X1 _12643_ ( .A1(_04888_ ), .A2(_04889_ ), .ZN(_04890_ ) );
XNOR2_X1 _12644_ ( .A(_04890_ ), .B(_02543_ ), .ZN(_04891_ ) );
OAI21_X1 _12645_ ( .A(_04773_ ), .B1(_04186_ ), .B2(_04187_ ), .ZN(_04892_ ) );
NAND2_X1 _12646_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [6] ), .ZN(_04893_ ) );
AND2_X2 _12647_ ( .A1(_04892_ ), .A2(_04893_ ), .ZN(_04894_ ) );
OR2_X1 _12648_ ( .A1(_04894_ ), .A2(_04189_ ), .ZN(_04895_ ) );
NAND3_X1 _12649_ ( .A1(_04892_ ), .A2(_04189_ ), .A3(_04893_ ), .ZN(_04896_ ) );
AOI21_X1 _12650_ ( .A(_04891_ ), .B1(_04895_ ), .B2(_04896_ ), .ZN(_04897_ ) );
NAND2_X1 _12651_ ( .A1(_04234_ ), .A2(_04773_ ), .ZN(_04898_ ) );
OR2_X1 _12652_ ( .A1(_04772_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04899_ ) );
NAND2_X1 _12653_ ( .A1(_04898_ ), .A2(_04899_ ), .ZN(_04900_ ) );
INV_X1 _12654_ ( .A(_02589_ ), .ZN(_04901_ ) );
XNOR2_X1 _12655_ ( .A(_04900_ ), .B(_04901_ ), .ZN(_04902_ ) );
INV_X1 _12656_ ( .A(_04902_ ), .ZN(_04903_ ) );
NAND3_X1 _12657_ ( .A1(_04259_ ), .A2(_04774_ ), .A3(_04279_ ), .ZN(_04904_ ) );
NAND2_X1 _12658_ ( .A1(_02612_ ), .A2(fanout_net_6 ), .ZN(_04905_ ) );
NAND2_X1 _12659_ ( .A1(_04904_ ), .A2(_04905_ ), .ZN(_04906_ ) );
XNOR2_X1 _12660_ ( .A(_04906_ ), .B(_02611_ ), .ZN(_04907_ ) );
INV_X1 _12661_ ( .A(_04907_ ), .ZN(_04908_ ) );
NAND4_X1 _12662_ ( .A1(_04887_ ), .A2(_04897_ ), .A3(_04903_ ), .A4(_04908_ ), .ZN(_04909_ ) );
NAND3_X1 _12663_ ( .A1(_04892_ ), .A2(_02565_ ), .A3(_04893_ ), .ZN(_04910_ ) );
NOR2_X1 _12664_ ( .A1(_04891_ ), .A2(_04910_ ), .ZN(_04911_ ) );
NAND3_X1 _12665_ ( .A1(_04903_ ), .A2(_02611_ ), .A3(_04906_ ), .ZN(_04912_ ) );
OAI21_X1 _12666_ ( .A(_04912_ ), .B1(_04901_ ), .B2(_04900_ ), .ZN(_04913_ ) );
AOI221_X4 _12667_ ( .A(_04911_ ), .B1(_02543_ ), .B2(_04890_ ), .C1(_04913_ ), .C2(_04897_ ), .ZN(_04914_ ) );
AOI21_X1 _12668_ ( .A(_04859_ ), .B1(_04909_ ), .B2(_04914_ ), .ZN(_04915_ ) );
INV_X1 _12669_ ( .A(_04858_ ), .ZN(_04916_ ) );
AND2_X1 _12670_ ( .A1(_04842_ ), .A2(_04024_ ), .ZN(_04917_ ) );
NOR2_X1 _12671_ ( .A1(_04842_ ), .A2(_04024_ ), .ZN(_04918_ ) );
OAI211_X1 _12672_ ( .A(_02789_ ), .B(_04847_ ), .C1(_04917_ ), .C2(_04918_ ), .ZN(_04919_ ) );
OAI211_X1 _12673_ ( .A(_02812_ ), .B(_04841_ ), .C1(_04047_ ), .C2(fanout_net_6 ), .ZN(_04920_ ) );
AOI21_X1 _12674_ ( .A(_04916_ ), .B1(_04919_ ), .B2(_04920_ ), .ZN(_04921_ ) );
INV_X1 _12675_ ( .A(_04853_ ), .ZN(_04922_ ) );
NAND3_X1 _12676_ ( .A1(_04922_ ), .A2(_02742_ ), .A3(_04856_ ), .ZN(_04923_ ) );
INV_X1 _12677_ ( .A(_04852_ ), .ZN(_04924_ ) );
OAI21_X1 _12678_ ( .A(_04923_ ), .B1(_03916_ ), .B2(_04924_ ), .ZN(_04925_ ) );
OAI21_X1 _12679_ ( .A(_04839_ ), .B1(_04921_ ), .B2(_04925_ ), .ZN(_04926_ ) );
AOI22_X1 _12680_ ( .A1(_04829_ ), .A2(_04830_ ), .B1(_02667_ ), .B2(_02668_ ), .ZN(_04927_ ) );
INV_X1 _12681_ ( .A(_04836_ ), .ZN(_04928_ ) );
NOR3_X1 _12682_ ( .A1(_04832_ ), .A2(_04079_ ), .A3(_04928_ ), .ZN(_04929_ ) );
OAI21_X1 _12683_ ( .A(_04828_ ), .B1(_04927_ ), .B2(_04929_ ), .ZN(_04930_ ) );
INV_X1 _12684_ ( .A(_04821_ ), .ZN(_04931_ ) );
NAND3_X1 _12685_ ( .A1(_04931_ ), .A2(_02718_ ), .A3(_04824_ ), .ZN(_04932_ ) );
NAND2_X1 _12686_ ( .A1(_04820_ ), .A2(_02694_ ), .ZN(_04933_ ) );
NAND4_X1 _12687_ ( .A1(_04926_ ), .A2(_04930_ ), .A3(_04932_ ), .A4(_04933_ ), .ZN(_04934_ ) );
OR2_X1 _12688_ ( .A1(_04915_ ), .A2(_04934_ ), .ZN(_04935_ ) );
OR2_X1 _12689_ ( .A1(_04561_ ), .A2(fanout_net_6 ), .ZN(_04936_ ) );
NAND2_X1 _12690_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [22] ), .ZN(_04937_ ) );
AND2_X2 _12691_ ( .A1(_04936_ ), .A2(_04937_ ), .ZN(_04938_ ) );
XNOR2_X1 _12692_ ( .A(_04938_ ), .B(_02270_ ), .ZN(_04939_ ) );
OR2_X1 _12693_ ( .A1(_04536_ ), .A2(fanout_net_6 ), .ZN(_04940_ ) );
NAND2_X1 _12694_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [23] ), .ZN(_04941_ ) );
AND2_X1 _12695_ ( .A1(_04940_ ), .A2(_04941_ ), .ZN(_04942_ ) );
INV_X1 _12696_ ( .A(_02247_ ), .ZN(_04943_ ) );
NOR2_X1 _12697_ ( .A1(_04942_ ), .A2(_04943_ ), .ZN(_04944_ ) );
AND3_X1 _12698_ ( .A1(_04940_ ), .A2(_04943_ ), .A3(_04941_ ), .ZN(_04945_ ) );
NOR2_X2 _12699_ ( .A1(_04944_ ), .A2(_04945_ ), .ZN(_04946_ ) );
OR2_X1 _12700_ ( .A1(_04939_ ), .A2(_04946_ ), .ZN(_04947_ ) );
OAI21_X1 _12701_ ( .A(_04774_ ), .B1(_04507_ ), .B2(_04509_ ), .ZN(_04948_ ) );
NAND2_X1 _12702_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [21] ), .ZN(_04949_ ) );
AND2_X2 _12703_ ( .A1(_04948_ ), .A2(_04949_ ), .ZN(_04950_ ) );
XNOR2_X1 _12704_ ( .A(_04950_ ), .B(_04511_ ), .ZN(_04951_ ) );
NAND3_X1 _12705_ ( .A1(_04463_ ), .A2(_04774_ ), .A3(_04486_ ), .ZN(_04952_ ) );
NAND2_X1 _12706_ ( .A1(\ID_EX_typ [4] ), .A2(\ID_EX_imm [20] ), .ZN(_04953_ ) );
AND2_X1 _12707_ ( .A1(_04952_ ), .A2(_04953_ ), .ZN(_04954_ ) );
XNOR2_X1 _12708_ ( .A(_04954_ ), .B(_02294_ ), .ZN(_04955_ ) );
NOR3_X1 _12709_ ( .A1(_04947_ ), .A2(_04951_ ), .A3(_04955_ ), .ZN(_04956_ ) );
OR2_X1 _12710_ ( .A1(_04405_ ), .A2(\ID_EX_typ [4] ), .ZN(_04957_ ) );
NAND2_X1 _12711_ ( .A1(\ID_EX_typ [4] ), .A2(\ID_EX_imm [19] ), .ZN(_04958_ ) );
AND2_X1 _12712_ ( .A1(_04957_ ), .A2(_04958_ ), .ZN(_04959_ ) );
XNOR2_X1 _12713_ ( .A(_04959_ ), .B(_02370_ ), .ZN(_04960_ ) );
NAND3_X1 _12714_ ( .A1(_04358_ ), .A2(_04774_ ), .A3(_04380_ ), .ZN(_04961_ ) );
NAND2_X1 _12715_ ( .A1(\ID_EX_typ [4] ), .A2(\ID_EX_imm [18] ), .ZN(_04962_ ) );
AND2_X1 _12716_ ( .A1(_04961_ ), .A2(_04962_ ), .ZN(_04963_ ) );
XNOR2_X1 _12717_ ( .A(_04963_ ), .B(_02346_ ), .ZN(_04964_ ) );
OAI21_X1 _12718_ ( .A(_04774_ ), .B1(_04426_ ), .B2(_04428_ ), .ZN(_04965_ ) );
NAND2_X1 _12719_ ( .A1(\ID_EX_typ [4] ), .A2(\ID_EX_imm [17] ), .ZN(_04966_ ) );
AND2_X1 _12720_ ( .A1(_04965_ ), .A2(_04966_ ), .ZN(_04967_ ) );
XNOR2_X1 _12721_ ( .A(_04967_ ), .B(_02394_ ), .ZN(_04968_ ) );
NAND3_X1 _12722_ ( .A1(_04433_ ), .A2(_04774_ ), .A3(_04458_ ), .ZN(_04969_ ) );
NAND2_X1 _12723_ ( .A1(\ID_EX_typ [4] ), .A2(\ID_EX_imm [16] ), .ZN(_04970_ ) );
AND2_X1 _12724_ ( .A1(_04969_ ), .A2(_04970_ ), .ZN(_04971_ ) );
XNOR2_X1 _12725_ ( .A(_04971_ ), .B(_02417_ ), .ZN(_04972_ ) );
NOR4_X1 _12726_ ( .A1(_04960_ ), .A2(_04964_ ), .A3(_04968_ ), .A4(_04972_ ), .ZN(_04973_ ) );
AND3_X2 _12727_ ( .A1(_04935_ ), .A2(_04956_ ), .A3(_04973_ ), .ZN(_04974_ ) );
INV_X1 _12728_ ( .A(_04938_ ), .ZN(_04975_ ) );
NOR3_X1 _12729_ ( .A1(_04946_ ), .A2(_04538_ ), .A3(_04975_ ), .ZN(_04976_ ) );
NAND3_X1 _12730_ ( .A1(_04948_ ), .A2(_04511_ ), .A3(_04949_ ), .ZN(_04977_ ) );
INV_X1 _12731_ ( .A(_04511_ ), .ZN(_04978_ ) );
AND2_X1 _12732_ ( .A1(_04950_ ), .A2(_04978_ ), .ZN(_04979_ ) );
NOR2_X1 _12733_ ( .A1(_04950_ ), .A2(_04978_ ), .ZN(_04980_ ) );
OAI211_X1 _12734_ ( .A(_02294_ ), .B(_04954_ ), .C1(_04979_ ), .C2(_04980_ ), .ZN(_04981_ ) );
AOI21_X1 _12735_ ( .A(_04947_ ), .B1(_04977_ ), .B2(_04981_ ), .ZN(_04982_ ) );
AOI211_X1 _12736_ ( .A(_04976_ ), .B(_04982_ ), .C1(_02247_ ), .C2(_04942_ ), .ZN(_04983_ ) );
NOR2_X1 _12737_ ( .A1(_04960_ ), .A2(_04964_ ), .ZN(_04984_ ) );
NAND3_X1 _12738_ ( .A1(_04969_ ), .A2(_02417_ ), .A3(_04970_ ), .ZN(_04985_ ) );
NOR2_X1 _12739_ ( .A1(_04968_ ), .A2(_04985_ ), .ZN(_04986_ ) );
AND3_X1 _12740_ ( .A1(_04965_ ), .A2(_02394_ ), .A3(_04966_ ), .ZN(_04987_ ) );
OAI21_X1 _12741_ ( .A(_04984_ ), .B1(_04986_ ), .B2(_04987_ ), .ZN(_04988_ ) );
INV_X1 _12742_ ( .A(_04959_ ), .ZN(_04989_ ) );
OAI21_X1 _12743_ ( .A(_04988_ ), .B1(_04383_ ), .B2(_04989_ ), .ZN(_04990_ ) );
INV_X1 _12744_ ( .A(_04963_ ), .ZN(_04991_ ) );
NOR3_X1 _12745_ ( .A1(_04960_ ), .A2(_04357_ ), .A3(_04991_ ), .ZN(_04992_ ) );
OAI21_X1 _12746_ ( .A(_04956_ ), .B1(_04990_ ), .B2(_04992_ ), .ZN(_04993_ ) );
NAND2_X1 _12747_ ( .A1(_04983_ ), .A2(_04993_ ), .ZN(_04994_ ) );
OAI21_X1 _12748_ ( .A(_04817_ ), .B1(_04974_ ), .B2(_04994_ ), .ZN(_04995_ ) );
NAND2_X1 _12749_ ( .A1(_04813_ ), .A2(_02899_ ), .ZN(_04996_ ) );
OAI211_X1 _12750_ ( .A(_02876_ ), .B(_04806_ ), .C1(_04814_ ), .C2(_04815_ ), .ZN(_04997_ ) );
AOI21_X1 _12751_ ( .A(_04803_ ), .B1(_04996_ ), .B2(_04997_ ), .ZN(_04998_ ) );
INV_X1 _12752_ ( .A(_04790_ ), .ZN(_04999_ ) );
NOR3_X1 _12753_ ( .A1(_04801_ ), .A2(_04791_ ), .A3(_04999_ ), .ZN(_05000_ ) );
AOI21_X1 _12754_ ( .A(_04708_ ), .B1(_04796_ ), .B2(_04797_ ), .ZN(_05001_ ) );
NOR3_X1 _12755_ ( .A1(_04998_ ), .A2(_05000_ ), .A3(_05001_ ), .ZN(_05002_ ) );
AOI21_X1 _12756_ ( .A(_04786_ ), .B1(_04995_ ), .B2(_05002_ ), .ZN(_05003_ ) );
NAND3_X1 _12757_ ( .A1(_04612_ ), .A2(_04787_ ), .A3(_04632_ ), .ZN(_05004_ ) );
OR2_X1 _12758_ ( .A1(_04787_ ), .A2(\ID_EX_imm [31] ), .ZN(_05005_ ) );
NAND2_X1 _12759_ ( .A1(_05004_ ), .A2(_05005_ ), .ZN(_05006_ ) );
INV_X1 _12760_ ( .A(_02990_ ), .ZN(_05007_ ) );
XNOR2_X1 _12761_ ( .A(_05006_ ), .B(_05007_ ), .ZN(_05008_ ) );
INV_X1 _12762_ ( .A(_05008_ ), .ZN(_05009_ ) );
NAND3_X1 _12763_ ( .A1(_04635_ ), .A2(_04787_ ), .A3(_04655_ ), .ZN(_05010_ ) );
OR2_X1 _12764_ ( .A1(_04787_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05011_ ) );
NAND2_X1 _12765_ ( .A1(_05010_ ), .A2(_05011_ ), .ZN(_05012_ ) );
XNOR2_X1 _12766_ ( .A(_02963_ ), .B(_05012_ ), .ZN(_05013_ ) );
NOR2_X1 _12767_ ( .A1(_05009_ ), .A2(_05013_ ), .ZN(_05014_ ) );
NAND2_X1 _12768_ ( .A1(_05003_ ), .A2(_05014_ ), .ZN(_05015_ ) );
NOR2_X1 _12769_ ( .A1(_02963_ ), .A2(_05012_ ), .ZN(_05016_ ) );
AND2_X1 _12770_ ( .A1(_05008_ ), .A2(_05016_ ), .ZN(_05017_ ) );
INV_X1 _12771_ ( .A(_05006_ ), .ZN(_05018_ ) );
INV_X1 _12772_ ( .A(_04777_ ), .ZN(_05019_ ) );
OAI211_X1 _12773_ ( .A(_02167_ ), .B(_05019_ ), .C1(_04784_ ), .C2(_04785_ ), .ZN(_05020_ ) );
OAI21_X1 _12774_ ( .A(_05020_ ), .B1(_02940_ ), .B2(_04783_ ), .ZN(_05021_ ) );
AOI221_X4 _12775_ ( .A(_05017_ ), .B1(_05007_ ), .B2(_05018_ ), .C1(_05021_ ), .C2(_05014_ ), .ZN(_05022_ ) );
AOI21_X1 _12776_ ( .A(_04771_ ), .B1(_05015_ ), .B2(_05022_ ), .ZN(_05023_ ) );
AND2_X1 _12777_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_5 ), .ZN(_05024_ ) );
AND2_X2 _12778_ ( .A1(_05024_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_05025_ ) );
INV_X2 _12779_ ( .A(_05025_ ), .ZN(_05026_ ) );
NAND2_X1 _12780_ ( .A1(_04256_ ), .A2(_02464_ ), .ZN(_05027_ ) );
INV_X2 _12781_ ( .A(_04257_ ), .ZN(_05028_ ) );
AOI21_X1 _12782_ ( .A(_04353_ ), .B1(_02488_ ), .B2(_02468_ ), .ZN(_05029_ ) );
OAI21_X4 _12783_ ( .A(_05027_ ), .B1(_05028_ ), .B2(_05029_ ), .ZN(_05030_ ) );
NAND2_X1 _12784_ ( .A1(_05030_ ), .A2(_04306_ ), .ZN(_05031_ ) );
INV_X1 _12785_ ( .A(_04304_ ), .ZN(_05032_ ) );
AOI22_X1 _12786_ ( .A1(_05031_ ), .A2(_05032_ ), .B1(_02520_ ), .B2(_04328_ ), .ZN(_05033_ ) );
NOR2_X1 _12787_ ( .A1(_02520_ ), .A2(_04328_ ), .ZN(_05034_ ) );
OR2_X2 _12788_ ( .A1(_05033_ ), .A2(_05034_ ), .ZN(_05035_ ) );
NAND4_X4 _12789_ ( .A1(_05035_ ), .A2(_04214_ ), .A3(_04235_ ), .A4(_04281_ ), .ZN(_05036_ ) );
AND3_X1 _12790_ ( .A1(_04213_ ), .A2(_02565_ ), .A3(_04188_ ), .ZN(_05037_ ) );
NAND3_X1 _12791_ ( .A1(_04235_ ), .A2(_02611_ ), .A3(_04280_ ), .ZN(_05038_ ) );
OAI21_X1 _12792_ ( .A(_05038_ ), .B1(_04901_ ), .B2(_04234_ ), .ZN(_05039_ ) );
AOI221_X2 _12793_ ( .A(_05037_ ), .B1(_02543_ ), .B2(_04212_ ), .C1(_05039_ ), .C2(_04214_ ), .ZN(_05040_ ) );
AND2_X4 _12794_ ( .A1(_05036_ ), .A2(_05040_ ), .ZN(_05041_ ) );
INV_X4 _12795_ ( .A(_05041_ ), .ZN(_05042_ ) );
NAND2_X4 _12796_ ( .A1(_05042_ ), .A2(_04167_ ), .ZN(_05043_ ) );
AND3_X1 _12797_ ( .A1(_04133_ ), .A2(_02718_ ), .A3(_04164_ ), .ZN(_05044_ ) );
NAND2_X1 _12798_ ( .A1(_04106_ ), .A2(_02647_ ), .ZN(_05045_ ) );
NOR3_X1 _12799_ ( .A1(_04076_ ), .A2(_04077_ ), .A3(_05045_ ), .ZN(_05046_ ) );
OR2_X1 _12800_ ( .A1(_05046_ ), .A2(_04076_ ), .ZN(_05047_ ) );
NAND3_X1 _12801_ ( .A1(_05047_ ), .A2(_04133_ ), .A3(_04165_ ), .ZN(_05048_ ) );
AND2_X1 _12802_ ( .A1(_04021_ ), .A2(_02789_ ), .ZN(_05049_ ) );
AOI21_X1 _12803_ ( .A(_05049_ ), .B1(_02812_ ), .B2(_04047_ ), .ZN(_05050_ ) );
NOR2_X1 _12804_ ( .A1(_04047_ ), .A2(_02812_ ), .ZN(_05051_ ) );
NOR2_X1 _12805_ ( .A1(_05050_ ), .A2(_05051_ ), .ZN(_05052_ ) );
AND2_X1 _12806_ ( .A1(_05052_ ), .A2(_03993_ ), .ZN(_05053_ ) );
AND3_X1 _12807_ ( .A1(_02765_ ), .A2(_03963_ ), .A3(_03928_ ), .ZN(_05054_ ) );
AND3_X1 _12808_ ( .A1(_03965_ ), .A2(_02742_ ), .A3(_03991_ ), .ZN(_05055_ ) );
NOR3_X4 _12809_ ( .A1(_05053_ ), .A2(_05054_ ), .A3(_05055_ ), .ZN(_05056_ ) );
OAI21_X1 _12810_ ( .A(_05048_ ), .B1(_05056_ ), .B2(_04166_ ), .ZN(_05057_ ) );
AOI211_X2 _12811_ ( .A(_05044_ ), .B(_05057_ ), .C1(_02694_ ), .C2(_04132_ ), .ZN(_05058_ ) );
AND2_X1 _12812_ ( .A1(_05043_ ), .A2(_05058_ ), .ZN(_05059_ ) );
INV_X1 _12813_ ( .A(_04762_ ), .ZN(_05060_ ) );
OR2_X4 _12814_ ( .A1(_05059_ ), .A2(_05060_ ), .ZN(_05061_ ) );
NOR2_X1 _12815_ ( .A1(_04778_ ), .A2(_04609_ ), .ZN(_05062_ ) );
NOR2_X1 _12816_ ( .A1(_04586_ ), .A2(_05062_ ), .ZN(_05063_ ) );
NOR2_X1 _12817_ ( .A1(_05063_ ), .A2(_04587_ ), .ZN(_05064_ ) );
AND3_X1 _12818_ ( .A1(_05064_ ), .A2(_04634_ ), .A3(_04658_ ), .ZN(_05065_ ) );
NOR2_X1 _12819_ ( .A1(_02963_ ), .A2(_04656_ ), .ZN(_05066_ ) );
NAND2_X1 _12820_ ( .A1(_04634_ ), .A2(_05066_ ), .ZN(_05067_ ) );
NOR2_X1 _12821_ ( .A1(_04733_ ), .A2(_04807_ ), .ZN(_05068_ ) );
NAND3_X1 _12822_ ( .A1(_05068_ ), .A2(_04758_ ), .A3(_04757_ ), .ZN(_05069_ ) );
NAND2_X1 _12823_ ( .A1(_05069_ ), .A2(_04758_ ), .ZN(_05070_ ) );
NAND4_X1 _12824_ ( .A1(_05070_ ), .A2(_04709_ ), .A3(_04710_ ), .A4(_04685_ ), .ZN(_05071_ ) );
NOR2_X1 _12825_ ( .A1(_04684_ ), .A2(_04791_ ), .ZN(_05072_ ) );
NAND3_X1 _12826_ ( .A1(_04709_ ), .A2(_04710_ ), .A3(_05072_ ), .ZN(_05073_ ) );
AND3_X1 _12827_ ( .A1(_05071_ ), .A2(_04709_ ), .A3(_05073_ ), .ZN(_05074_ ) );
INV_X1 _12828_ ( .A(_04659_ ), .ZN(_05075_ ) );
OAI221_X1 _12829_ ( .A(_05067_ ), .B1(_05007_ ), .B2(_04633_ ), .C1(_05074_ ), .C2(_05075_ ), .ZN(_05076_ ) );
AND2_X1 _12830_ ( .A1(_04459_ ), .A2(_02417_ ), .ZN(_05077_ ) );
NAND2_X1 _12831_ ( .A1(_04431_ ), .A2(_05077_ ), .ZN(_05078_ ) );
AND2_X1 _12832_ ( .A1(_04429_ ), .A2(_02394_ ), .ZN(_05079_ ) );
INV_X1 _12833_ ( .A(_05079_ ), .ZN(_05080_ ) );
NAND2_X1 _12834_ ( .A1(_05078_ ), .A2(_05080_ ), .ZN(_05081_ ) );
AND2_X1 _12835_ ( .A1(_04407_ ), .A2(_05081_ ), .ZN(_05082_ ) );
AND3_X1 _12836_ ( .A1(_02370_ ), .A2(_04404_ ), .A3(_04385_ ), .ZN(_05083_ ) );
AND3_X1 _12837_ ( .A1(_04406_ ), .A2(_02346_ ), .A3(_04381_ ), .ZN(_05084_ ) );
NOR3_X1 _12838_ ( .A1(_05082_ ), .A2(_05083_ ), .A3(_05084_ ), .ZN(_05085_ ) );
NOR2_X1 _12839_ ( .A1(_05085_ ), .A2(_04563_ ), .ZN(_05086_ ) );
AND2_X1 _12840_ ( .A1(_04487_ ), .A2(_02294_ ), .ZN(_05087_ ) );
NOR2_X1 _12841_ ( .A1(_04512_ ), .A2(_05087_ ), .ZN(_05088_ ) );
NOR2_X1 _12842_ ( .A1(_05088_ ), .A2(_04513_ ), .ZN(_05089_ ) );
AND3_X1 _12843_ ( .A1(_05089_ ), .A2(_04537_ ), .A3(_04562_ ), .ZN(_05090_ ) );
OR2_X1 _12844_ ( .A1(_05086_ ), .A2(_05090_ ), .ZN(_05091_ ) );
AND2_X1 _12845_ ( .A1(_02247_ ), .A2(_04536_ ), .ZN(_05092_ ) );
AND2_X1 _12846_ ( .A1(_04561_ ), .A2(_02270_ ), .ZN(_05093_ ) );
AND2_X1 _12847_ ( .A1(_04537_ ), .A2(_05093_ ), .ZN(_05094_ ) );
NOR3_X1 _12848_ ( .A1(_05091_ ), .A2(_05092_ ), .A3(_05094_ ), .ZN(_05095_ ) );
INV_X1 _12849_ ( .A(_05095_ ), .ZN(_05096_ ) );
AOI211_X1 _12850_ ( .A(_05065_ ), .B(_05076_ ), .C1(_05096_ ), .C2(_04761_ ), .ZN(_05097_ ) );
AOI21_X1 _12851_ ( .A(_05026_ ), .B1(_05061_ ), .B2(_05097_ ), .ZN(_05098_ ) );
AND2_X2 _12852_ ( .A1(_04764_ ), .A2(\ID_EX_typ [2] ), .ZN(_05099_ ) );
AND3_X1 _12853_ ( .A1(_05061_ ), .A2(_05097_ ), .A3(_05099_ ), .ZN(_05100_ ) );
OR4_X2 _12854_ ( .A1(_05023_ ), .A2(_04765_ ), .A3(_05098_ ), .A4(_05100_ ), .ZN(_05101_ ) );
AND2_X1 _12855_ ( .A1(_05015_ ), .A2(_05022_ ), .ZN(_05102_ ) );
AND3_X1 _12856_ ( .A1(_05102_ ), .A2(\ID_EX_typ [2] ), .A3(_03913_ ), .ZN(_05103_ ) );
OAI221_X2 _12857_ ( .A(_03915_ ), .B1(_04763_ ), .B2(_04766_ ), .C1(_05101_ ), .C2(_05103_ ), .ZN(_05104_ ) );
NAND4_X1 _12858_ ( .A1(_04167_ ), .A2(_04214_ ), .A3(_04235_ ), .A4(_04355_ ), .ZN(_05105_ ) );
OAI21_X1 _12859_ ( .A(_03914_ ), .B1(_05060_ ), .B2(_05105_ ), .ZN(_05106_ ) );
AOI21_X1 _12860_ ( .A(_03912_ ), .B1(_05104_ ), .B2(_05106_ ), .ZN(_05107_ ) );
XOR2_X1 _12861_ ( .A(\ID_EX_pc [25] ), .B(\ID_EX_imm [25] ), .Z(_05108_ ) );
XOR2_X1 _12862_ ( .A(\ID_EX_pc [24] ), .B(\ID_EX_imm [24] ), .Z(_05109_ ) );
XOR2_X1 _12863_ ( .A(\ID_EX_pc [4] ), .B(\ID_EX_imm [4] ), .Z(_05110_ ) );
INV_X1 _12864_ ( .A(_05110_ ), .ZN(_05111_ ) );
XOR2_X1 _12865_ ( .A(\ID_EX_pc [2] ), .B(\ID_EX_imm [2] ), .Z(_05112_ ) );
XOR2_X1 _12866_ ( .A(\ID_EX_pc [1] ), .B(\ID_EX_imm [1] ), .Z(_05113_ ) );
AND2_X1 _12867_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_05114_ ) );
AND2_X1 _12868_ ( .A1(_05113_ ), .A2(_05114_ ), .ZN(_05115_ ) );
AND2_X1 _12869_ ( .A1(\ID_EX_pc [1] ), .A2(\ID_EX_imm [1] ), .ZN(_05116_ ) );
OAI21_X1 _12870_ ( .A(_05112_ ), .B1(_05115_ ), .B2(_05116_ ), .ZN(_05117_ ) );
NAND2_X1 _12871_ ( .A1(\ID_EX_pc [2] ), .A2(\ID_EX_imm [2] ), .ZN(_05118_ ) );
NAND2_X1 _12872_ ( .A1(_05117_ ), .A2(_05118_ ), .ZN(_05119_ ) );
OAI21_X1 _12873_ ( .A(_05119_ ), .B1(\ID_EX_pc [3] ), .B2(\ID_EX_imm [3] ), .ZN(_05120_ ) );
AND2_X1 _12874_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_05121_ ) );
INV_X1 _12875_ ( .A(_05121_ ), .ZN(_05122_ ) );
AOI21_X1 _12876_ ( .A(_05111_ ), .B1(_05120_ ), .B2(_05122_ ), .ZN(_05123_ ) );
AND2_X1 _12877_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_05124_ ) );
AND2_X1 _12878_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_05125_ ) );
NOR3_X1 _12879_ ( .A1(_05123_ ), .A2(_05124_ ), .A3(_05125_ ), .ZN(_05126_ ) );
NOR2_X1 _12880_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_05127_ ) );
NOR2_X1 _12881_ ( .A1(_05126_ ), .A2(_05127_ ), .ZN(_05128_ ) );
XOR2_X1 _12882_ ( .A(\ID_EX_pc [6] ), .B(\ID_EX_imm [6] ), .Z(_05129_ ) );
NAND2_X1 _12883_ ( .A1(_05128_ ), .A2(_05129_ ), .ZN(_05130_ ) );
NAND2_X1 _12884_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_05131_ ) );
NAND2_X1 _12885_ ( .A1(_05130_ ), .A2(_05131_ ), .ZN(_05132_ ) );
OAI21_X1 _12886_ ( .A(_05132_ ), .B1(\ID_EX_pc [7] ), .B2(\ID_EX_imm [7] ), .ZN(_05133_ ) );
AND2_X1 _12887_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_05134_ ) );
INV_X1 _12888_ ( .A(_05134_ ), .ZN(_05135_ ) );
NAND2_X1 _12889_ ( .A1(_05133_ ), .A2(_05135_ ), .ZN(_05136_ ) );
XOR2_X1 _12890_ ( .A(\ID_EX_pc [11] ), .B(\ID_EX_imm [11] ), .Z(_05137_ ) );
XOR2_X1 _12891_ ( .A(\ID_EX_pc [10] ), .B(\ID_EX_imm [10] ), .Z(_05138_ ) );
AND2_X1 _12892_ ( .A1(_05137_ ), .A2(_05138_ ), .ZN(_05139_ ) );
XOR2_X1 _12893_ ( .A(\ID_EX_pc [8] ), .B(\ID_EX_imm [8] ), .Z(_05140_ ) );
XOR2_X1 _12894_ ( .A(\ID_EX_pc [9] ), .B(\ID_EX_imm [9] ), .Z(_05141_ ) );
AND2_X1 _12895_ ( .A1(_05140_ ), .A2(_05141_ ), .ZN(_05142_ ) );
AND3_X1 _12896_ ( .A1(_05136_ ), .A2(_05139_ ), .A3(_05142_ ), .ZN(_05143_ ) );
AND2_X1 _12897_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_05144_ ) );
AND2_X1 _12898_ ( .A1(_05137_ ), .A2(_05144_ ), .ZN(_05145_ ) );
AOI21_X1 _12899_ ( .A(_05145_ ), .B1(\ID_EX_pc [11] ), .B2(\ID_EX_imm [11] ), .ZN(_05146_ ) );
AND2_X1 _12900_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_imm [8] ), .ZN(_05147_ ) );
AND2_X1 _12901_ ( .A1(_05141_ ), .A2(_05147_ ), .ZN(_05148_ ) );
AOI21_X1 _12902_ ( .A(_05148_ ), .B1(\ID_EX_pc [9] ), .B2(\ID_EX_imm [9] ), .ZN(_05149_ ) );
INV_X1 _12903_ ( .A(_05139_ ), .ZN(_05150_ ) );
OAI21_X1 _12904_ ( .A(_05146_ ), .B1(_05149_ ), .B2(_05150_ ), .ZN(_05151_ ) );
OR2_X1 _12905_ ( .A1(_05143_ ), .A2(_05151_ ), .ZN(_05152_ ) );
XOR2_X1 _12906_ ( .A(\ID_EX_pc [15] ), .B(\ID_EX_imm [15] ), .Z(_05153_ ) );
XOR2_X1 _12907_ ( .A(\ID_EX_pc [14] ), .B(\ID_EX_imm [14] ), .Z(_05154_ ) );
XOR2_X1 _12908_ ( .A(\ID_EX_pc [12] ), .B(\ID_EX_imm [12] ), .Z(_05155_ ) );
XOR2_X1 _12909_ ( .A(\ID_EX_pc [13] ), .B(\ID_EX_imm [13] ), .Z(_05156_ ) );
AND2_X1 _12910_ ( .A1(_05155_ ), .A2(_05156_ ), .ZN(_05157_ ) );
NAND4_X1 _12911_ ( .A1(_05152_ ), .A2(_05153_ ), .A3(_05154_ ), .A4(_05157_ ), .ZN(_05158_ ) );
AND2_X1 _12912_ ( .A1(\ID_EX_pc [12] ), .A2(\ID_EX_imm [12] ), .ZN(_05159_ ) );
AND2_X1 _12913_ ( .A1(_05156_ ), .A2(_05159_ ), .ZN(_05160_ ) );
AOI21_X1 _12914_ ( .A(_05160_ ), .B1(\ID_EX_pc [13] ), .B2(\ID_EX_imm [13] ), .ZN(_05161_ ) );
NAND2_X1 _12915_ ( .A1(_05153_ ), .A2(_05154_ ), .ZN(_05162_ ) );
NOR2_X1 _12916_ ( .A1(_05161_ ), .A2(_05162_ ), .ZN(_05163_ ) );
AND2_X1 _12917_ ( .A1(\ID_EX_pc [15] ), .A2(\ID_EX_imm [15] ), .ZN(_05164_ ) );
AND2_X1 _12918_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_05165_ ) );
AND2_X1 _12919_ ( .A1(_05153_ ), .A2(_05165_ ), .ZN(_05166_ ) );
NOR3_X1 _12920_ ( .A1(_05163_ ), .A2(_05164_ ), .A3(_05166_ ), .ZN(_05167_ ) );
NAND2_X1 _12921_ ( .A1(_05158_ ), .A2(_05167_ ), .ZN(_05168_ ) );
XOR2_X1 _12922_ ( .A(\ID_EX_pc [23] ), .B(\ID_EX_imm [23] ), .Z(_05169_ ) );
XOR2_X1 _12923_ ( .A(\ID_EX_pc [22] ), .B(\ID_EX_imm [22] ), .Z(_05170_ ) );
AND2_X1 _12924_ ( .A1(_05169_ ), .A2(_05170_ ), .ZN(_05171_ ) );
XOR2_X1 _12925_ ( .A(\ID_EX_pc [21] ), .B(\ID_EX_imm [21] ), .Z(_05172_ ) );
XOR2_X1 _12926_ ( .A(\ID_EX_pc [20] ), .B(\ID_EX_imm [20] ), .Z(_05173_ ) );
AND2_X1 _12927_ ( .A1(_05172_ ), .A2(_05173_ ), .ZN(_05174_ ) );
AND2_X1 _12928_ ( .A1(_05171_ ), .A2(_05174_ ), .ZN(_05175_ ) );
XOR2_X1 _12929_ ( .A(\ID_EX_pc [19] ), .B(\ID_EX_imm [19] ), .Z(_05176_ ) );
XOR2_X1 _12930_ ( .A(\ID_EX_pc [18] ), .B(\ID_EX_imm [18] ), .Z(_05177_ ) );
AND2_X1 _12931_ ( .A1(_05176_ ), .A2(_05177_ ), .ZN(_05178_ ) );
XOR2_X1 _12932_ ( .A(\ID_EX_pc [16] ), .B(\ID_EX_imm [16] ), .Z(_05179_ ) );
XOR2_X1 _12933_ ( .A(\ID_EX_pc [17] ), .B(\ID_EX_imm [17] ), .Z(_05180_ ) );
AND2_X1 _12934_ ( .A1(_05179_ ), .A2(_05180_ ), .ZN(_05181_ ) );
AND2_X1 _12935_ ( .A1(_05178_ ), .A2(_05181_ ), .ZN(_05182_ ) );
AND3_X1 _12936_ ( .A1(_05168_ ), .A2(_05175_ ), .A3(_05182_ ), .ZN(_05183_ ) );
AND2_X1 _12937_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_05184_ ) );
AND2_X1 _12938_ ( .A1(_05176_ ), .A2(_05184_ ), .ZN(_05185_ ) );
AOI21_X1 _12939_ ( .A(_05185_ ), .B1(\ID_EX_pc [19] ), .B2(\ID_EX_imm [19] ), .ZN(_05186_ ) );
AND2_X1 _12940_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_05187_ ) );
AND2_X1 _12941_ ( .A1(_05180_ ), .A2(_05187_ ), .ZN(_05188_ ) );
AOI21_X1 _12942_ ( .A(_05188_ ), .B1(\ID_EX_pc [17] ), .B2(\ID_EX_imm [17] ), .ZN(_05189_ ) );
INV_X1 _12943_ ( .A(_05178_ ), .ZN(_05190_ ) );
OAI21_X1 _12944_ ( .A(_05186_ ), .B1(_05189_ ), .B2(_05190_ ), .ZN(_05191_ ) );
NAND2_X1 _12945_ ( .A1(_05191_ ), .A2(_05175_ ), .ZN(_05192_ ) );
AND2_X1 _12946_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_05193_ ) );
AND2_X1 _12947_ ( .A1(_05169_ ), .A2(_05193_ ), .ZN(_05194_ ) );
AOI21_X1 _12948_ ( .A(_05194_ ), .B1(\ID_EX_pc [23] ), .B2(\ID_EX_imm [23] ), .ZN(_05195_ ) );
INV_X1 _12949_ ( .A(_05171_ ), .ZN(_05196_ ) );
AND3_X1 _12950_ ( .A1(_05172_ ), .A2(\ID_EX_pc [20] ), .A3(\ID_EX_imm [20] ), .ZN(_05197_ ) );
AOI21_X1 _12951_ ( .A(_05197_ ), .B1(\ID_EX_pc [21] ), .B2(\ID_EX_imm [21] ), .ZN(_05198_ ) );
OAI211_X1 _12952_ ( .A(_05192_ ), .B(_05195_ ), .C1(_05196_ ), .C2(_05198_ ), .ZN(_05199_ ) );
OAI211_X1 _12953_ ( .A(_05108_ ), .B(_05109_ ), .C1(_05183_ ), .C2(_05199_ ), .ZN(_05200_ ) );
AND2_X1 _12954_ ( .A1(\ID_EX_pc [24] ), .A2(\ID_EX_imm [24] ), .ZN(_05201_ ) );
AND2_X1 _12955_ ( .A1(_05108_ ), .A2(_05201_ ), .ZN(_05202_ ) );
AOI21_X1 _12956_ ( .A(_05202_ ), .B1(\ID_EX_pc [25] ), .B2(\ID_EX_imm [25] ), .ZN(_05203_ ) );
AND2_X1 _12957_ ( .A1(_05200_ ), .A2(_05203_ ), .ZN(_05204_ ) );
INV_X1 _12958_ ( .A(_05204_ ), .ZN(_05205_ ) );
XOR2_X1 _12959_ ( .A(\ID_EX_pc [27] ), .B(\ID_EX_imm [27] ), .Z(_05206_ ) );
XOR2_X1 _12960_ ( .A(\ID_EX_pc [26] ), .B(\ID_EX_imm [26] ), .Z(_05207_ ) );
AND3_X1 _12961_ ( .A1(_05205_ ), .A2(_05206_ ), .A3(_05207_ ), .ZN(_05208_ ) );
NAND3_X1 _12962_ ( .A1(_05206_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_imm [26] ), .ZN(_05209_ ) );
INV_X1 _12963_ ( .A(\ID_EX_pc [27] ), .ZN(_05210_ ) );
OAI21_X1 _12964_ ( .A(_05209_ ), .B1(_05210_ ), .B2(_02200_ ), .ZN(_05211_ ) );
NOR2_X1 _12965_ ( .A1(_05208_ ), .A2(_05211_ ), .ZN(_05212_ ) );
AND2_X1 _12966_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_05213_ ) );
NOR2_X1 _12967_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_05214_ ) );
NOR3_X1 _12968_ ( .A1(_05212_ ), .A2(_05213_ ), .A3(_05214_ ), .ZN(_05215_ ) );
NOR2_X1 _12969_ ( .A1(_05215_ ), .A2(_05213_ ), .ZN(_05216_ ) );
INV_X1 _12970_ ( .A(\ID_EX_pc [29] ), .ZN(_05217_ ) );
OAI21_X1 _12971_ ( .A(_05216_ ), .B1(_05217_ ), .B2(_02935_ ), .ZN(_05218_ ) );
NAND2_X1 _12972_ ( .A1(_05217_ ), .A2(_02935_ ), .ZN(_05219_ ) );
NAND2_X1 _12973_ ( .A1(_05218_ ), .A2(_05219_ ), .ZN(_05220_ ) );
XNOR2_X1 _12974_ ( .A(\ID_EX_pc [30] ), .B(\ID_EX_imm [30] ), .ZN(_05221_ ) );
XOR2_X1 _12975_ ( .A(_05220_ ), .B(_05221_ ), .Z(_05222_ ) );
AND2_X4 _12976_ ( .A1(_05104_ ), .A2(_05106_ ), .ZN(_05223_ ) );
BUF_X8 _12977_ ( .A(_05223_ ), .Z(_05224_ ) );
AOI211_X1 _12978_ ( .A(\ID_EX_typ [3] ), .B(_05107_ ), .C1(_05222_ ), .C2(_05224_ ), .ZN(_05225_ ) );
INV_X1 _12979_ ( .A(\EX_LS_result_csreg_mem [30] ), .ZN(_05226_ ) );
INV_X1 _12980_ ( .A(\ID_EX_csr [9] ), .ZN(_05227_ ) );
INV_X1 _12981_ ( .A(\ID_EX_csr [8] ), .ZN(_05228_ ) );
OR3_X1 _12982_ ( .A1(_05227_ ), .A2(_05228_ ), .A3(\ID_EX_csr [11] ), .ZN(_05229_ ) );
NOR2_X1 _12983_ ( .A1(_05229_ ), .A2(\ID_EX_csr [10] ), .ZN(_05230_ ) );
NOR2_X1 _12984_ ( .A1(\ID_EX_csr [7] ), .A2(\ID_EX_csr [6] ), .ZN(_05231_ ) );
NOR2_X1 _12985_ ( .A1(\ID_EX_csr [5] ), .A2(\ID_EX_csr [4] ), .ZN(_05232_ ) );
AND3_X1 _12986_ ( .A1(_05230_ ), .A2(_05231_ ), .A3(_05232_ ), .ZN(_05233_ ) );
BUF_X4 _12987_ ( .A(_05233_ ), .Z(_05234_ ) );
BUF_X4 _12988_ ( .A(_05234_ ), .Z(_05235_ ) );
BUF_X2 _12989_ ( .A(_05235_ ), .Z(_05236_ ) );
INV_X1 _12990_ ( .A(\ID_EX_csr [3] ), .ZN(_05237_ ) );
INV_X1 _12991_ ( .A(\ID_EX_csr [2] ), .ZN(_05238_ ) );
NAND2_X1 _12992_ ( .A1(_05237_ ), .A2(_05238_ ), .ZN(_05239_ ) );
NOR3_X1 _12993_ ( .A1(_05239_ ), .A2(\ID_EX_csr [1] ), .A3(\ID_EX_csr [0] ), .ZN(_05240_ ) );
BUF_X4 _12994_ ( .A(_05240_ ), .Z(_05241_ ) );
BUF_X4 _12995_ ( .A(_05241_ ), .Z(_05242_ ) );
NAND3_X1 _12996_ ( .A1(_05236_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_05242_ ), .ZN(_05243_ ) );
INV_X1 _12997_ ( .A(\ID_EX_csr [7] ), .ZN(_05244_ ) );
AND3_X1 _12998_ ( .A1(_05232_ ), .A2(_05244_ ), .A3(\ID_EX_csr [6] ), .ZN(_05245_ ) );
AND2_X2 _12999_ ( .A1(_05230_ ), .A2(_05245_ ), .ZN(_05246_ ) );
BUF_X4 _13000_ ( .A(_05246_ ), .Z(_05247_ ) );
BUF_X4 _13001_ ( .A(_05247_ ), .Z(_05248_ ) );
INV_X1 _13002_ ( .A(\ID_EX_csr [1] ), .ZN(_05249_ ) );
NAND2_X1 _13003_ ( .A1(_05249_ ), .A2(\ID_EX_csr [0] ), .ZN(_05250_ ) );
NOR2_X1 _13004_ ( .A1(_05239_ ), .A2(_05250_ ), .ZN(_05251_ ) );
BUF_X4 _13005_ ( .A(_05251_ ), .Z(_05252_ ) );
BUF_X4 _13006_ ( .A(_05252_ ), .Z(_05253_ ) );
NAND3_X1 _13007_ ( .A1(_05248_ ), .A2(\mepc [30] ), .A3(_05253_ ), .ZN(_05254_ ) );
NAND3_X1 _13008_ ( .A1(_05237_ ), .A2(_05238_ ), .A3(\ID_EX_csr [1] ), .ZN(_05255_ ) );
NOR2_X1 _13009_ ( .A1(_05255_ ), .A2(\ID_EX_csr [0] ), .ZN(_05256_ ) );
BUF_X2 _13010_ ( .A(_05256_ ), .Z(_05257_ ) );
NAND3_X1 _13011_ ( .A1(_05248_ ), .A2(\mycsreg.CSReg[3][30] ), .A3(_05257_ ), .ZN(_05258_ ) );
NAND3_X1 _13012_ ( .A1(_05243_ ), .A2(_05254_ ), .A3(_05258_ ), .ZN(_05259_ ) );
BUF_X2 _13013_ ( .A(_05234_ ), .Z(_05260_ ) );
NOR3_X1 _13014_ ( .A1(_05250_ ), .A2(\ID_EX_csr [3] ), .A3(_05238_ ), .ZN(_05261_ ) );
BUF_X2 _13015_ ( .A(_05261_ ), .Z(_05262_ ) );
AND3_X1 _13016_ ( .A1(_05260_ ), .A2(\mtvec [30] ), .A3(_05262_ ), .ZN(_05263_ ) );
INV_X1 _13017_ ( .A(\ID_EX_csr [5] ), .ZN(_05264_ ) );
AND4_X1 _13018_ ( .A1(\ID_EX_csr [10] ), .A2(_05264_ ), .A3(\ID_EX_csr [4] ), .A4(\ID_EX_csr [11] ), .ZN(_05265_ ) );
AND2_X1 _13019_ ( .A1(\ID_EX_csr [9] ), .A2(\ID_EX_csr [8] ), .ZN(_05266_ ) );
AND3_X1 _13020_ ( .A1(_05265_ ), .A2(_05266_ ), .A3(_05231_ ), .ZN(_05267_ ) );
AND2_X2 _13021_ ( .A1(_05267_ ), .A2(_05251_ ), .ZN(_05268_ ) );
NOR3_X1 _13022_ ( .A1(_05259_ ), .A2(_05263_ ), .A3(_05268_ ), .ZN(_05269_ ) );
AOI22_X1 _13023_ ( .A1(\EX_LS_dest_csreg_mem [9] ), .A2(_05227_ ), .B1(_05228_ ), .B2(\EX_LS_dest_csreg_mem [8] ), .ZN(_05270_ ) );
XNOR2_X1 _13024_ ( .A(\EX_LS_dest_csreg_mem [4] ), .B(\ID_EX_csr [4] ), .ZN(_05271_ ) );
XNOR2_X1 _13025_ ( .A(\EX_LS_dest_csreg_mem [3] ), .B(\ID_EX_csr [3] ), .ZN(_05272_ ) );
INV_X1 _13026_ ( .A(\EX_LS_dest_csreg_mem [9] ), .ZN(_05273_ ) );
INV_X1 _13027_ ( .A(\EX_LS_dest_csreg_mem [8] ), .ZN(_05274_ ) );
AOI22_X1 _13028_ ( .A1(_05273_ ), .A2(\ID_EX_csr [9] ), .B1(_05274_ ), .B2(\ID_EX_csr [8] ), .ZN(_05275_ ) );
AND4_X1 _13029_ ( .A1(_05270_ ), .A2(_05271_ ), .A3(_05272_ ), .A4(_05275_ ), .ZN(_05276_ ) );
XNOR2_X1 _13030_ ( .A(\EX_LS_dest_csreg_mem [10] ), .B(\ID_EX_csr [10] ), .ZN(_05277_ ) );
XNOR2_X1 _13031_ ( .A(\EX_LS_dest_csreg_mem [7] ), .B(\ID_EX_csr [7] ), .ZN(_05278_ ) );
AND3_X1 _13032_ ( .A1(_05276_ ), .A2(_05277_ ), .A3(_05278_ ), .ZN(_05279_ ) );
XNOR2_X1 _13033_ ( .A(\EX_LS_dest_csreg_mem [5] ), .B(\ID_EX_csr [5] ), .ZN(_05280_ ) );
XNOR2_X1 _13034_ ( .A(fanout_net_3 ), .B(\ID_EX_csr [0] ), .ZN(_05281_ ) );
XNOR2_X1 _13035_ ( .A(\EX_LS_dest_csreg_mem [11] ), .B(\ID_EX_csr [11] ), .ZN(_05282_ ) );
XNOR2_X1 _13036_ ( .A(\EX_LS_dest_csreg_mem [6] ), .B(\ID_EX_csr [6] ), .ZN(_05283_ ) );
NAND4_X1 _13037_ ( .A1(_05280_ ), .A2(_05281_ ), .A3(_05282_ ), .A4(_05283_ ), .ZN(_05284_ ) );
BUF_X4 _13038_ ( .A(_02093_ ), .Z(_05285_ ) );
XNOR2_X1 _13039_ ( .A(fanout_net_4 ), .B(\ID_EX_csr [1] ), .ZN(_05286_ ) );
INV_X1 _13040_ ( .A(_05286_ ), .ZN(_05287_ ) );
XOR2_X1 _13041_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .Z(_05288_ ) );
NOR4_X1 _13042_ ( .A1(_05284_ ), .A2(_05285_ ), .A3(_05287_ ), .A4(_05288_ ), .ZN(_05289_ ) );
AND2_X1 _13043_ ( .A1(_05279_ ), .A2(_05289_ ), .ZN(_05290_ ) );
BUF_X4 _13044_ ( .A(_05290_ ), .Z(_05291_ ) );
INV_X1 _13045_ ( .A(_05291_ ), .ZN(_05292_ ) );
BUF_X4 _13046_ ( .A(_05292_ ), .Z(_05293_ ) );
MUX2_X1 _13047_ ( .A(_05226_ ), .B(_05269_ ), .S(_05293_ ), .Z(_05294_ ) );
AOI211_X1 _13048_ ( .A(_03892_ ), .B(_05225_ ), .C1(\ID_EX_typ [3] ), .C2(_05294_ ), .ZN(_05295_ ) );
OAI21_X1 _13049_ ( .A(_03892_ ), .B1(_05222_ ), .B2(fanout_net_5 ), .ZN(_05296_ ) );
AOI21_X1 _13050_ ( .A(_05296_ ), .B1(_02995_ ), .B2(fanout_net_5 ), .ZN(_05297_ ) );
NOR2_X1 _13051_ ( .A1(_05295_ ), .A2(_05297_ ), .ZN(_05298_ ) );
INV_X2 _13052_ ( .A(_03886_ ), .ZN(_05299_ ) );
BUF_X4 _13053_ ( .A(_05299_ ), .Z(_05300_ ) );
NOR2_X1 _13054_ ( .A1(_05298_ ), .A2(_05300_ ), .ZN(_00122_ ) );
INV_X1 _13055_ ( .A(_05223_ ), .ZN(_05301_ ) );
BUF_X4 _13056_ ( .A(_05301_ ), .Z(_05302_ ) );
NAND4_X1 _13057_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_pc [16] ), .A3(\ID_EX_pc [15] ), .A4(\ID_EX_pc [14] ), .ZN(_05303_ ) );
NAND2_X1 _13058_ ( .A1(\ID_EX_pc [13] ), .A2(\ID_EX_pc [12] ), .ZN(_05304_ ) );
INV_X1 _13059_ ( .A(\ID_EX_pc [11] ), .ZN(_05305_ ) );
INV_X1 _13060_ ( .A(\ID_EX_pc [10] ), .ZN(_05306_ ) );
NOR4_X1 _13061_ ( .A1(_05303_ ), .A2(_05304_ ), .A3(_05305_ ), .A4(_05306_ ), .ZN(_05307_ ) );
AND2_X1 _13062_ ( .A1(_03899_ ), .A2(_05307_ ), .ZN(_05308_ ) );
AND4_X1 _13063_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_pc [23] ), .A4(\ID_EX_pc [22] ), .ZN(_05309_ ) );
AND2_X1 _13064_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_pc [18] ), .ZN(_05310_ ) );
AND4_X1 _13065_ ( .A1(\ID_EX_pc [21] ), .A2(_05309_ ), .A3(\ID_EX_pc [20] ), .A4(_05310_ ), .ZN(_05311_ ) );
AND2_X1 _13066_ ( .A1(_05308_ ), .A2(_05311_ ), .ZN(_05312_ ) );
NAND3_X1 _13067_ ( .A1(_05312_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_05313_ ) );
INV_X1 _13068_ ( .A(\ID_EX_pc [28] ), .ZN(_05314_ ) );
NOR2_X1 _13069_ ( .A1(_05313_ ), .A2(_05314_ ), .ZN(_05315_ ) );
XNOR2_X1 _13070_ ( .A(_05315_ ), .B(_05217_ ), .ZN(_05316_ ) );
NAND2_X1 _13071_ ( .A1(_05302_ ), .A2(_05316_ ), .ZN(_05317_ ) );
INV_X2 _13072_ ( .A(\ID_EX_typ [3] ), .ZN(_05318_ ) );
BUF_X4 _13073_ ( .A(_05318_ ), .Z(_05319_ ) );
BUF_X4 _13074_ ( .A(_05301_ ), .Z(_05320_ ) );
XNOR2_X1 _13075_ ( .A(\ID_EX_pc [29] ), .B(\ID_EX_imm [29] ), .ZN(_05321_ ) );
XNOR2_X1 _13076_ ( .A(_05216_ ), .B(_05321_ ), .ZN(_05322_ ) );
OAI211_X1 _13077_ ( .A(_05317_ ), .B(_05319_ ), .C1(_05320_ ), .C2(_05322_ ), .ZN(_05323_ ) );
INV_X2 _13078_ ( .A(_03876_ ), .ZN(_05324_ ) );
BUF_X4 _13079_ ( .A(_05324_ ), .Z(_05325_ ) );
BUF_X4 _13080_ ( .A(_05319_ ), .Z(_05326_ ) );
BUF_X4 _13081_ ( .A(_05234_ ), .Z(_05327_ ) );
BUF_X4 _13082_ ( .A(_05327_ ), .Z(_05328_ ) );
NAND3_X1 _13083_ ( .A1(_05328_ ), .A2(\mycsreg.CSReg[0][29] ), .A3(_05242_ ), .ZN(_05329_ ) );
BUF_X2 _13084_ ( .A(_05261_ ), .Z(_05330_ ) );
BUF_X2 _13085_ ( .A(_05330_ ), .Z(_05331_ ) );
NAND3_X1 _13086_ ( .A1(_05328_ ), .A2(\mtvec [29] ), .A3(_05331_ ), .ZN(_05332_ ) );
BUF_X2 _13087_ ( .A(_05230_ ), .Z(_05333_ ) );
BUF_X2 _13088_ ( .A(_05245_ ), .Z(_05334_ ) );
NAND4_X1 _13089_ ( .A1(_05333_ ), .A2(_05334_ ), .A3(_05253_ ), .A4(\mepc [29] ), .ZN(_05335_ ) );
BUF_X4 _13090_ ( .A(_05246_ ), .Z(_05336_ ) );
BUF_X4 _13091_ ( .A(_05336_ ), .Z(_05337_ ) );
BUF_X4 _13092_ ( .A(_05256_ ), .Z(_05338_ ) );
BUF_X4 _13093_ ( .A(_05338_ ), .Z(_05339_ ) );
NAND3_X1 _13094_ ( .A1(_05337_ ), .A2(\mycsreg.CSReg[3][29] ), .A3(_05339_ ), .ZN(_05340_ ) );
NAND4_X1 _13095_ ( .A1(_05329_ ), .A2(_05332_ ), .A3(_05335_ ), .A4(_05340_ ), .ZN(_05341_ ) );
NOR3_X1 _13096_ ( .A1(_05341_ ), .A2(_05291_ ), .A3(_05268_ ), .ZN(_05342_ ) );
NOR2_X1 _13097_ ( .A1(_05293_ ), .A2(\EX_LS_result_csreg_mem [29] ), .ZN(_05343_ ) );
NOR2_X1 _13098_ ( .A1(_05342_ ), .A2(_05343_ ), .ZN(_05344_ ) );
OAI211_X1 _13099_ ( .A(_05323_ ), .B(_05325_ ), .C1(_05326_ ), .C2(_05344_ ), .ZN(_05345_ ) );
MUX2_X1 _13100_ ( .A(_05322_ ), .B(_03032_ ), .S(fanout_net_5 ), .Z(_05346_ ) );
BUF_X2 _13101_ ( .A(_05324_ ), .Z(_05347_ ) );
OR2_X1 _13102_ ( .A1(_05346_ ), .A2(_05347_ ), .ZN(_05348_ ) );
AOI21_X1 _13103_ ( .A(_05300_ ), .B1(_05345_ ), .B2(_05348_ ), .ZN(_00123_ ) );
NAND3_X1 _13104_ ( .A1(_03899_ ), .A2(_05307_ ), .A3(_05310_ ), .ZN(_05349_ ) );
XNOR2_X1 _13105_ ( .A(_05349_ ), .B(\ID_EX_pc [20] ), .ZN(_05350_ ) );
AOI21_X1 _13106_ ( .A(\ID_EX_typ [3] ), .B1(_05302_ ), .B2(_05350_ ), .ZN(_05351_ ) );
AND2_X1 _13107_ ( .A1(_05168_ ), .A2(_05182_ ), .ZN(_05352_ ) );
OR2_X1 _13108_ ( .A1(_05352_ ), .A2(_05191_ ), .ZN(_05353_ ) );
XOR2_X1 _13109_ ( .A(_05353_ ), .B(_05173_ ), .Z(_05354_ ) );
INV_X1 _13110_ ( .A(_05354_ ), .ZN(_05355_ ) );
OAI21_X1 _13111_ ( .A(_05351_ ), .B1(_05320_ ), .B2(_05355_ ), .ZN(_05356_ ) );
AND3_X1 _13112_ ( .A1(_05234_ ), .A2(\mtvec [20] ), .A3(_05261_ ), .ZN(_05357_ ) );
AND2_X1 _13113_ ( .A1(_05267_ ), .A2(_05256_ ), .ZN(_05358_ ) );
BUF_X4 _13114_ ( .A(_05358_ ), .Z(_05359_ ) );
NOR3_X1 _13115_ ( .A1(_05357_ ), .A2(_05268_ ), .A3(_05359_ ), .ZN(_05360_ ) );
NAND3_X1 _13116_ ( .A1(_05234_ ), .A2(\mycsreg.CSReg[0][20] ), .A3(_05240_ ), .ZN(_05361_ ) );
NAND3_X1 _13117_ ( .A1(_05246_ ), .A2(\mepc [20] ), .A3(_05251_ ), .ZN(_05362_ ) );
NAND3_X1 _13118_ ( .A1(_05246_ ), .A2(\mycsreg.CSReg[3][20] ), .A3(_05338_ ), .ZN(_05363_ ) );
AND3_X1 _13119_ ( .A1(_05361_ ), .A2(_05362_ ), .A3(_05363_ ), .ZN(_05364_ ) );
AOI21_X1 _13120_ ( .A(_05291_ ), .B1(_05360_ ), .B2(_05364_ ), .ZN(_05365_ ) );
BUF_X2 _13121_ ( .A(_05279_ ), .Z(_05366_ ) );
BUF_X2 _13122_ ( .A(_05289_ ), .Z(_05367_ ) );
AND3_X1 _13123_ ( .A1(_05366_ ), .A2(_05367_ ), .A3(\EX_LS_result_csreg_mem [20] ), .ZN(_05368_ ) );
OR2_X1 _13124_ ( .A1(_05365_ ), .A2(_05368_ ), .ZN(_05369_ ) );
OAI211_X1 _13125_ ( .A(_05356_ ), .B(_05325_ ), .C1(_05326_ ), .C2(_05369_ ), .ZN(_05370_ ) );
AND2_X2 _13126_ ( .A1(_03876_ ), .A2(fanout_net_5 ), .ZN(_05371_ ) );
AND3_X1 _13127_ ( .A1(_03001_ ), .A2(_02998_ ), .A3(_05371_ ), .ZN(_05372_ ) );
BUF_X4 _13128_ ( .A(_03878_ ), .Z(_05373_ ) );
BUF_X4 _13129_ ( .A(_05373_ ), .Z(_05374_ ) );
AOI21_X1 _13130_ ( .A(_05372_ ), .B1(_05374_ ), .B2(_05354_ ), .ZN(_05375_ ) );
AOI21_X1 _13131_ ( .A(_05300_ ), .B1(_05370_ ), .B2(_05375_ ), .ZN(_00124_ ) );
BUF_X4 _13132_ ( .A(_05324_ ), .Z(_05376_ ) );
BUF_X4 _13133_ ( .A(_05318_ ), .Z(_05377_ ) );
BUF_X2 _13134_ ( .A(_05240_ ), .Z(_05378_ ) );
NAND3_X1 _13135_ ( .A1(_05327_ ), .A2(\mycsreg.CSReg[0][19] ), .A3(_05378_ ), .ZN(_05379_ ) );
NAND3_X1 _13136_ ( .A1(_05327_ ), .A2(\mtvec [19] ), .A3(_05262_ ), .ZN(_05380_ ) );
NAND3_X1 _13137_ ( .A1(_05336_ ), .A2(\mycsreg.CSReg[3][19] ), .A3(_05257_ ), .ZN(_05381_ ) );
AND3_X1 _13138_ ( .A1(_05379_ ), .A2(_05380_ ), .A3(_05381_ ), .ZN(_05382_ ) );
BUF_X2 _13139_ ( .A(_05251_ ), .Z(_05383_ ) );
AND3_X1 _13140_ ( .A1(_05336_ ), .A2(\mepc [19] ), .A3(_05383_ ), .ZN(_05384_ ) );
NOR2_X1 _13141_ ( .A1(_05384_ ), .A2(_05359_ ), .ZN(_05385_ ) );
BUF_X2 _13142_ ( .A(_05366_ ), .Z(_05386_ ) );
BUF_X2 _13143_ ( .A(_05367_ ), .Z(_05387_ ) );
AOI22_X1 _13144_ ( .A1(_05382_ ), .A2(_05385_ ), .B1(_05386_ ), .B2(_05387_ ), .ZN(_05388_ ) );
AND3_X1 _13145_ ( .A1(_05386_ ), .A2(_05387_ ), .A3(\EX_LS_result_csreg_mem [19] ), .ZN(_05389_ ) );
NOR2_X1 _13146_ ( .A1(_05388_ ), .A2(_05389_ ), .ZN(_05390_ ) );
INV_X1 _13147_ ( .A(_05390_ ), .ZN(_05391_ ) );
INV_X1 _13148_ ( .A(_05177_ ), .ZN(_05392_ ) );
NAND2_X1 _13149_ ( .A1(_05168_ ), .A2(_05181_ ), .ZN(_05393_ ) );
AOI21_X1 _13150_ ( .A(_05392_ ), .B1(_05393_ ), .B2(_05189_ ), .ZN(_05394_ ) );
OR2_X1 _13151_ ( .A1(_05394_ ), .A2(_05184_ ), .ZN(_05395_ ) );
XNOR2_X1 _13152_ ( .A(_05395_ ), .B(_05176_ ), .ZN(_05396_ ) );
OAI21_X1 _13153_ ( .A(_05377_ ), .B1(_05320_ ), .B2(_05396_ ), .ZN(_05397_ ) );
NAND3_X1 _13154_ ( .A1(_03899_ ), .A2(\ID_EX_pc [18] ), .A3(_05307_ ), .ZN(_05398_ ) );
INV_X1 _13155_ ( .A(\ID_EX_pc [19] ), .ZN(_05399_ ) );
XNOR2_X1 _13156_ ( .A(_05398_ ), .B(_05399_ ), .ZN(_05400_ ) );
AOI21_X1 _13157_ ( .A(_05400_ ), .B1(_05104_ ), .B2(_05106_ ), .ZN(_05401_ ) );
OAI221_X1 _13158_ ( .A(_05376_ ), .B1(_05377_ ), .B2(_05391_ ), .C1(_05397_ ), .C2(_05401_ ), .ZN(_05402_ ) );
INV_X1 _13159_ ( .A(_05371_ ), .ZN(_05403_ ) );
NOR2_X1 _13160_ ( .A1(_03010_ ), .A2(_05403_ ), .ZN(_05404_ ) );
NOR2_X1 _13161_ ( .A1(_05396_ ), .A2(_03879_ ), .ZN(_05405_ ) );
NOR2_X1 _13162_ ( .A1(_05404_ ), .A2(_05405_ ), .ZN(_05406_ ) );
AOI21_X1 _13163_ ( .A(_05300_ ), .B1(_05402_ ), .B2(_05406_ ), .ZN(_00125_ ) );
BUF_X4 _13164_ ( .A(_05324_ ), .Z(_05407_ ) );
BUF_X2 _13165_ ( .A(_05234_ ), .Z(_05408_ ) );
NAND3_X1 _13166_ ( .A1(_05408_ ), .A2(\mycsreg.CSReg[0][18] ), .A3(_05241_ ), .ZN(_05409_ ) );
NAND3_X1 _13167_ ( .A1(_05408_ ), .A2(\mtvec [18] ), .A3(_05330_ ), .ZN(_05410_ ) );
NAND3_X1 _13168_ ( .A1(_05336_ ), .A2(\mycsreg.CSReg[3][18] ), .A3(_05338_ ), .ZN(_05411_ ) );
AND3_X1 _13169_ ( .A1(_05409_ ), .A2(_05410_ ), .A3(_05411_ ), .ZN(_05412_ ) );
NAND3_X1 _13170_ ( .A1(_05336_ ), .A2(\mepc [18] ), .A3(_05252_ ), .ZN(_05413_ ) );
INV_X1 _13171_ ( .A(_05359_ ), .ZN(_05414_ ) );
AND2_X1 _13172_ ( .A1(_05413_ ), .A2(_05414_ ), .ZN(_05415_ ) );
AOI22_X1 _13173_ ( .A1(_05412_ ), .A2(_05415_ ), .B1(_05386_ ), .B2(_05387_ ), .ZN(_05416_ ) );
AND3_X1 _13174_ ( .A1(_05366_ ), .A2(_05367_ ), .A3(\EX_LS_result_csreg_mem [18] ), .ZN(_05417_ ) );
NOR2_X1 _13175_ ( .A1(_05416_ ), .A2(_05417_ ), .ZN(_05418_ ) );
INV_X1 _13176_ ( .A(_05418_ ), .ZN(_05419_ ) );
NAND2_X1 _13177_ ( .A1(_05393_ ), .A2(_05189_ ), .ZN(_05420_ ) );
XNOR2_X1 _13178_ ( .A(_05420_ ), .B(_05392_ ), .ZN(_05421_ ) );
INV_X1 _13179_ ( .A(_05421_ ), .ZN(_05422_ ) );
OAI21_X1 _13180_ ( .A(_05377_ ), .B1(_05320_ ), .B2(_05422_ ), .ZN(_05423_ ) );
XNOR2_X1 _13181_ ( .A(_05308_ ), .B(\ID_EX_pc [18] ), .ZN(_05424_ ) );
AOI21_X1 _13182_ ( .A(_05424_ ), .B1(_05104_ ), .B2(_05106_ ), .ZN(_05425_ ) );
OAI221_X1 _13183_ ( .A(_05407_ ), .B1(_05377_ ), .B2(_05419_ ), .C1(_05423_ ), .C2(_05425_ ), .ZN(_05426_ ) );
BUF_X4 _13184_ ( .A(_05371_ ), .Z(_05427_ ) );
AOI22_X1 _13185_ ( .A1(_03012_ ), .A2(_05427_ ), .B1(_05374_ ), .B2(_05421_ ), .ZN(_05428_ ) );
AOI21_X1 _13186_ ( .A(_05300_ ), .B1(_05426_ ), .B2(_05428_ ), .ZN(_00126_ ) );
AND2_X1 _13187_ ( .A1(_03903_ ), .A2(\ID_EX_pc [16] ), .ZN(_05429_ ) );
XNOR2_X1 _13188_ ( .A(_05429_ ), .B(\ID_EX_pc [17] ), .ZN(_05430_ ) );
AND2_X1 _13189_ ( .A1(_05168_ ), .A2(_05179_ ), .ZN(_05431_ ) );
OR2_X1 _13190_ ( .A1(_05431_ ), .A2(_05187_ ), .ZN(_05432_ ) );
XNOR2_X1 _13191_ ( .A(_05432_ ), .B(_05180_ ), .ZN(_05433_ ) );
MUX2_X1 _13192_ ( .A(_05430_ ), .B(_05433_ ), .S(_05224_ ), .Z(_05434_ ) );
NAND2_X1 _13193_ ( .A1(_05434_ ), .A2(_05377_ ), .ZN(_05435_ ) );
BUF_X4 _13194_ ( .A(_05324_ ), .Z(_05436_ ) );
NAND3_X1 _13195_ ( .A1(_05408_ ), .A2(\mtvec [17] ), .A3(_05330_ ), .ZN(_05437_ ) );
NAND3_X1 _13196_ ( .A1(_05336_ ), .A2(\mycsreg.CSReg[3][17] ), .A3(_05338_ ), .ZN(_05438_ ) );
AND2_X1 _13197_ ( .A1(_05437_ ), .A2(_05438_ ), .ZN(_05439_ ) );
NAND3_X1 _13198_ ( .A1(_05408_ ), .A2(\mycsreg.CSReg[0][17] ), .A3(_05241_ ), .ZN(_05440_ ) );
NAND3_X1 _13199_ ( .A1(_05336_ ), .A2(\mepc [17] ), .A3(_05252_ ), .ZN(_05441_ ) );
AND2_X1 _13200_ ( .A1(_05440_ ), .A2(_05441_ ), .ZN(_05442_ ) );
NOR2_X1 _13201_ ( .A1(_05268_ ), .A2(_05359_ ), .ZN(_05443_ ) );
BUF_X4 _13202_ ( .A(_05443_ ), .Z(_05444_ ) );
NAND4_X1 _13203_ ( .A1(_05293_ ), .A2(_05439_ ), .A3(_05442_ ), .A4(_05444_ ), .ZN(_05445_ ) );
INV_X1 _13204_ ( .A(\EX_LS_result_csreg_mem [17] ), .ZN(_05446_ ) );
NAND3_X1 _13205_ ( .A1(_05386_ ), .A2(_05387_ ), .A3(_05446_ ), .ZN(_05447_ ) );
AND2_X1 _13206_ ( .A1(_05445_ ), .A2(_05447_ ), .ZN(_05448_ ) );
OAI211_X1 _13207_ ( .A(_05435_ ), .B(_05436_ ), .C1(_05326_ ), .C2(_05448_ ), .ZN(_05449_ ) );
NOR2_X1 _13208_ ( .A1(_03014_ ), .A2(_05403_ ), .ZN(_05450_ ) );
NOR2_X1 _13209_ ( .A1(_05433_ ), .A2(_03879_ ), .ZN(_05451_ ) );
NOR2_X1 _13210_ ( .A1(_05450_ ), .A2(_05451_ ), .ZN(_05452_ ) );
AOI21_X1 _13211_ ( .A(_05300_ ), .B1(_05449_ ), .B2(_05452_ ), .ZN(_00127_ ) );
INV_X1 _13212_ ( .A(\ID_EX_pc [16] ), .ZN(_05453_ ) );
XNOR2_X1 _13213_ ( .A(_03903_ ), .B(_05453_ ), .ZN(_05454_ ) );
AOI21_X1 _13214_ ( .A(\ID_EX_typ [3] ), .B1(_05301_ ), .B2(_05454_ ), .ZN(_05455_ ) );
XOR2_X1 _13215_ ( .A(_05168_ ), .B(_05179_ ), .Z(_05456_ ) );
INV_X1 _13216_ ( .A(_05456_ ), .ZN(_05457_ ) );
OAI21_X1 _13217_ ( .A(_05455_ ), .B1(_05320_ ), .B2(_05457_ ), .ZN(_05458_ ) );
NAND3_X1 _13218_ ( .A1(_05327_ ), .A2(\mycsreg.CSReg[0][16] ), .A3(_05378_ ), .ZN(_05459_ ) );
NAND4_X1 _13219_ ( .A1(_05333_ ), .A2(_05334_ ), .A3(_05383_ ), .A4(\mepc [16] ), .ZN(_05460_ ) );
AND4_X1 _13220_ ( .A1(_02092_ ), .A2(_05270_ ), .A3(_05275_ ), .A4(_05282_ ), .ZN(_05461_ ) );
AND4_X1 _13221_ ( .A1(_05271_ ), .A2(_05286_ ), .A3(_05280_ ), .A4(_05281_ ), .ZN(_05462_ ) );
NAND2_X1 _13222_ ( .A1(_05461_ ), .A2(_05462_ ), .ZN(_05463_ ) );
AND3_X1 _13223_ ( .A1(_05277_ ), .A2(_05278_ ), .A3(_05283_ ), .ZN(_05464_ ) );
XNOR2_X1 _13224_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .ZN(_05465_ ) );
NAND3_X1 _13225_ ( .A1(_05464_ ), .A2(_05272_ ), .A3(_05465_ ), .ZN(_05466_ ) );
OAI211_X1 _13226_ ( .A(_05459_ ), .B(_05460_ ), .C1(_05463_ ), .C2(_05466_ ), .ZN(_05467_ ) );
NAND3_X1 _13227_ ( .A1(_05327_ ), .A2(\mtvec [16] ), .A3(_05262_ ), .ZN(_05468_ ) );
BUF_X2 _13228_ ( .A(_05246_ ), .Z(_05469_ ) );
NAND3_X1 _13229_ ( .A1(_05469_ ), .A2(\mycsreg.CSReg[3][16] ), .A3(_05257_ ), .ZN(_05470_ ) );
NAND3_X1 _13230_ ( .A1(_05443_ ), .A2(_05468_ ), .A3(_05470_ ), .ZN(_05471_ ) );
NOR2_X1 _13231_ ( .A1(_05467_ ), .A2(_05471_ ), .ZN(_05472_ ) );
BUF_X2 _13232_ ( .A(_05463_ ), .Z(_05473_ ) );
CLKBUF_X2 _13233_ ( .A(_05466_ ), .Z(_05474_ ) );
NOR3_X1 _13234_ ( .A1(_05473_ ), .A2(_05474_ ), .A3(\EX_LS_result_csreg_mem [16] ), .ZN(_05475_ ) );
NOR2_X1 _13235_ ( .A1(_05472_ ), .A2(_05475_ ), .ZN(_05476_ ) );
OAI211_X1 _13236_ ( .A(_05458_ ), .B(_05436_ ), .C1(_05326_ ), .C2(_05476_ ), .ZN(_05477_ ) );
NOR3_X1 _13237_ ( .A1(_03015_ ), .A2(_03005_ ), .A3(_05403_ ), .ZN(_05478_ ) );
AOI21_X1 _13238_ ( .A(_05478_ ), .B1(_05374_ ), .B2(_05456_ ), .ZN(_05479_ ) );
AOI21_X1 _13239_ ( .A(_05300_ ), .B1(_05477_ ), .B2(_05479_ ), .ZN(_00128_ ) );
BUF_X4 _13240_ ( .A(_05224_ ), .Z(_05480_ ) );
INV_X1 _13241_ ( .A(_05154_ ), .ZN(_05481_ ) );
OAI21_X1 _13242_ ( .A(_05157_ ), .B1(_05143_ ), .B2(_05151_ ), .ZN(_05482_ ) );
AOI21_X1 _13243_ ( .A(_05481_ ), .B1(_05482_ ), .B2(_05161_ ), .ZN(_05483_ ) );
NOR2_X1 _13244_ ( .A1(_05483_ ), .A2(_05165_ ), .ZN(_05484_ ) );
XNOR2_X1 _13245_ ( .A(_05484_ ), .B(_05153_ ), .ZN(_05485_ ) );
AOI21_X1 _13246_ ( .A(\ID_EX_typ [3] ), .B1(_05480_ ), .B2(_05485_ ), .ZN(_05486_ ) );
AND2_X1 _13247_ ( .A1(_03902_ ), .A2(\ID_EX_pc [14] ), .ZN(_05487_ ) );
XNOR2_X1 _13248_ ( .A(_05487_ ), .B(\ID_EX_pc [15] ), .ZN(_05488_ ) );
OAI21_X1 _13249_ ( .A(_05486_ ), .B1(_05480_ ), .B2(_05488_ ), .ZN(_05489_ ) );
NAND3_X1 _13250_ ( .A1(_05260_ ), .A2(\mycsreg.CSReg[0][15] ), .A3(_05378_ ), .ZN(_05490_ ) );
NAND3_X1 _13251_ ( .A1(_05260_ ), .A2(\mtvec [15] ), .A3(_05262_ ), .ZN(_05491_ ) );
NAND3_X1 _13252_ ( .A1(_05469_ ), .A2(\mycsreg.CSReg[3][15] ), .A3(_05257_ ), .ZN(_05492_ ) );
AND3_X1 _13253_ ( .A1(_05490_ ), .A2(_05491_ ), .A3(_05492_ ), .ZN(_05493_ ) );
AND3_X1 _13254_ ( .A1(_05469_ ), .A2(\mepc [15] ), .A3(_05383_ ), .ZN(_05494_ ) );
NOR2_X1 _13255_ ( .A1(_05494_ ), .A2(_05359_ ), .ZN(_05495_ ) );
CLKBUF_X2 _13256_ ( .A(_05366_ ), .Z(_05496_ ) );
CLKBUF_X2 _13257_ ( .A(_05367_ ), .Z(_05497_ ) );
AOI22_X1 _13258_ ( .A1(_05493_ ), .A2(_05495_ ), .B1(_05496_ ), .B2(_05497_ ), .ZN(_05498_ ) );
AND3_X1 _13259_ ( .A1(_05386_ ), .A2(_05387_ ), .A3(\EX_LS_result_csreg_mem [15] ), .ZN(_05499_ ) );
NOR2_X1 _13260_ ( .A1(_05498_ ), .A2(_05499_ ), .ZN(_05500_ ) );
INV_X1 _13261_ ( .A(_05500_ ), .ZN(_05501_ ) );
OAI211_X1 _13262_ ( .A(_05489_ ), .B(_05436_ ), .C1(_05326_ ), .C2(_05501_ ), .ZN(_05502_ ) );
NOR2_X1 _13263_ ( .A1(_03025_ ), .A2(_05403_ ), .ZN(_05503_ ) );
AOI21_X1 _13264_ ( .A(_05503_ ), .B1(_05374_ ), .B2(_05485_ ), .ZN(_05504_ ) );
AOI21_X1 _13265_ ( .A(_05300_ ), .B1(_05502_ ), .B2(_05504_ ), .ZN(_00129_ ) );
INV_X1 _13266_ ( .A(\ID_EX_pc [14] ), .ZN(_05505_ ) );
XNOR2_X1 _13267_ ( .A(_03902_ ), .B(_05505_ ), .ZN(_05506_ ) );
AND3_X1 _13268_ ( .A1(_05482_ ), .A2(_05481_ ), .A3(_05161_ ), .ZN(_05507_ ) );
NOR2_X1 _13269_ ( .A1(_05507_ ), .A2(_05483_ ), .ZN(_05508_ ) );
MUX2_X1 _13270_ ( .A(_05506_ ), .B(_05508_ ), .S(_05224_ ), .Z(_05509_ ) );
OR2_X1 _13271_ ( .A1(_05509_ ), .A2(\ID_EX_typ [3] ), .ZN(_05510_ ) );
NAND3_X1 _13272_ ( .A1(_05327_ ), .A2(\mycsreg.CSReg[0][14] ), .A3(_05378_ ), .ZN(_05511_ ) );
NAND4_X1 _13273_ ( .A1(_05333_ ), .A2(_05334_ ), .A3(_05383_ ), .A4(\mepc [14] ), .ZN(_05512_ ) );
OAI211_X1 _13274_ ( .A(_05511_ ), .B(_05512_ ), .C1(_05463_ ), .C2(_05466_ ), .ZN(_05513_ ) );
NAND3_X1 _13275_ ( .A1(_05327_ ), .A2(\mtvec [14] ), .A3(_05262_ ), .ZN(_05514_ ) );
NAND3_X1 _13276_ ( .A1(_05469_ ), .A2(\mycsreg.CSReg[3][14] ), .A3(_05257_ ), .ZN(_05515_ ) );
NAND3_X1 _13277_ ( .A1(_05443_ ), .A2(_05514_ ), .A3(_05515_ ), .ZN(_05516_ ) );
NOR2_X1 _13278_ ( .A1(_05513_ ), .A2(_05516_ ), .ZN(_05517_ ) );
NOR3_X1 _13279_ ( .A1(_05473_ ), .A2(_05474_ ), .A3(\EX_LS_result_csreg_mem [14] ), .ZN(_05518_ ) );
NOR2_X1 _13280_ ( .A1(_05517_ ), .A2(_05518_ ), .ZN(_05519_ ) );
OAI211_X1 _13281_ ( .A(_05510_ ), .B(_05436_ ), .C1(_05326_ ), .C2(_05519_ ), .ZN(_05520_ ) );
AOI22_X1 _13282_ ( .A1(_03026_ ), .A2(_05427_ ), .B1(_05374_ ), .B2(_05508_ ), .ZN(_05521_ ) );
AOI21_X1 _13283_ ( .A(_05300_ ), .B1(_05520_ ), .B2(_05521_ ), .ZN(_00130_ ) );
BUF_X4 _13284_ ( .A(_05299_ ), .Z(_05522_ ) );
AND2_X1 _13285_ ( .A1(_05152_ ), .A2(_05155_ ), .ZN(_05523_ ) );
NOR2_X1 _13286_ ( .A1(_05523_ ), .A2(_05159_ ), .ZN(_05524_ ) );
XNOR2_X1 _13287_ ( .A(_05524_ ), .B(_05156_ ), .ZN(_05525_ ) );
AOI21_X1 _13288_ ( .A(\ID_EX_typ [3] ), .B1(_05480_ ), .B2(_05525_ ), .ZN(_05526_ ) );
AND2_X1 _13289_ ( .A1(_03901_ ), .A2(\ID_EX_pc [12] ), .ZN(_05527_ ) );
XNOR2_X1 _13290_ ( .A(_05527_ ), .B(\ID_EX_pc [13] ), .ZN(_05528_ ) );
OAI21_X1 _13291_ ( .A(_05526_ ), .B1(_05480_ ), .B2(_05528_ ), .ZN(_05529_ ) );
NOR2_X1 _13292_ ( .A1(_05463_ ), .A2(_05466_ ), .ZN(_05530_ ) );
INV_X1 _13293_ ( .A(_05530_ ), .ZN(_05531_ ) );
NAND3_X1 _13294_ ( .A1(_05234_ ), .A2(\mycsreg.CSReg[0][13] ), .A3(_05240_ ), .ZN(_05532_ ) );
NAND4_X1 _13295_ ( .A1(_05333_ ), .A2(_05334_ ), .A3(_05251_ ), .A4(\mepc [13] ), .ZN(_05533_ ) );
AND2_X1 _13296_ ( .A1(_05532_ ), .A2(_05533_ ), .ZN(_05534_ ) );
AND3_X1 _13297_ ( .A1(_05234_ ), .A2(\mtvec [13] ), .A3(_05261_ ), .ZN(_05535_ ) );
INV_X1 _13298_ ( .A(_05535_ ), .ZN(_05536_ ) );
AND3_X1 _13299_ ( .A1(_05246_ ), .A2(\mycsreg.CSReg[3][13] ), .A3(_05256_ ), .ZN(_05537_ ) );
NOR2_X1 _13300_ ( .A1(_05537_ ), .A2(_05268_ ), .ZN(_05538_ ) );
NAND4_X1 _13301_ ( .A1(_05531_ ), .A2(_05534_ ), .A3(_05536_ ), .A4(_05538_ ), .ZN(_05539_ ) );
NOR3_X1 _13302_ ( .A1(_05463_ ), .A2(_05466_ ), .A3(\EX_LS_result_csreg_mem [13] ), .ZN(_05540_ ) );
INV_X1 _13303_ ( .A(_05540_ ), .ZN(_05541_ ) );
AND2_X1 _13304_ ( .A1(_05539_ ), .A2(_05541_ ), .ZN(_05542_ ) );
OAI211_X1 _13305_ ( .A(_05529_ ), .B(_05436_ ), .C1(_05326_ ), .C2(_05542_ ), .ZN(_05543_ ) );
NOR2_X1 _13306_ ( .A1(_03029_ ), .A2(_05403_ ), .ZN(_05544_ ) );
AOI21_X1 _13307_ ( .A(_05544_ ), .B1(_05374_ ), .B2(_05525_ ), .ZN(_05545_ ) );
AOI21_X1 _13308_ ( .A(_05522_ ), .B1(_05543_ ), .B2(_05545_ ), .ZN(_00131_ ) );
INV_X1 _13309_ ( .A(\ID_EX_pc [12] ), .ZN(_05546_ ) );
XNOR2_X1 _13310_ ( .A(_03901_ ), .B(_05546_ ), .ZN(_05547_ ) );
XOR2_X1 _13311_ ( .A(_05152_ ), .B(_05155_ ), .Z(_05548_ ) );
MUX2_X1 _13312_ ( .A(_05547_ ), .B(_05548_ ), .S(_05224_ ), .Z(_05549_ ) );
OR2_X1 _13313_ ( .A1(_05549_ ), .A2(\ID_EX_typ [3] ), .ZN(_05550_ ) );
NAND3_X1 _13314_ ( .A1(_05235_ ), .A2(\mycsreg.CSReg[0][12] ), .A3(_05241_ ), .ZN(_05551_ ) );
NAND4_X1 _13315_ ( .A1(_05333_ ), .A2(_05334_ ), .A3(_05252_ ), .A4(\mepc [12] ), .ZN(_05552_ ) );
AND2_X1 _13316_ ( .A1(_05551_ ), .A2(_05552_ ), .ZN(_05553_ ) );
NAND3_X1 _13317_ ( .A1(_05235_ ), .A2(\mtvec [12] ), .A3(_05330_ ), .ZN(_05554_ ) );
NAND3_X1 _13318_ ( .A1(_05247_ ), .A2(\mycsreg.CSReg[3][12] ), .A3(_05338_ ), .ZN(_05555_ ) );
AND2_X1 _13319_ ( .A1(_05554_ ), .A2(_05555_ ), .ZN(_05556_ ) );
NAND4_X1 _13320_ ( .A1(_05292_ ), .A2(_05553_ ), .A3(_05556_ ), .A4(_05443_ ), .ZN(_05557_ ) );
INV_X1 _13321_ ( .A(\EX_LS_result_csreg_mem [12] ), .ZN(_05558_ ) );
NAND3_X1 _13322_ ( .A1(_05366_ ), .A2(_05387_ ), .A3(_05558_ ), .ZN(_05559_ ) );
AND2_X1 _13323_ ( .A1(_05557_ ), .A2(_05559_ ), .ZN(_05560_ ) );
OAI211_X1 _13324_ ( .A(_05550_ ), .B(_05436_ ), .C1(_05326_ ), .C2(_05560_ ), .ZN(_05561_ ) );
AND3_X1 _13325_ ( .A1(_03030_ ), .A2(_03027_ ), .A3(_05371_ ), .ZN(_05562_ ) );
AOI21_X1 _13326_ ( .A(_05562_ ), .B1(_05374_ ), .B2(_05548_ ), .ZN(_05563_ ) );
AOI21_X1 _13327_ ( .A(_05522_ ), .B1(_05561_ ), .B2(_05563_ ), .ZN(_00132_ ) );
INV_X1 _13328_ ( .A(_05138_ ), .ZN(_05564_ ) );
NAND2_X1 _13329_ ( .A1(_05136_ ), .A2(_05142_ ), .ZN(_05565_ ) );
AOI21_X1 _13330_ ( .A(_05564_ ), .B1(_05565_ ), .B2(_05149_ ), .ZN(_05566_ ) );
NOR2_X1 _13331_ ( .A1(_05566_ ), .A2(_05144_ ), .ZN(_05567_ ) );
XNOR2_X1 _13332_ ( .A(_05567_ ), .B(_05137_ ), .ZN(_05568_ ) );
AOI21_X1 _13333_ ( .A(\ID_EX_typ [3] ), .B1(_05480_ ), .B2(_05568_ ), .ZN(_05569_ ) );
XNOR2_X1 _13334_ ( .A(_03900_ ), .B(\ID_EX_pc [11] ), .ZN(_05570_ ) );
OAI21_X1 _13335_ ( .A(_05569_ ), .B1(_05480_ ), .B2(_05570_ ), .ZN(_05571_ ) );
INV_X1 _13336_ ( .A(_05443_ ), .ZN(_05572_ ) );
NOR2_X1 _13337_ ( .A1(_05291_ ), .A2(_05572_ ), .ZN(_05573_ ) );
NAND3_X1 _13338_ ( .A1(_05469_ ), .A2(\mycsreg.CSReg[3][11] ), .A3(_05257_ ), .ZN(_05574_ ) );
NAND3_X1 _13339_ ( .A1(_05260_ ), .A2(\mtvec [11] ), .A3(_05262_ ), .ZN(_05575_ ) );
NAND3_X1 _13340_ ( .A1(_05260_ ), .A2(\mycsreg.CSReg[0][11] ), .A3(_05378_ ), .ZN(_05576_ ) );
NAND3_X1 _13341_ ( .A1(_05469_ ), .A2(\mepc [11] ), .A3(_05383_ ), .ZN(_05577_ ) );
AND4_X1 _13342_ ( .A1(_05574_ ), .A2(_05575_ ), .A3(_05576_ ), .A4(_05577_ ), .ZN(_05578_ ) );
AND2_X1 _13343_ ( .A1(_05573_ ), .A2(_05578_ ), .ZN(_05579_ ) );
INV_X1 _13344_ ( .A(\EX_LS_result_csreg_mem [11] ), .ZN(_05580_ ) );
AND3_X1 _13345_ ( .A1(_05496_ ), .A2(_05497_ ), .A3(_05580_ ), .ZN(_05581_ ) );
NOR2_X1 _13346_ ( .A1(_05579_ ), .A2(_05581_ ), .ZN(_05582_ ) );
OAI211_X1 _13347_ ( .A(_05571_ ), .B(_05436_ ), .C1(_05326_ ), .C2(_05582_ ), .ZN(_05583_ ) );
AOI21_X1 _13348_ ( .A(_02822_ ), .B1(_02626_ ), .B2(_02815_ ), .ZN(_05584_ ) );
AND3_X1 _13349_ ( .A1(_02721_ ), .A2(_02743_ ), .A3(_02740_ ), .ZN(_05585_ ) );
NOR3_X1 _13350_ ( .A1(_05584_ ), .A2(_02825_ ), .A3(_05585_ ), .ZN(_05586_ ) );
NOR2_X1 _13351_ ( .A1(_05586_ ), .A2(_02825_ ), .ZN(_05587_ ) );
XNOR2_X1 _13352_ ( .A(_05587_ ), .B(_02767_ ), .ZN(_05588_ ) );
AOI22_X1 _13353_ ( .A1(_05588_ ), .A2(_05427_ ), .B1(_05374_ ), .B2(_05568_ ), .ZN(_05589_ ) );
AOI21_X1 _13354_ ( .A(_05522_ ), .B1(_05583_ ), .B2(_05589_ ), .ZN(_00133_ ) );
XNOR2_X1 _13355_ ( .A(_05313_ ), .B(\ID_EX_pc [28] ), .ZN(_05590_ ) );
AND2_X1 _13356_ ( .A1(_05301_ ), .A2(_05590_ ), .ZN(_05591_ ) );
XOR2_X1 _13357_ ( .A(\ID_EX_pc [28] ), .B(\ID_EX_imm [28] ), .Z(_05592_ ) );
XNOR2_X1 _13358_ ( .A(_05212_ ), .B(_05592_ ), .ZN(_05593_ ) );
AOI211_X1 _13359_ ( .A(\ID_EX_typ [3] ), .B(_05591_ ), .C1(_05224_ ), .C2(_05593_ ), .ZN(_05594_ ) );
NAND3_X1 _13360_ ( .A1(_05327_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_05378_ ), .ZN(_05595_ ) );
NAND4_X1 _13361_ ( .A1(_05333_ ), .A2(_05334_ ), .A3(_05383_ ), .A4(\mepc [28] ), .ZN(_05596_ ) );
AND2_X1 _13362_ ( .A1(_05595_ ), .A2(_05596_ ), .ZN(_05597_ ) );
AND3_X1 _13363_ ( .A1(_05336_ ), .A2(\mycsreg.CSReg[3][28] ), .A3(_05257_ ), .ZN(_05598_ ) );
NOR2_X1 _13364_ ( .A1(_05598_ ), .A2(_05268_ ), .ZN(_05599_ ) );
AND3_X1 _13365_ ( .A1(_05408_ ), .A2(\mtvec [28] ), .A3(_05262_ ), .ZN(_05600_ ) );
INV_X1 _13366_ ( .A(_05600_ ), .ZN(_05601_ ) );
NAND4_X1 _13367_ ( .A1(_05597_ ), .A2(_05599_ ), .A3(_05531_ ), .A4(_05601_ ), .ZN(_05602_ ) );
CLKBUF_X2 _13368_ ( .A(_05466_ ), .Z(_05603_ ) );
OR3_X1 _13369_ ( .A1(_05473_ ), .A2(\EX_LS_result_csreg_mem [28] ), .A3(_05603_ ), .ZN(_05604_ ) );
NAND2_X1 _13370_ ( .A1(_05602_ ), .A2(_05604_ ), .ZN(_05605_ ) );
AOI21_X1 _13371_ ( .A(_05594_ ), .B1(\ID_EX_typ [3] ), .B2(_05605_ ), .ZN(_05606_ ) );
NAND2_X1 _13372_ ( .A1(_05606_ ), .A2(_05325_ ), .ZN(_05607_ ) );
OAI21_X1 _13373_ ( .A(fanout_net_5 ), .B1(_03033_ ), .B2(_02913_ ), .ZN(_05608_ ) );
CLKBUF_X2 _13374_ ( .A(_03876_ ), .Z(_05609_ ) );
BUF_X4 _13375_ ( .A(_05609_ ), .Z(_05610_ ) );
OAI211_X1 _13376_ ( .A(_05608_ ), .B(_05610_ ), .C1(fanout_net_5 ), .C2(_05593_ ), .ZN(_05611_ ) );
AOI21_X1 _13377_ ( .A(_05522_ ), .B1(_05607_ ), .B2(_05611_ ), .ZN(_00134_ ) );
AND3_X1 _13378_ ( .A1(_05408_ ), .A2(\mtvec [10] ), .A3(_05330_ ), .ZN(_05612_ ) );
NOR2_X1 _13379_ ( .A1(_05612_ ), .A2(_05359_ ), .ZN(_05613_ ) );
NAND3_X1 _13380_ ( .A1(_05235_ ), .A2(\mycsreg.CSReg[0][10] ), .A3(_05241_ ), .ZN(_05614_ ) );
NAND3_X1 _13381_ ( .A1(_05247_ ), .A2(\mepc [10] ), .A3(_05252_ ), .ZN(_05615_ ) );
NAND3_X1 _13382_ ( .A1(_05247_ ), .A2(\mycsreg.CSReg[3][10] ), .A3(_05338_ ), .ZN(_05616_ ) );
AND3_X1 _13383_ ( .A1(_05614_ ), .A2(_05615_ ), .A3(_05616_ ), .ZN(_05617_ ) );
AOI21_X1 _13384_ ( .A(_05291_ ), .B1(_05613_ ), .B2(_05617_ ), .ZN(_05618_ ) );
AND3_X1 _13385_ ( .A1(_05366_ ), .A2(_05367_ ), .A3(\EX_LS_result_csreg_mem [10] ), .ZN(_05619_ ) );
NOR2_X1 _13386_ ( .A1(_05618_ ), .A2(_05619_ ), .ZN(_05620_ ) );
INV_X1 _13387_ ( .A(_05620_ ), .ZN(_05621_ ) );
XNOR2_X1 _13388_ ( .A(_03899_ ), .B(_05306_ ), .ZN(_05622_ ) );
AND3_X1 _13389_ ( .A1(_05565_ ), .A2(_05564_ ), .A3(_05149_ ), .ZN(_05623_ ) );
NOR2_X1 _13390_ ( .A1(_05623_ ), .A2(_05566_ ), .ZN(_05624_ ) );
MUX2_X1 _13391_ ( .A(_05622_ ), .B(_05624_ ), .S(_05223_ ), .Z(_05625_ ) );
MUX2_X1 _13392_ ( .A(_05621_ ), .B(_05625_ ), .S(_05318_ ), .Z(_05626_ ) );
NAND2_X1 _13393_ ( .A1(_05626_ ), .A2(_05325_ ), .ZN(_05627_ ) );
XNOR2_X1 _13394_ ( .A(_05584_ ), .B(_02744_ ), .ZN(_05628_ ) );
AOI22_X1 _13395_ ( .A1(_05628_ ), .A2(_05427_ ), .B1(_05373_ ), .B2(_05624_ ), .ZN(_05629_ ) );
AOI21_X1 _13396_ ( .A(_05522_ ), .B1(_05627_ ), .B2(_05629_ ), .ZN(_00135_ ) );
INV_X1 _13397_ ( .A(\ID_EX_pc [9] ), .ZN(_05630_ ) );
XNOR2_X1 _13398_ ( .A(_03898_ ), .B(_05630_ ), .ZN(_05631_ ) );
AND2_X1 _13399_ ( .A1(_05136_ ), .A2(_05140_ ), .ZN(_05632_ ) );
NOR2_X1 _13400_ ( .A1(_05632_ ), .A2(_05147_ ), .ZN(_05633_ ) );
XNOR2_X1 _13401_ ( .A(_05633_ ), .B(_05141_ ), .ZN(_05634_ ) );
MUX2_X1 _13402_ ( .A(_05631_ ), .B(_05634_ ), .S(_05224_ ), .Z(_05635_ ) );
OR2_X1 _13403_ ( .A1(_05635_ ), .A2(\ID_EX_typ [3] ), .ZN(_05636_ ) );
AND3_X1 _13404_ ( .A1(_05496_ ), .A2(_05497_ ), .A3(\EX_LS_result_csreg_mem [9] ), .ZN(_05637_ ) );
INV_X1 _13405_ ( .A(_05637_ ), .ZN(_05638_ ) );
AND3_X1 _13406_ ( .A1(_05236_ ), .A2(\mtvec [9] ), .A3(_05331_ ), .ZN(_05639_ ) );
NOR2_X1 _13407_ ( .A1(_05639_ ), .A2(_05359_ ), .ZN(_05640_ ) );
NAND3_X1 _13408_ ( .A1(_05337_ ), .A2(\mepc [9] ), .A3(_05253_ ), .ZN(_05641_ ) );
NAND3_X1 _13409_ ( .A1(_05248_ ), .A2(\mycsreg.CSReg[3][9] ), .A3(_05339_ ), .ZN(_05642_ ) );
AND3_X1 _13410_ ( .A1(_05260_ ), .A2(\mycsreg.CSReg[0][9] ), .A3(_05378_ ), .ZN(_05643_ ) );
INV_X1 _13411_ ( .A(_05643_ ), .ZN(_05644_ ) );
AND4_X1 _13412_ ( .A1(_05640_ ), .A2(_05641_ ), .A3(_05642_ ), .A4(_05644_ ), .ZN(_05645_ ) );
OAI21_X1 _13413_ ( .A(_05638_ ), .B1(_05645_ ), .B2(_05291_ ), .ZN(_05646_ ) );
OAI211_X1 _13414_ ( .A(_05636_ ), .B(_05436_ ), .C1(_05326_ ), .C2(_05646_ ), .ZN(_05647_ ) );
AND2_X1 _13415_ ( .A1(_02626_ ), .A2(_02791_ ), .ZN(_05648_ ) );
OR2_X1 _13416_ ( .A1(_05648_ ), .A2(_02819_ ), .ZN(_05649_ ) );
XNOR2_X1 _13417_ ( .A(_05649_ ), .B(_02814_ ), .ZN(_05650_ ) );
NOR2_X1 _13418_ ( .A1(_05650_ ), .A2(_05403_ ), .ZN(_05651_ ) );
AOI21_X1 _13419_ ( .A(_05651_ ), .B1(_05374_ ), .B2(_05634_ ), .ZN(_05652_ ) );
AOI21_X1 _13420_ ( .A(_05522_ ), .B1(_05647_ ), .B2(_05652_ ), .ZN(_00136_ ) );
INV_X1 _13421_ ( .A(\EX_LS_result_csreg_mem [8] ), .ZN(_05653_ ) );
AND3_X1 _13422_ ( .A1(_05496_ ), .A2(_05497_ ), .A3(_05653_ ), .ZN(_05654_ ) );
NAND3_X1 _13423_ ( .A1(_05327_ ), .A2(\mycsreg.CSReg[0][8] ), .A3(_05378_ ), .ZN(_05655_ ) );
NAND3_X1 _13424_ ( .A1(_05260_ ), .A2(\mtvec [8] ), .A3(_05262_ ), .ZN(_05656_ ) );
NAND4_X1 _13425_ ( .A1(_05333_ ), .A2(_05334_ ), .A3(_05383_ ), .A4(\mepc [8] ), .ZN(_05657_ ) );
NAND3_X1 _13426_ ( .A1(_05469_ ), .A2(\mycsreg.CSReg[3][8] ), .A3(_05257_ ), .ZN(_05658_ ) );
AND4_X1 _13427_ ( .A1(_05655_ ), .A2(_05656_ ), .A3(_05657_ ), .A4(_05658_ ), .ZN(_05659_ ) );
AOI21_X1 _13428_ ( .A(_05654_ ), .B1(_05573_ ), .B2(_05659_ ), .ZN(_05660_ ) );
XNOR2_X1 _13429_ ( .A(_03897_ ), .B(\ID_EX_pc [8] ), .ZN(_05661_ ) );
OAI21_X1 _13430_ ( .A(_05377_ ), .B1(_05480_ ), .B2(_05661_ ), .ZN(_05662_ ) );
XOR2_X1 _13431_ ( .A(_05136_ ), .B(_05140_ ), .Z(_05663_ ) );
AND3_X1 _13432_ ( .A1(_05104_ ), .A2(_05106_ ), .A3(_05663_ ), .ZN(_05664_ ) );
OAI221_X1 _13433_ ( .A(_05407_ ), .B1(_05377_ ), .B2(_05660_ ), .C1(_05662_ ), .C2(_05664_ ), .ZN(_05665_ ) );
XNOR2_X1 _13434_ ( .A(_02625_ ), .B(_02791_ ), .ZN(_05666_ ) );
AOI22_X1 _13435_ ( .A1(_05666_ ), .A2(_05427_ ), .B1(_05373_ ), .B2(_05663_ ), .ZN(_05667_ ) );
AOI21_X1 _13436_ ( .A(_05522_ ), .B1(_05665_ ), .B2(_05667_ ), .ZN(_00137_ ) );
AND3_X1 _13437_ ( .A1(_05366_ ), .A2(_05367_ ), .A3(\EX_LS_result_csreg_mem [7] ), .ZN(_05668_ ) );
INV_X1 _13438_ ( .A(_05668_ ), .ZN(_05669_ ) );
NAND3_X1 _13439_ ( .A1(_05248_ ), .A2(\mycsreg.CSReg[3][7] ), .A3(_05339_ ), .ZN(_05670_ ) );
NAND3_X1 _13440_ ( .A1(_05236_ ), .A2(\mtvec [7] ), .A3(_05331_ ), .ZN(_05671_ ) );
NAND3_X1 _13441_ ( .A1(_05236_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_05242_ ), .ZN(_05672_ ) );
NAND3_X1 _13442_ ( .A1(_05248_ ), .A2(\mepc [7] ), .A3(_05253_ ), .ZN(_05673_ ) );
AND4_X1 _13443_ ( .A1(_05670_ ), .A2(_05671_ ), .A3(_05672_ ), .A4(_05673_ ), .ZN(_05674_ ) );
OAI21_X1 _13444_ ( .A(_05669_ ), .B1(_05674_ ), .B2(_05291_ ), .ZN(_05675_ ) );
INV_X1 _13445_ ( .A(\ID_EX_pc [7] ), .ZN(_05676_ ) );
XNOR2_X1 _13446_ ( .A(_03896_ ), .B(_05676_ ), .ZN(_05677_ ) );
XNOR2_X1 _13447_ ( .A(\ID_EX_pc [7] ), .B(\ID_EX_imm [7] ), .ZN(_05678_ ) );
XNOR2_X1 _13448_ ( .A(_05132_ ), .B(_05678_ ), .ZN(_05679_ ) );
MUX2_X1 _13449_ ( .A(_05677_ ), .B(_05679_ ), .S(_05223_ ), .Z(_05680_ ) );
MUX2_X1 _13450_ ( .A(_05675_ ), .B(_05680_ ), .S(_05318_ ), .Z(_05681_ ) );
NAND2_X1 _13451_ ( .A1(_05681_ ), .A2(_05325_ ), .ZN(_05682_ ) );
AOI21_X1 _13452_ ( .A(_02614_ ), .B1(_02519_ ), .B2(_02521_ ), .ZN(_05683_ ) );
NAND2_X1 _13453_ ( .A1(_05683_ ), .A2(_02620_ ), .ZN(_05684_ ) );
NAND2_X1 _13454_ ( .A1(_05684_ ), .A2(_02622_ ), .ZN(_05685_ ) );
NAND2_X1 _13455_ ( .A1(_05685_ ), .A2(_02566_ ), .ZN(_05686_ ) );
NAND2_X1 _13456_ ( .A1(_05686_ ), .A2(_02617_ ), .ZN(_05687_ ) );
XNOR2_X1 _13457_ ( .A(_05687_ ), .B(_02544_ ), .ZN(_05688_ ) );
AOI22_X1 _13458_ ( .A1(_05688_ ), .A2(_05427_ ), .B1(_05373_ ), .B2(_05679_ ), .ZN(_05689_ ) );
AOI21_X1 _13459_ ( .A(_05522_ ), .B1(_05682_ ), .B2(_05689_ ), .ZN(_00138_ ) );
XOR2_X1 _13460_ ( .A(_05128_ ), .B(_05129_ ), .Z(_05690_ ) );
AOI21_X1 _13461_ ( .A(\ID_EX_typ [3] ), .B1(_05480_ ), .B2(_05690_ ), .ZN(_05691_ ) );
XNOR2_X1 _13462_ ( .A(_03895_ ), .B(\ID_EX_pc [6] ), .ZN(_05692_ ) );
OAI21_X1 _13463_ ( .A(_05691_ ), .B1(_05480_ ), .B2(_05692_ ), .ZN(_05693_ ) );
BUF_X4 _13464_ ( .A(_05319_ ), .Z(_05694_ ) );
NOR2_X1 _13465_ ( .A1(_05290_ ), .A2(_05268_ ), .ZN(_05695_ ) );
AND3_X1 _13466_ ( .A1(_05246_ ), .A2(\mycsreg.CSReg[3][6] ), .A3(_05256_ ), .ZN(_05696_ ) );
AND3_X1 _13467_ ( .A1(_05246_ ), .A2(\mepc [6] ), .A3(_05251_ ), .ZN(_05697_ ) );
NOR2_X1 _13468_ ( .A1(_05696_ ), .A2(_05697_ ), .ZN(_05698_ ) );
AND3_X1 _13469_ ( .A1(_05234_ ), .A2(\mtvec [6] ), .A3(_05261_ ), .ZN(_05699_ ) );
AND3_X1 _13470_ ( .A1(_05234_ ), .A2(\mycsreg.CSReg[0][6] ), .A3(_05240_ ), .ZN(_05700_ ) );
NOR2_X1 _13471_ ( .A1(_05699_ ), .A2(_05700_ ), .ZN(_05701_ ) );
NAND3_X1 _13472_ ( .A1(_05695_ ), .A2(_05698_ ), .A3(_05701_ ), .ZN(_05702_ ) );
INV_X1 _13473_ ( .A(\EX_LS_result_csreg_mem [6] ), .ZN(_05703_ ) );
NAND3_X1 _13474_ ( .A1(_05366_ ), .A2(_05367_ ), .A3(_05703_ ), .ZN(_05704_ ) );
AND2_X1 _13475_ ( .A1(_05702_ ), .A2(_05704_ ), .ZN(_05705_ ) );
OAI211_X1 _13476_ ( .A(_05693_ ), .B(_05436_ ), .C1(_05694_ ), .C2(_05705_ ), .ZN(_05706_ ) );
XNOR2_X1 _13477_ ( .A(_05685_ ), .B(_02567_ ), .ZN(_05707_ ) );
AOI22_X1 _13478_ ( .A1(_05707_ ), .A2(_05427_ ), .B1(_05373_ ), .B2(_05690_ ), .ZN(_05708_ ) );
AOI21_X1 _13479_ ( .A(_05522_ ), .B1(_05706_ ), .B2(_05708_ ), .ZN(_00139_ ) );
INV_X1 _13480_ ( .A(\ID_EX_pc [5] ), .ZN(_05709_ ) );
XNOR2_X1 _13481_ ( .A(_03894_ ), .B(_05709_ ), .ZN(_05710_ ) );
AOI21_X1 _13482_ ( .A(\ID_EX_typ [3] ), .B1(_05301_ ), .B2(_05710_ ), .ZN(_05711_ ) );
OR2_X1 _13483_ ( .A1(_05123_ ), .A2(_05125_ ), .ZN(_05712_ ) );
NOR2_X1 _13484_ ( .A1(_05124_ ), .A2(_05127_ ), .ZN(_05713_ ) );
XNOR2_X1 _13485_ ( .A(_05712_ ), .B(_05713_ ), .ZN(_05714_ ) );
OAI21_X1 _13486_ ( .A(_05711_ ), .B1(_05320_ ), .B2(_05714_ ), .ZN(_05715_ ) );
NAND3_X1 _13487_ ( .A1(_05235_ ), .A2(\mycsreg.CSReg[0][5] ), .A3(_05241_ ), .ZN(_05716_ ) );
NAND3_X1 _13488_ ( .A1(_05235_ ), .A2(\mtvec [5] ), .A3(_05330_ ), .ZN(_05717_ ) );
AND2_X1 _13489_ ( .A1(_05716_ ), .A2(_05717_ ), .ZN(_05718_ ) );
INV_X1 _13490_ ( .A(_05268_ ), .ZN(_05719_ ) );
NAND3_X1 _13491_ ( .A1(_05247_ ), .A2(\mycsreg.CSReg[3][5] ), .A3(_05338_ ), .ZN(_05720_ ) );
NAND3_X1 _13492_ ( .A1(_05247_ ), .A2(\mepc [5] ), .A3(_05252_ ), .ZN(_05721_ ) );
AND2_X1 _13493_ ( .A1(_05720_ ), .A2(_05721_ ), .ZN(_05722_ ) );
NAND4_X1 _13494_ ( .A1(_05293_ ), .A2(_05718_ ), .A3(_05719_ ), .A4(_05722_ ), .ZN(_05723_ ) );
INV_X1 _13495_ ( .A(\EX_LS_result_csreg_mem [5] ), .ZN(_05724_ ) );
NAND3_X1 _13496_ ( .A1(_05386_ ), .A2(_05387_ ), .A3(_05724_ ), .ZN(_05725_ ) );
AND2_X1 _13497_ ( .A1(_05723_ ), .A2(_05725_ ), .ZN(_05726_ ) );
OAI211_X1 _13498_ ( .A(_05715_ ), .B(_05436_ ), .C1(_05694_ ), .C2(_05726_ ), .ZN(_05727_ ) );
NOR2_X1 _13499_ ( .A1(_05714_ ), .A2(_03879_ ), .ZN(_05728_ ) );
NOR2_X1 _13500_ ( .A1(_05683_ ), .A2(_02621_ ), .ZN(_05729_ ) );
XNOR2_X1 _13501_ ( .A(_05729_ ), .B(_02620_ ), .ZN(_05730_ ) );
AOI21_X1 _13502_ ( .A(_05728_ ), .B1(_05730_ ), .B2(_05427_ ), .ZN(_05731_ ) );
AOI21_X1 _13503_ ( .A(_05522_ ), .B1(_05727_ ), .B2(_05731_ ), .ZN(_00140_ ) );
BUF_X4 _13504_ ( .A(_05299_ ), .Z(_05732_ ) );
NAND3_X1 _13505_ ( .A1(_05469_ ), .A2(\mycsreg.CSReg[3][4] ), .A3(_05257_ ), .ZN(_05733_ ) );
NAND3_X1 _13506_ ( .A1(_05260_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_05378_ ), .ZN(_05734_ ) );
NAND3_X1 _13507_ ( .A1(_05327_ ), .A2(\mtvec [4] ), .A3(_05262_ ), .ZN(_05735_ ) );
NAND3_X1 _13508_ ( .A1(_05469_ ), .A2(\mepc [4] ), .A3(_05383_ ), .ZN(_05736_ ) );
AND4_X1 _13509_ ( .A1(_05733_ ), .A2(_05734_ ), .A3(_05735_ ), .A4(_05736_ ), .ZN(_05737_ ) );
AND2_X1 _13510_ ( .A1(_05737_ ), .A2(_05695_ ), .ZN(_05738_ ) );
INV_X1 _13511_ ( .A(\EX_LS_result_csreg_mem [4] ), .ZN(_05739_ ) );
AND3_X1 _13512_ ( .A1(_05386_ ), .A2(_05387_ ), .A3(_05739_ ), .ZN(_05740_ ) );
NOR2_X1 _13513_ ( .A1(_05738_ ), .A2(_05740_ ), .ZN(_05741_ ) );
XNOR2_X1 _13514_ ( .A(_03893_ ), .B(\ID_EX_pc [4] ), .ZN(_05742_ ) );
OAI21_X1 _13515_ ( .A(_05319_ ), .B1(_05480_ ), .B2(_05742_ ), .ZN(_05743_ ) );
AND3_X1 _13516_ ( .A1(_05120_ ), .A2(_05122_ ), .A3(_05111_ ), .ZN(_05744_ ) );
NOR2_X1 _13517_ ( .A1(_05744_ ), .A2(_05123_ ), .ZN(_05745_ ) );
AND3_X1 _13518_ ( .A1(_05104_ ), .A2(_05106_ ), .A3(_05745_ ), .ZN(_05746_ ) );
OAI221_X1 _13519_ ( .A(_05407_ ), .B1(_05377_ ), .B2(_05741_ ), .C1(_05743_ ), .C2(_05746_ ), .ZN(_05747_ ) );
XNOR2_X1 _13520_ ( .A(_02522_ ), .B(_02613_ ), .ZN(_05748_ ) );
AOI22_X1 _13521_ ( .A1(_05748_ ), .A2(_05427_ ), .B1(_05373_ ), .B2(_05745_ ), .ZN(_05749_ ) );
AOI21_X1 _13522_ ( .A(_05732_ ), .B1(_05747_ ), .B2(_05749_ ), .ZN(_00141_ ) );
XOR2_X1 _13523_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_pc [2] ), .Z(_05750_ ) );
XNOR2_X1 _13524_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_imm [3] ), .ZN(_05751_ ) );
XNOR2_X1 _13525_ ( .A(_05119_ ), .B(_05751_ ), .ZN(_05752_ ) );
MUX2_X1 _13526_ ( .A(_05750_ ), .B(_05752_ ), .S(_05224_ ), .Z(_05753_ ) );
OR2_X1 _13527_ ( .A1(_05753_ ), .A2(\ID_EX_typ [3] ), .ZN(_05754_ ) );
INV_X1 _13528_ ( .A(\EX_LS_result_csreg_mem [3] ), .ZN(_05755_ ) );
AND3_X1 _13529_ ( .A1(_05496_ ), .A2(_05497_ ), .A3(_05755_ ), .ZN(_05756_ ) );
NAND3_X1 _13530_ ( .A1(_05337_ ), .A2(\mycsreg.CSReg[3][3] ), .A3(_05339_ ), .ZN(_05757_ ) );
NAND3_X1 _13531_ ( .A1(_05328_ ), .A2(\mtvec [3] ), .A3(_05331_ ), .ZN(_05758_ ) );
NAND3_X1 _13532_ ( .A1(_05328_ ), .A2(\mycsreg.CSReg[0][3] ), .A3(_05242_ ), .ZN(_05759_ ) );
NAND3_X1 _13533_ ( .A1(_05337_ ), .A2(\mepc [3] ), .A3(_05253_ ), .ZN(_05760_ ) );
AND4_X1 _13534_ ( .A1(_05757_ ), .A2(_05758_ ), .A3(_05759_ ), .A4(_05760_ ), .ZN(_05761_ ) );
AOI21_X1 _13535_ ( .A(_05756_ ), .B1(_05761_ ), .B2(_05695_ ), .ZN(_05762_ ) );
OAI211_X1 _13536_ ( .A(_05754_ ), .B(_05376_ ), .C1(_05694_ ), .C2(_05762_ ), .ZN(_05763_ ) );
XNOR2_X1 _13537_ ( .A(_02494_ ), .B(_02517_ ), .ZN(_05764_ ) );
AOI22_X1 _13538_ ( .A1(_05764_ ), .A2(_05427_ ), .B1(_05373_ ), .B2(_05752_ ), .ZN(_05765_ ) );
AOI21_X1 _13539_ ( .A(_05732_ ), .B1(_05763_ ), .B2(_05765_ ), .ZN(_00142_ ) );
OR3_X1 _13540_ ( .A1(_05115_ ), .A2(_05116_ ), .A3(_05112_ ), .ZN(_05766_ ) );
AND2_X1 _13541_ ( .A1(_05766_ ), .A2(_05117_ ), .ZN(_05767_ ) );
MUX2_X1 _13542_ ( .A(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .B(_05767_ ), .S(_05223_ ), .Z(_05768_ ) );
OR2_X1 _13543_ ( .A1(_05768_ ), .A2(\ID_EX_typ [3] ), .ZN(_05769_ ) );
AND3_X1 _13544_ ( .A1(_05496_ ), .A2(_05497_ ), .A3(\EX_LS_result_csreg_mem [2] ), .ZN(_05770_ ) );
INV_X1 _13545_ ( .A(_05770_ ), .ZN(_05771_ ) );
NAND3_X1 _13546_ ( .A1(_05236_ ), .A2(\mycsreg.CSReg[0][2] ), .A3(_05242_ ), .ZN(_05772_ ) );
NAND4_X1 _13547_ ( .A1(_05333_ ), .A2(_05334_ ), .A3(_05383_ ), .A4(\mepc [2] ), .ZN(_05773_ ) );
NAND2_X1 _13548_ ( .A1(_05772_ ), .A2(_05773_ ), .ZN(_05774_ ) );
AND3_X1 _13549_ ( .A1(_05236_ ), .A2(\mtvec [2] ), .A3(_05331_ ), .ZN(_05775_ ) );
AND4_X1 _13550_ ( .A1(\mycsreg.CSReg[3][2] ), .A2(_05333_ ), .A3(_05334_ ), .A4(_05257_ ), .ZN(_05776_ ) );
NOR4_X1 _13551_ ( .A1(_05774_ ), .A2(_05775_ ), .A3(_05359_ ), .A4(_05776_ ), .ZN(_05777_ ) );
BUF_X4 _13552_ ( .A(_05291_ ), .Z(_05778_ ) );
OAI21_X1 _13553_ ( .A(_05771_ ), .B1(_05777_ ), .B2(_05778_ ), .ZN(_05779_ ) );
OAI211_X1 _13554_ ( .A(_05769_ ), .B(_05376_ ), .C1(_05694_ ), .C2(_05779_ ), .ZN(_05780_ ) );
OR3_X1 _13555_ ( .A1(_02490_ ), .A2(_02491_ ), .A3(_02443_ ), .ZN(_05781_ ) );
AND2_X1 _13556_ ( .A1(_05781_ ), .A2(_02492_ ), .ZN(_05782_ ) );
AOI22_X1 _13557_ ( .A1(_05782_ ), .A2(_05371_ ), .B1(_05373_ ), .B2(_05767_ ), .ZN(_05783_ ) );
AOI21_X1 _13558_ ( .A(_05732_ ), .B1(_05780_ ), .B2(_05783_ ), .ZN(_00143_ ) );
AND3_X1 _13559_ ( .A1(_05386_ ), .A2(_05387_ ), .A3(\EX_LS_result_csreg_mem [1] ), .ZN(_05784_ ) );
INV_X1 _13560_ ( .A(_05784_ ), .ZN(_05785_ ) );
NAND3_X1 _13561_ ( .A1(_05337_ ), .A2(\mycsreg.CSReg[3][1] ), .A3(_05339_ ), .ZN(_05786_ ) );
NAND3_X1 _13562_ ( .A1(_05328_ ), .A2(\mtvec [1] ), .A3(_05331_ ), .ZN(_05787_ ) );
NAND3_X1 _13563_ ( .A1(_05236_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_05242_ ), .ZN(_05788_ ) );
NAND3_X1 _13564_ ( .A1(_05248_ ), .A2(\mepc [1] ), .A3(_05253_ ), .ZN(_05789_ ) );
AND4_X1 _13565_ ( .A1(_05786_ ), .A2(_05787_ ), .A3(_05788_ ), .A4(_05789_ ), .ZN(_05790_ ) );
OAI21_X1 _13566_ ( .A(_05785_ ), .B1(_05790_ ), .B2(_05291_ ), .ZN(_05791_ ) );
XOR2_X1 _13567_ ( .A(_05113_ ), .B(_05114_ ), .Z(_05792_ ) );
INV_X1 _13568_ ( .A(_05792_ ), .ZN(_05793_ ) );
OAI21_X1 _13569_ ( .A(_05319_ ), .B1(_05320_ ), .B2(_05793_ ), .ZN(_05794_ ) );
INV_X1 _13570_ ( .A(\ID_EX_pc [1] ), .ZN(_05795_ ) );
AOI21_X1 _13571_ ( .A(_05795_ ), .B1(_05104_ ), .B2(_05106_ ), .ZN(_05796_ ) );
OAI221_X1 _13572_ ( .A(_05407_ ), .B1(_05377_ ), .B2(_05791_ ), .C1(_05794_ ), .C2(_05796_ ), .ZN(_05797_ ) );
XOR2_X1 _13573_ ( .A(_02466_ ), .B(_02489_ ), .Z(_05798_ ) );
AOI22_X1 _13574_ ( .A1(_05798_ ), .A2(_05371_ ), .B1(_05373_ ), .B2(_05792_ ), .ZN(_05799_ ) );
AOI21_X1 _13575_ ( .A(_05732_ ), .B1(_05797_ ), .B2(_05799_ ), .ZN(_00144_ ) );
NAND3_X1 _13576_ ( .A1(_05308_ ), .A2(\ID_EX_pc [26] ), .A3(_05311_ ), .ZN(_05800_ ) );
XNOR2_X1 _13577_ ( .A(_05800_ ), .B(_05210_ ), .ZN(_05801_ ) );
OR2_X1 _13578_ ( .A1(_05224_ ), .A2(_05801_ ), .ZN(_05802_ ) );
NAND2_X1 _13579_ ( .A1(_05205_ ), .A2(_05207_ ), .ZN(_05803_ ) );
NAND2_X1 _13580_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_05804_ ) );
NAND2_X1 _13581_ ( .A1(_05803_ ), .A2(_05804_ ), .ZN(_05805_ ) );
XNOR2_X1 _13582_ ( .A(_05805_ ), .B(_05206_ ), .ZN(_05806_ ) );
OAI211_X1 _13583_ ( .A(_05802_ ), .B(_05319_ ), .C1(_05320_ ), .C2(_05806_ ), .ZN(_05807_ ) );
NAND3_X1 _13584_ ( .A1(_05408_ ), .A2(\mycsreg.CSReg[0][27] ), .A3(_05241_ ), .ZN(_05808_ ) );
NAND3_X1 _13585_ ( .A1(_05336_ ), .A2(\mycsreg.CSReg[3][27] ), .A3(_05338_ ), .ZN(_05809_ ) );
AND2_X1 _13586_ ( .A1(_05808_ ), .A2(_05809_ ), .ZN(_05810_ ) );
NAND3_X1 _13587_ ( .A1(_05408_ ), .A2(\mtvec [27] ), .A3(_05330_ ), .ZN(_05811_ ) );
NAND3_X1 _13588_ ( .A1(_05247_ ), .A2(\mepc [27] ), .A3(_05252_ ), .ZN(_05812_ ) );
AND2_X1 _13589_ ( .A1(_05811_ ), .A2(_05812_ ), .ZN(_05813_ ) );
NAND4_X1 _13590_ ( .A1(_05292_ ), .A2(_05719_ ), .A3(_05810_ ), .A4(_05813_ ), .ZN(_05814_ ) );
INV_X1 _13591_ ( .A(\EX_LS_result_csreg_mem [27] ), .ZN(_05815_ ) );
NAND3_X1 _13592_ ( .A1(_05386_ ), .A2(_05387_ ), .A3(_05815_ ), .ZN(_05816_ ) );
AND2_X1 _13593_ ( .A1(_05814_ ), .A2(_05816_ ), .ZN(_05817_ ) );
OAI211_X1 _13594_ ( .A(_05807_ ), .B(_05376_ ), .C1(_05694_ ), .C2(_05817_ ), .ZN(_05818_ ) );
MUX2_X1 _13595_ ( .A(_05806_ ), .B(_03036_ ), .S(fanout_net_5 ), .Z(_05819_ ) );
OR2_X1 _13596_ ( .A1(_05819_ ), .A2(_05347_ ), .ZN(_05820_ ) );
AOI21_X1 _13597_ ( .A(_05732_ ), .B1(_05818_ ), .B2(_05820_ ), .ZN(_00145_ ) );
AND4_X1 _13598_ ( .A1(\mycsreg.CSReg[3][0] ), .A2(_05230_ ), .A3(_05245_ ), .A4(_05256_ ), .ZN(_05821_ ) );
NOR2_X1 _13599_ ( .A1(_05359_ ), .A2(_05821_ ), .ZN(_05822_ ) );
NAND3_X1 _13600_ ( .A1(_05336_ ), .A2(\mepc [0] ), .A3(_05252_ ), .ZN(_05823_ ) );
NAND3_X1 _13601_ ( .A1(_05408_ ), .A2(\mtvec [0] ), .A3(_05330_ ), .ZN(_05824_ ) );
NAND3_X1 _13602_ ( .A1(_05408_ ), .A2(\mycsreg.CSReg[0][0] ), .A3(_05241_ ), .ZN(_05825_ ) );
NAND4_X1 _13603_ ( .A1(_05822_ ), .A2(_05823_ ), .A3(_05824_ ), .A4(_05825_ ), .ZN(_05826_ ) );
NAND2_X1 _13604_ ( .A1(_05826_ ), .A2(_05292_ ), .ZN(_05827_ ) );
NAND3_X1 _13605_ ( .A1(_05366_ ), .A2(_05367_ ), .A3(\EX_LS_result_csreg_mem [0] ), .ZN(_05828_ ) );
AND2_X1 _13606_ ( .A1(_05827_ ), .A2(_05828_ ), .ZN(_05829_ ) );
INV_X1 _13607_ ( .A(_05829_ ), .ZN(_05830_ ) );
XOR2_X1 _13608_ ( .A(\ID_EX_pc [0] ), .B(\ID_EX_imm [0] ), .Z(_05831_ ) );
MUX2_X1 _13609_ ( .A(\ID_EX_pc [0] ), .B(_05831_ ), .S(_05223_ ), .Z(_05832_ ) );
MUX2_X1 _13610_ ( .A(_05830_ ), .B(_05832_ ), .S(_05318_ ), .Z(_05833_ ) );
AOI22_X1 _13611_ ( .A1(_05833_ ), .A2(_05325_ ), .B1(_05374_ ), .B2(_05831_ ), .ZN(_05834_ ) );
NOR2_X1 _13612_ ( .A1(_05834_ ), .A2(_05300_ ), .ZN(_00146_ ) );
XOR2_X1 _13613_ ( .A(_05312_ ), .B(\ID_EX_pc [26] ), .Z(_05835_ ) );
NAND2_X1 _13614_ ( .A1(_05302_ ), .A2(_05835_ ), .ZN(_05836_ ) );
XNOR2_X1 _13615_ ( .A(_05204_ ), .B(_05207_ ), .ZN(_05837_ ) );
INV_X1 _13616_ ( .A(_05837_ ), .ZN(_05838_ ) );
OAI211_X1 _13617_ ( .A(_05836_ ), .B(_05319_ ), .C1(_05302_ ), .C2(_05838_ ), .ZN(_05839_ ) );
BUF_X2 _13618_ ( .A(_05496_ ), .Z(_05840_ ) );
BUF_X2 _13619_ ( .A(_05497_ ), .Z(_05841_ ) );
NAND3_X1 _13620_ ( .A1(_05840_ ), .A2(_05841_ ), .A3(\EX_LS_result_csreg_mem [26] ), .ZN(_05842_ ) );
NAND3_X1 _13621_ ( .A1(_05337_ ), .A2(\mycsreg.CSReg[3][26] ), .A3(_05339_ ), .ZN(_05843_ ) );
NAND3_X1 _13622_ ( .A1(_05328_ ), .A2(\mtvec [26] ), .A3(_05331_ ), .ZN(_05844_ ) );
NAND3_X1 _13623_ ( .A1(_05236_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_05242_ ), .ZN(_05845_ ) );
NAND3_X1 _13624_ ( .A1(_05248_ ), .A2(\mepc [26] ), .A3(_05253_ ), .ZN(_05846_ ) );
AND4_X1 _13625_ ( .A1(_05843_ ), .A2(_05844_ ), .A3(_05845_ ), .A4(_05846_ ), .ZN(_05847_ ) );
OAI21_X1 _13626_ ( .A(_05842_ ), .B1(_05847_ ), .B2(_05778_ ), .ZN(_05848_ ) );
OAI211_X1 _13627_ ( .A(_05839_ ), .B(_05376_ ), .C1(_05694_ ), .C2(_05848_ ), .ZN(_05849_ ) );
BUF_X4 _13628_ ( .A(_03877_ ), .Z(_05850_ ) );
BUF_X4 _13629_ ( .A(_05850_ ), .Z(_05851_ ) );
AOI21_X1 _13630_ ( .A(_05851_ ), .B1(_03037_ ), .B2(_03034_ ), .ZN(_05852_ ) );
OAI21_X1 _13631_ ( .A(_03892_ ), .B1(_05837_ ), .B2(fanout_net_5 ), .ZN(_05853_ ) );
OR2_X1 _13632_ ( .A1(_05852_ ), .A2(_05853_ ), .ZN(_05854_ ) );
AOI21_X1 _13633_ ( .A(_05732_ ), .B1(_05849_ ), .B2(_05854_ ), .ZN(_00147_ ) );
AND3_X1 _13634_ ( .A1(_05310_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_05855_ ) );
AND2_X1 _13635_ ( .A1(_05308_ ), .A2(_05855_ ), .ZN(_05856_ ) );
AND3_X1 _13636_ ( .A1(_05856_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_05857_ ) );
NAND2_X1 _13637_ ( .A1(_05857_ ), .A2(\ID_EX_pc [24] ), .ZN(_05858_ ) );
XNOR2_X1 _13638_ ( .A(_05858_ ), .B(\ID_EX_pc [25] ), .ZN(_05859_ ) );
NAND2_X1 _13639_ ( .A1(_05302_ ), .A2(_05859_ ), .ZN(_05860_ ) );
OR2_X1 _13640_ ( .A1(_05183_ ), .A2(_05199_ ), .ZN(_05861_ ) );
AND2_X1 _13641_ ( .A1(_05861_ ), .A2(_05109_ ), .ZN(_05862_ ) );
OR2_X1 _13642_ ( .A1(_05862_ ), .A2(_05201_ ), .ZN(_05863_ ) );
XNOR2_X1 _13643_ ( .A(_05863_ ), .B(_05108_ ), .ZN(_05864_ ) );
OAI211_X1 _13644_ ( .A(_05860_ ), .B(_05319_ ), .C1(_05302_ ), .C2(_05864_ ), .ZN(_05865_ ) );
NAND3_X1 _13645_ ( .A1(_05496_ ), .A2(_05497_ ), .A3(\EX_LS_result_csreg_mem [25] ), .ZN(_05866_ ) );
NAND3_X1 _13646_ ( .A1(_05248_ ), .A2(\mycsreg.CSReg[3][25] ), .A3(_05339_ ), .ZN(_05867_ ) );
NAND3_X1 _13647_ ( .A1(_05236_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_05242_ ), .ZN(_05868_ ) );
NAND3_X1 _13648_ ( .A1(_05236_ ), .A2(\mtvec [25] ), .A3(_05331_ ), .ZN(_05869_ ) );
NAND3_X1 _13649_ ( .A1(_05248_ ), .A2(\mepc [25] ), .A3(_05253_ ), .ZN(_05870_ ) );
AND4_X1 _13650_ ( .A1(_05867_ ), .A2(_05868_ ), .A3(_05869_ ), .A4(_05870_ ), .ZN(_05871_ ) );
OAI21_X1 _13651_ ( .A(_05866_ ), .B1(_05871_ ), .B2(_05778_ ), .ZN(_05872_ ) );
OAI211_X1 _13652_ ( .A(_05865_ ), .B(_05376_ ), .C1(_05694_ ), .C2(_05872_ ), .ZN(_05873_ ) );
MUX2_X1 _13653_ ( .A(_05864_ ), .B(_03040_ ), .S(fanout_net_5 ), .Z(_05874_ ) );
OR2_X1 _13654_ ( .A1(_05874_ ), .A2(_05347_ ), .ZN(_05875_ ) );
AOI21_X1 _13655_ ( .A(_05732_ ), .B1(_05873_ ), .B2(_05875_ ), .ZN(_00148_ ) );
NAND3_X1 _13656_ ( .A1(_05856_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_05876_ ) );
XNOR2_X1 _13657_ ( .A(_05876_ ), .B(\ID_EX_pc [24] ), .ZN(_05877_ ) );
AOI21_X1 _13658_ ( .A(\ID_EX_typ [3] ), .B1(_05301_ ), .B2(_05877_ ), .ZN(_05878_ ) );
XOR2_X1 _13659_ ( .A(_05861_ ), .B(_05109_ ), .Z(_05879_ ) );
INV_X1 _13660_ ( .A(_05879_ ), .ZN(_05880_ ) );
OAI21_X1 _13661_ ( .A(_05878_ ), .B1(_05320_ ), .B2(_05880_ ), .ZN(_05881_ ) );
NAND3_X1 _13662_ ( .A1(_05248_ ), .A2(\mycsreg.CSReg[3][24] ), .A3(_05339_ ), .ZN(_05882_ ) );
NAND3_X1 _13663_ ( .A1(_05260_ ), .A2(\mycsreg.CSReg[0][24] ), .A3(_05378_ ), .ZN(_05883_ ) );
NAND3_X1 _13664_ ( .A1(_05260_ ), .A2(\mtvec [24] ), .A3(_05262_ ), .ZN(_05884_ ) );
NAND3_X1 _13665_ ( .A1(_05469_ ), .A2(\mepc [24] ), .A3(_05383_ ), .ZN(_05885_ ) );
AND4_X1 _13666_ ( .A1(_05882_ ), .A2(_05883_ ), .A3(_05884_ ), .A4(_05885_ ), .ZN(_05886_ ) );
AND2_X1 _13667_ ( .A1(_05573_ ), .A2(_05886_ ), .ZN(_05887_ ) );
INV_X1 _13668_ ( .A(\EX_LS_result_csreg_mem [24] ), .ZN(_05888_ ) );
AND3_X1 _13669_ ( .A1(_05386_ ), .A2(_05367_ ), .A3(_05888_ ), .ZN(_05889_ ) );
NOR2_X1 _13670_ ( .A1(_05887_ ), .A2(_05889_ ), .ZN(_05890_ ) );
OAI211_X1 _13671_ ( .A(_05881_ ), .B(_05376_ ), .C1(_05694_ ), .C2(_05890_ ), .ZN(_05891_ ) );
AOI22_X1 _13672_ ( .A1(_03041_ ), .A2(_05371_ ), .B1(_05373_ ), .B2(_05879_ ), .ZN(_05892_ ) );
AOI21_X1 _13673_ ( .A(_05732_ ), .B1(_05891_ ), .B2(_05892_ ), .ZN(_00149_ ) );
NAND3_X1 _13674_ ( .A1(_05308_ ), .A2(\ID_EX_pc [22] ), .A3(_05855_ ), .ZN(_05893_ ) );
XNOR2_X1 _13675_ ( .A(_05893_ ), .B(\ID_EX_pc [23] ), .ZN(_05894_ ) );
NAND2_X1 _13676_ ( .A1(_05302_ ), .A2(_05894_ ), .ZN(_05895_ ) );
INV_X1 _13677_ ( .A(_05170_ ), .ZN(_05896_ ) );
OAI21_X1 _13678_ ( .A(_05174_ ), .B1(_05352_ ), .B2(_05191_ ), .ZN(_05897_ ) );
AOI21_X1 _13679_ ( .A(_05896_ ), .B1(_05897_ ), .B2(_05198_ ), .ZN(_05898_ ) );
OR2_X1 _13680_ ( .A1(_05898_ ), .A2(_05193_ ), .ZN(_05899_ ) );
XNOR2_X1 _13681_ ( .A(_05899_ ), .B(_05169_ ), .ZN(_05900_ ) );
OAI211_X1 _13682_ ( .A(_05895_ ), .B(_05319_ ), .C1(_05302_ ), .C2(_05900_ ), .ZN(_05901_ ) );
NAND3_X1 _13683_ ( .A1(_05496_ ), .A2(_05497_ ), .A3(\EX_LS_result_csreg_mem [23] ), .ZN(_05902_ ) );
NAND3_X1 _13684_ ( .A1(_05337_ ), .A2(\mycsreg.CSReg[3][23] ), .A3(_05339_ ), .ZN(_05903_ ) );
NAND3_X1 _13685_ ( .A1(_05328_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_05242_ ), .ZN(_05904_ ) );
NAND3_X1 _13686_ ( .A1(_05328_ ), .A2(\mtvec [23] ), .A3(_05331_ ), .ZN(_05905_ ) );
NAND3_X1 _13687_ ( .A1(_05337_ ), .A2(\mepc [23] ), .A3(_05253_ ), .ZN(_05906_ ) );
AND4_X1 _13688_ ( .A1(_05903_ ), .A2(_05904_ ), .A3(_05905_ ), .A4(_05906_ ), .ZN(_05907_ ) );
OAI21_X1 _13689_ ( .A(_05902_ ), .B1(_05907_ ), .B2(_05291_ ), .ZN(_05908_ ) );
OAI211_X1 _13690_ ( .A(_05901_ ), .B(_05376_ ), .C1(_05694_ ), .C2(_05908_ ), .ZN(_05909_ ) );
MUX2_X1 _13691_ ( .A(_05900_ ), .B(_03048_ ), .S(fanout_net_5 ), .Z(_05910_ ) );
OR2_X1 _13692_ ( .A1(_05910_ ), .A2(_05347_ ), .ZN(_05911_ ) );
AOI21_X1 _13693_ ( .A(_05732_ ), .B1(_05909_ ), .B2(_05911_ ), .ZN(_00150_ ) );
INV_X1 _13694_ ( .A(\ID_EX_pc [22] ), .ZN(_05912_ ) );
XNOR2_X1 _13695_ ( .A(_05856_ ), .B(_05912_ ), .ZN(_05913_ ) );
NAND2_X1 _13696_ ( .A1(_05302_ ), .A2(_05913_ ), .ZN(_05914_ ) );
NAND2_X1 _13697_ ( .A1(_05897_ ), .A2(_05198_ ), .ZN(_05915_ ) );
XNOR2_X1 _13698_ ( .A(_05915_ ), .B(_05896_ ), .ZN(_05916_ ) );
INV_X1 _13699_ ( .A(_05916_ ), .ZN(_05917_ ) );
OAI211_X1 _13700_ ( .A(_05914_ ), .B(_05319_ ), .C1(_05302_ ), .C2(_05917_ ), .ZN(_05918_ ) );
INV_X1 _13701_ ( .A(\EX_LS_result_csreg_mem [22] ), .ZN(_05919_ ) );
AND3_X1 _13702_ ( .A1(_05496_ ), .A2(_05497_ ), .A3(_05919_ ), .ZN(_05920_ ) );
NAND3_X1 _13703_ ( .A1(_05337_ ), .A2(\mycsreg.CSReg[3][22] ), .A3(_05339_ ), .ZN(_05921_ ) );
NAND3_X1 _13704_ ( .A1(_05328_ ), .A2(\mycsreg.CSReg[0][22] ), .A3(_05242_ ), .ZN(_05922_ ) );
NAND3_X1 _13705_ ( .A1(_05328_ ), .A2(\mtvec [22] ), .A3(_05331_ ), .ZN(_05923_ ) );
NAND3_X1 _13706_ ( .A1(_05337_ ), .A2(\mepc [22] ), .A3(_05253_ ), .ZN(_05924_ ) );
AND4_X1 _13707_ ( .A1(_05921_ ), .A2(_05922_ ), .A3(_05923_ ), .A4(_05924_ ), .ZN(_05925_ ) );
AOI21_X1 _13708_ ( .A(_05920_ ), .B1(_05573_ ), .B2(_05925_ ), .ZN(_05926_ ) );
OAI211_X1 _13709_ ( .A(_05918_ ), .B(_05376_ ), .C1(_05694_ ), .C2(_05926_ ), .ZN(_05927_ ) );
BUF_X4 _13710_ ( .A(_05324_ ), .Z(_05928_ ) );
BUF_X4 _13711_ ( .A(_05850_ ), .Z(_05929_ ) );
BUF_X4 _13712_ ( .A(_05929_ ), .Z(_05930_ ) );
AOI21_X1 _13713_ ( .A(_05928_ ), .B1(_05917_ ), .B2(_05930_ ), .ZN(_05931_ ) );
BUF_X4 _13714_ ( .A(_05929_ ), .Z(_05932_ ) );
OAI21_X1 _13715_ ( .A(_05931_ ), .B1(_03049_ ), .B2(_05932_ ), .ZN(_05933_ ) );
AOI21_X1 _13716_ ( .A(_05732_ ), .B1(_05927_ ), .B2(_05933_ ), .ZN(_00151_ ) );
INV_X1 _13717_ ( .A(\ID_EX_pc [20] ), .ZN(_05934_ ) );
NOR2_X1 _13718_ ( .A1(_05349_ ), .A2(_05934_ ), .ZN(_05935_ ) );
INV_X1 _13719_ ( .A(\ID_EX_pc [21] ), .ZN(_05936_ ) );
XNOR2_X1 _13720_ ( .A(_05935_ ), .B(_05936_ ), .ZN(_05937_ ) );
AOI21_X1 _13721_ ( .A(\ID_EX_typ [3] ), .B1(_05301_ ), .B2(_05937_ ), .ZN(_05938_ ) );
OAI21_X1 _13722_ ( .A(_05173_ ), .B1(_05352_ ), .B2(_05191_ ), .ZN(_05939_ ) );
NAND2_X1 _13723_ ( .A1(\ID_EX_pc [20] ), .A2(\ID_EX_imm [20] ), .ZN(_05940_ ) );
NAND2_X1 _13724_ ( .A1(_05939_ ), .A2(_05940_ ), .ZN(_05941_ ) );
XNOR2_X1 _13725_ ( .A(_05941_ ), .B(_05172_ ), .ZN(_05942_ ) );
OAI21_X1 _13726_ ( .A(_05938_ ), .B1(_05320_ ), .B2(_05942_ ), .ZN(_05943_ ) );
NAND3_X1 _13727_ ( .A1(_05235_ ), .A2(\mycsreg.CSReg[0][21] ), .A3(_05241_ ), .ZN(_05944_ ) );
NAND4_X1 _13728_ ( .A1(_05333_ ), .A2(_05334_ ), .A3(_05252_ ), .A4(\mepc [21] ), .ZN(_05945_ ) );
AND2_X1 _13729_ ( .A1(_05944_ ), .A2(_05945_ ), .ZN(_05946_ ) );
AND3_X1 _13730_ ( .A1(_05235_ ), .A2(\mtvec [21] ), .A3(_05330_ ), .ZN(_05947_ ) );
INV_X1 _13731_ ( .A(_05947_ ), .ZN(_05948_ ) );
AND3_X1 _13732_ ( .A1(_05247_ ), .A2(\mycsreg.CSReg[3][21] ), .A3(_05338_ ), .ZN(_05949_ ) );
NOR2_X1 _13733_ ( .A1(_05949_ ), .A2(_05268_ ), .ZN(_05950_ ) );
NAND4_X1 _13734_ ( .A1(_05531_ ), .A2(_05946_ ), .A3(_05948_ ), .A4(_05950_ ), .ZN(_05951_ ) );
NOR3_X1 _13735_ ( .A1(_05463_ ), .A2(_05466_ ), .A3(\EX_LS_result_csreg_mem [21] ), .ZN(_05952_ ) );
INV_X1 _13736_ ( .A(_05952_ ), .ZN(_05953_ ) );
AND2_X1 _13737_ ( .A1(_05951_ ), .A2(_05953_ ), .ZN(_05954_ ) );
OAI211_X1 _13738_ ( .A(_05943_ ), .B(_05376_ ), .C1(_05377_ ), .C2(_05954_ ), .ZN(_05955_ ) );
NOR2_X1 _13739_ ( .A1(_03000_ ), .A2(_05403_ ), .ZN(_05956_ ) );
NOR2_X1 _13740_ ( .A1(_05942_ ), .A2(_03879_ ), .ZN(_05957_ ) );
NOR2_X1 _13741_ ( .A1(_05956_ ), .A2(_05957_ ), .ZN(_05958_ ) );
AOI21_X1 _13742_ ( .A(_05299_ ), .B1(_05955_ ), .B2(_05958_ ), .ZN(_00152_ ) );
NOR2_X1 _13743_ ( .A1(_02992_ ), .A2(_05403_ ), .ZN(_05959_ ) );
NOR2_X1 _13744_ ( .A1(_05220_ ), .A2(_05221_ ), .ZN(_05960_ ) );
AND2_X1 _13745_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_imm [30] ), .ZN(_05961_ ) );
NOR2_X1 _13746_ ( .A1(_05960_ ), .A2(_05961_ ), .ZN(_05962_ ) );
XNOR2_X1 _13747_ ( .A(\ID_EX_pc [31] ), .B(\ID_EX_imm [31] ), .ZN(_05963_ ) );
XNOR2_X1 _13748_ ( .A(_05962_ ), .B(_05963_ ), .ZN(_05964_ ) );
NAND3_X1 _13749_ ( .A1(_05235_ ), .A2(\mtvec [31] ), .A3(_05330_ ), .ZN(_05965_ ) );
NAND3_X1 _13750_ ( .A1(_05235_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_05241_ ), .ZN(_05966_ ) );
NAND3_X1 _13751_ ( .A1(_05247_ ), .A2(\mycsreg.CSReg[3][31] ), .A3(_05338_ ), .ZN(_05967_ ) );
NAND3_X1 _13752_ ( .A1(_05247_ ), .A2(\mepc [31] ), .A3(_05252_ ), .ZN(_05968_ ) );
NAND4_X1 _13753_ ( .A1(_05965_ ), .A2(_05966_ ), .A3(_05967_ ), .A4(_05968_ ), .ZN(_05969_ ) );
NAND2_X1 _13754_ ( .A1(_05292_ ), .A2(_05969_ ), .ZN(_05970_ ) );
NAND3_X1 _13755_ ( .A1(_05366_ ), .A2(_05367_ ), .A3(\EX_LS_result_csreg_mem [31] ), .ZN(_05971_ ) );
NAND3_X1 _13756_ ( .A1(_05970_ ), .A2(\ID_EX_typ [3] ), .A3(_05971_ ), .ZN(_05972_ ) );
NAND4_X1 _13757_ ( .A1(_05104_ ), .A2(_05324_ ), .A3(_05106_ ), .A4(_05972_ ), .ZN(_05973_ ) );
AOI21_X1 _13758_ ( .A(_05964_ ), .B1(_05973_ ), .B2(_03879_ ), .ZN(_05974_ ) );
NOR2_X1 _13759_ ( .A1(_03910_ ), .A2(_03911_ ), .ZN(_05975_ ) );
XNOR2_X1 _13760_ ( .A(_05975_ ), .B(\ID_EX_pc [31] ), .ZN(_05976_ ) );
OAI21_X2 _13761_ ( .A(_05318_ ), .B1(_05224_ ), .B2(_05976_ ), .ZN(_05977_ ) );
AND3_X2 _13762_ ( .A1(_05977_ ), .A2(_05324_ ), .A3(_05972_ ), .ZN(_05978_ ) );
OR4_X2 _13763_ ( .A1(_05299_ ), .A2(_05959_ ), .A3(_05974_ ), .A4(_05978_ ), .ZN(_00153_ ) );
AND3_X1 _13764_ ( .A1(_03891_ ), .A2(\ID_EX_pc [31] ), .A3(_03083_ ), .ZN(_00154_ ) );
AND3_X1 _13765_ ( .A1(_03891_ ), .A2(\ID_EX_pc [30] ), .A3(_03083_ ), .ZN(_00155_ ) );
CLKBUF_X2 _13766_ ( .A(_03065_ ), .Z(_05979_ ) );
AND3_X1 _13767_ ( .A1(_03891_ ), .A2(\ID_EX_pc [21] ), .A3(_05979_ ), .ZN(_00156_ ) );
AND3_X1 _13768_ ( .A1(_03891_ ), .A2(\ID_EX_pc [20] ), .A3(_05979_ ), .ZN(_00157_ ) );
AND3_X1 _13769_ ( .A1(_03891_ ), .A2(\ID_EX_pc [19] ), .A3(_05979_ ), .ZN(_00158_ ) );
CLKBUF_X2 _13770_ ( .A(_03890_ ), .Z(_05980_ ) );
AND3_X1 _13771_ ( .A1(_05980_ ), .A2(\ID_EX_pc [18] ), .A3(_05979_ ), .ZN(_00159_ ) );
AND3_X1 _13772_ ( .A1(_05980_ ), .A2(\ID_EX_pc [17] ), .A3(_05979_ ), .ZN(_00160_ ) );
AND3_X1 _13773_ ( .A1(_05980_ ), .A2(\ID_EX_pc [16] ), .A3(_05979_ ), .ZN(_00161_ ) );
AND3_X1 _13774_ ( .A1(_05980_ ), .A2(\ID_EX_pc [15] ), .A3(_05979_ ), .ZN(_00162_ ) );
AND3_X1 _13775_ ( .A1(_05980_ ), .A2(\ID_EX_pc [14] ), .A3(_05979_ ), .ZN(_00163_ ) );
AND3_X1 _13776_ ( .A1(_05980_ ), .A2(\ID_EX_pc [13] ), .A3(_05979_ ), .ZN(_00164_ ) );
AND3_X1 _13777_ ( .A1(_05980_ ), .A2(\ID_EX_pc [12] ), .A3(_05979_ ), .ZN(_00165_ ) );
CLKBUF_X2 _13778_ ( .A(_03065_ ), .Z(_05981_ ) );
AND3_X1 _13779_ ( .A1(_05980_ ), .A2(\ID_EX_pc [29] ), .A3(_05981_ ), .ZN(_00166_ ) );
AND3_X1 _13780_ ( .A1(_05980_ ), .A2(\ID_EX_pc [11] ), .A3(_05981_ ), .ZN(_00167_ ) );
AND3_X1 _13781_ ( .A1(_05980_ ), .A2(\ID_EX_pc [10] ), .A3(_05981_ ), .ZN(_00168_ ) );
CLKBUF_X2 _13782_ ( .A(_03885_ ), .Z(_05982_ ) );
AND3_X1 _13783_ ( .A1(_05982_ ), .A2(\ID_EX_pc [9] ), .A3(_05981_ ), .ZN(_00169_ ) );
AND3_X1 _13784_ ( .A1(_05982_ ), .A2(\ID_EX_pc [8] ), .A3(_05981_ ), .ZN(_00170_ ) );
AND3_X1 _13785_ ( .A1(_05982_ ), .A2(\ID_EX_pc [7] ), .A3(_05981_ ), .ZN(_00171_ ) );
AND3_X1 _13786_ ( .A1(_05982_ ), .A2(\ID_EX_pc [6] ), .A3(_05981_ ), .ZN(_00172_ ) );
AND3_X1 _13787_ ( .A1(_05982_ ), .A2(\ID_EX_pc [5] ), .A3(_05981_ ), .ZN(_00173_ ) );
AND3_X1 _13788_ ( .A1(_05982_ ), .A2(\ID_EX_pc [4] ), .A3(_05981_ ), .ZN(_00174_ ) );
AND3_X1 _13789_ ( .A1(_05982_ ), .A2(\ID_EX_pc [3] ), .A3(_05981_ ), .ZN(_00175_ ) );
CLKBUF_X2 _13790_ ( .A(_03065_ ), .Z(_05983_ ) );
AND3_X1 _13791_ ( .A1(_05982_ ), .A2(\ID_EX_pc [2] ), .A3(_05983_ ), .ZN(_00176_ ) );
AND3_X1 _13792_ ( .A1(_05982_ ), .A2(\ID_EX_pc [28] ), .A3(_05983_ ), .ZN(_00177_ ) );
AND3_X1 _13793_ ( .A1(_05982_ ), .A2(\ID_EX_pc [1] ), .A3(_05983_ ), .ZN(_00178_ ) );
CLKBUF_X2 _13794_ ( .A(_03885_ ), .Z(_05984_ ) );
AND3_X1 _13795_ ( .A1(_05984_ ), .A2(\ID_EX_pc [0] ), .A3(_05983_ ), .ZN(_00179_ ) );
AND3_X1 _13796_ ( .A1(_05984_ ), .A2(\ID_EX_pc [27] ), .A3(_05983_ ), .ZN(_00180_ ) );
AND3_X1 _13797_ ( .A1(_05984_ ), .A2(\ID_EX_pc [26] ), .A3(_05983_ ), .ZN(_00181_ ) );
AND3_X1 _13798_ ( .A1(_05984_ ), .A2(\ID_EX_pc [25] ), .A3(_05983_ ), .ZN(_00182_ ) );
AND3_X1 _13799_ ( .A1(_05984_ ), .A2(\ID_EX_pc [24] ), .A3(_05983_ ), .ZN(_00183_ ) );
AND3_X1 _13800_ ( .A1(_05984_ ), .A2(\ID_EX_pc [23] ), .A3(_05983_ ), .ZN(_00184_ ) );
AND3_X1 _13801_ ( .A1(_05984_ ), .A2(\ID_EX_pc [22] ), .A3(_05983_ ), .ZN(_00185_ ) );
CLKBUF_X2 _13802_ ( .A(_03065_ ), .Z(_05985_ ) );
AND3_X1 _13803_ ( .A1(_05984_ ), .A2(\ID_EX_typ [7] ), .A3(_05985_ ), .ZN(_00186_ ) );
INV_X1 _13804_ ( .A(io_master_awready ), .ZN(_05986_ ) );
NAND3_X1 _13805_ ( .A1(_02044_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .A3(_05986_ ), .ZN(_05987_ ) );
OAI21_X1 _13806_ ( .A(_05987_ ), .B1(\mylsu.state [4] ), .B2(\mylsu.state [0] ), .ZN(_05988_ ) );
OAI21_X1 _13807_ ( .A(_02069_ ), .B1(_03814_ ), .B2(io_master_arready ), .ZN(_05989_ ) );
INV_X1 _13808_ ( .A(_01966_ ), .ZN(_05990_ ) );
BUF_X2 _13809_ ( .A(_05990_ ), .Z(_05991_ ) );
NOR2_X1 _13810_ ( .A1(_05989_ ), .A2(_05991_ ), .ZN(_05992_ ) );
INV_X1 _13811_ ( .A(_05992_ ), .ZN(_05993_ ) );
AOI21_X1 _13812_ ( .A(_05988_ ), .B1(_05993_ ), .B2(_03844_ ), .ZN(_05994_ ) );
AND2_X1 _13813_ ( .A1(_03886_ ), .A2(EXU_valid_LSU ), .ZN(_05995_ ) );
INV_X1 _13814_ ( .A(_05995_ ), .ZN(_05996_ ) );
OAI22_X1 _13815_ ( .A1(_05994_ ), .A2(_05996_ ), .B1(_03873_ ), .B2(_05299_ ), .ZN(_00187_ ) );
AND3_X1 _13816_ ( .A1(_05984_ ), .A2(\ID_EX_typ [6] ), .A3(_05985_ ), .ZN(_00188_ ) );
AND3_X1 _13817_ ( .A1(_05984_ ), .A2(\ID_EX_typ [5] ), .A3(_05985_ ), .ZN(_00189_ ) );
AND3_X1 _13818_ ( .A1(_03890_ ), .A2(\ID_EX_typ [4] ), .A3(_05985_ ), .ZN(_00190_ ) );
AND3_X1 _13819_ ( .A1(_03890_ ), .A2(\ID_EX_typ [3] ), .A3(_05985_ ), .ZN(_00191_ ) );
AND3_X1 _13820_ ( .A1(_03890_ ), .A2(\ID_EX_typ [2] ), .A3(_05985_ ), .ZN(_00192_ ) );
AND3_X1 _13821_ ( .A1(_03890_ ), .A2(\ID_EX_typ [1] ), .A3(_05985_ ), .ZN(_00193_ ) );
AND3_X1 _13822_ ( .A1(_03890_ ), .A2(fanout_net_5 ), .A3(_05985_ ), .ZN(_00194_ ) );
AND2_X1 _13823_ ( .A1(_02059_ ), .A2(\myifu.myicache.valid_data_in ), .ZN(_05997_ ) );
CLKBUF_X2 _13824_ ( .A(_05997_ ), .Z(\myifu.wen_$_ANDNOT__A_Y ) );
NOR2_X2 _13825_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .ZN(_05998_ ) );
BUF_X2 _13826_ ( .A(_05998_ ), .Z(_05999_ ) );
AND3_X1 _13827_ ( .A1(_02059_ ), .A2(_05999_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(_00242_ ) );
AND3_X1 _13828_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_03745_ ), .A3(fanout_net_7 ), .ZN(_00243_ ) );
AND3_X1 _13829_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(fanout_net_11 ), .A3(_03753_ ), .ZN(_00244_ ) );
AND3_X1 _13830_ ( .A1(_03890_ ), .A2(\EX_LS_pc [2] ), .A3(_05985_ ), .ZN(_00282_ ) );
AND2_X1 _13831_ ( .A1(_03887_ ), .A2(\mylsu.state [3] ), .ZN(_00283_ ) );
INV_X1 _13832_ ( .A(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_06000_ ) );
AND3_X1 _13833_ ( .A1(_03885_ ), .A2(_06000_ ), .A3(_03065_ ), .ZN(_06001_ ) );
NOR2_X1 _13834_ ( .A1(\mylsu.state [3] ), .A2(\mylsu.state [1] ), .ZN(_06002_ ) );
NAND2_X1 _13835_ ( .A1(_06001_ ), .A2(_06002_ ), .ZN(_06003_ ) );
NOR2_X1 _13836_ ( .A1(_02041_ ), .A2(_03830_ ), .ZN(_06004_ ) );
OAI21_X1 _13837_ ( .A(_02042_ ), .B1(_02083_ ), .B2(_02084_ ), .ZN(_06005_ ) );
OR2_X1 _13838_ ( .A1(_06005_ ), .A2(_02087_ ), .ZN(_06006_ ) );
AOI21_X1 _13839_ ( .A(_03839_ ), .B1(_06006_ ), .B2(\EX_LS_flag [2] ), .ZN(_06007_ ) );
AOI21_X1 _13840_ ( .A(_06003_ ), .B1(_06004_ ), .B2(_06007_ ), .ZN(_00296_ ) );
NOR2_X1 _13841_ ( .A1(_02044_ ), .A2(_02049_ ), .ZN(_06008_ ) );
AOI21_X1 _13842_ ( .A(_02041_ ), .B1(_06006_ ), .B2(_06008_ ), .ZN(_06009_ ) );
AOI21_X1 _13843_ ( .A(_06003_ ), .B1(_06009_ ), .B2(_03845_ ), .ZN(_00297_ ) );
NOR2_X1 _13844_ ( .A1(_02085_ ), .A2(_02087_ ), .ZN(_06010_ ) );
NAND3_X1 _13845_ ( .A1(_06010_ ), .A2(\EX_LS_flag [2] ), .A3(_01989_ ), .ZN(_06011_ ) );
NOR2_X1 _13846_ ( .A1(_06011_ ), .A2(_06003_ ), .ZN(_00298_ ) );
NOR2_X1 _13847_ ( .A1(_02032_ ), .A2(_02033_ ), .ZN(_06012_ ) );
OR3_X1 _13848_ ( .A1(_06012_ ), .A2(\EX_LS_typ [4] ), .A3(_03862_ ), .ZN(_06013_ ) );
AND2_X1 _13849_ ( .A1(_06013_ ), .A2(_02040_ ), .ZN(_06014_ ) );
AOI21_X1 _13850_ ( .A(_06003_ ), .B1(_06014_ ), .B2(_03832_ ), .ZN(_00299_ ) );
AOI21_X1 _13851_ ( .A(_06003_ ), .B1(_03845_ ), .B2(_06011_ ), .ZN(_00300_ ) );
NAND3_X1 _13852_ ( .A1(_03887_ ), .A2(EXU_valid_LSU ), .A3(_06002_ ), .ZN(_06015_ ) );
OR3_X1 _13853_ ( .A1(_02054_ ), .A2(_03839_ ), .A3(_06015_ ), .ZN(_06016_ ) );
AND3_X1 _13854_ ( .A1(_06005_ ), .A2(_02086_ ), .A3(_06008_ ), .ZN(_06017_ ) );
AND2_X1 _13855_ ( .A1(_05993_ ), .A2(_06017_ ), .ZN(_06018_ ) );
OAI211_X1 _13856_ ( .A(_03844_ ), .B(_02035_ ), .C1(_06018_ ), .C2(_02039_ ), .ZN(_06019_ ) );
NOR2_X1 _13857_ ( .A1(_06017_ ), .A2(_02046_ ), .ZN(_06020_ ) );
AOI21_X1 _13858_ ( .A(_06016_ ), .B1(_06019_ ), .B2(_06020_ ), .ZN(_00301_ ) );
INV_X1 _13859_ ( .A(_00283_ ), .ZN(_06021_ ) );
INV_X1 _13860_ ( .A(_02046_ ), .ZN(_06022_ ) );
NAND3_X1 _13861_ ( .A1(_06022_ ), .A2(EXU_valid_LSU ), .A3(_06002_ ), .ZN(_06023_ ) );
OAI21_X1 _13862_ ( .A(_03887_ ), .B1(_03834_ ), .B2(_02090_ ), .ZN(_06024_ ) );
OAI21_X1 _13863_ ( .A(_06021_ ), .B1(_06023_ ), .B2(_06024_ ), .ZN(_00302_ ) );
BUF_X2 _13864_ ( .A(_02022_ ), .Z(\io_master_arburst [0] ) );
CLKBUF_X2 _13865_ ( .A(_01967_ ), .Z(_06025_ ) );
NOR3_X1 _13866_ ( .A1(_06025_ ), .A2(fanout_net_4 ), .A3(fanout_net_42 ), .ZN(_06026_ ) );
BUF_X4 _13867_ ( .A(_05991_ ), .Z(_06027_ ) );
BUF_X4 _13868_ ( .A(_06027_ ), .Z(_06028_ ) );
INV_X1 _13869_ ( .A(\mylsu.araddr_tmp [1] ), .ZN(_06029_ ) );
INV_X1 _13870_ ( .A(_01969_ ), .ZN(_06030_ ) );
AOI211_X1 _13871_ ( .A(_06026_ ), .B(_06028_ ), .C1(_06029_ ), .C2(_06030_ ), .ZN(\io_master_araddr [1] ) );
NOR3_X1 _13872_ ( .A1(_06025_ ), .A2(fanout_net_3 ), .A3(fanout_net_42 ), .ZN(_06031_ ) );
INV_X1 _13873_ ( .A(\mylsu.araddr_tmp [0] ), .ZN(_06032_ ) );
AOI211_X1 _13874_ ( .A(_06031_ ), .B(_06028_ ), .C1(_06032_ ), .C2(_06030_ ), .ZN(\io_master_araddr [0] ) );
OR3_X1 _13875_ ( .A1(_06025_ ), .A2(\EX_LS_dest_csreg_mem [15] ), .A3(fanout_net_42 ), .ZN(_06033_ ) );
BUF_X4 _13876_ ( .A(_01969_ ), .Z(_06034_ ) );
OAI21_X1 _13877_ ( .A(_06033_ ), .B1(_06034_ ), .B2(\mylsu.araddr_tmp [15] ), .ZN(_06035_ ) );
BUF_X4 _13878_ ( .A(_01972_ ), .Z(_06036_ ) );
BUF_X4 _13879_ ( .A(_06036_ ), .Z(_06037_ ) );
OAI22_X1 _13880_ ( .A1(_06028_ ), .A2(_06035_ ), .B1(_03653_ ), .B2(_06037_ ), .ZN(\io_master_araddr [15] ) );
OAI221_X1 _13881_ ( .A(\IF_ID_pc [14] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01947_ ), .C2(_01948_ ), .ZN(_06038_ ) );
INV_X1 _13882_ ( .A(_01956_ ), .ZN(_06039_ ) );
OR3_X1 _13883_ ( .A1(_06025_ ), .A2(\EX_LS_dest_csreg_mem [14] ), .A3(fanout_net_42 ), .ZN(_06040_ ) );
OAI211_X1 _13884_ ( .A(_06039_ ), .B(_06040_ ), .C1(\mylsu.araddr_tmp [14] ), .C2(_06034_ ), .ZN(_06041_ ) );
OAI21_X1 _13885_ ( .A(_06038_ ), .B1(\io_master_arburst [0] ), .B2(_06041_ ), .ZN(\io_master_araddr [14] ) );
OR3_X1 _13886_ ( .A1(_06025_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(fanout_net_42 ), .ZN(_06042_ ) );
OAI21_X1 _13887_ ( .A(_06042_ ), .B1(_06034_ ), .B2(\mylsu.araddr_tmp [5] ), .ZN(_06043_ ) );
OAI22_X1 _13888_ ( .A1(_06028_ ), .A2(_06043_ ), .B1(_03493_ ), .B2(_06037_ ), .ZN(\io_master_araddr [5] ) );
OR3_X1 _13889_ ( .A1(_06025_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(fanout_net_42 ), .ZN(_06044_ ) );
OAI21_X1 _13890_ ( .A(_06044_ ), .B1(_06034_ ), .B2(\mylsu.araddr_tmp [4] ), .ZN(_06045_ ) );
OAI22_X1 _13891_ ( .A1(_06028_ ), .A2(_06045_ ), .B1(_03745_ ), .B2(_06037_ ), .ZN(\io_master_araddr [4] ) );
OR3_X1 _13892_ ( .A1(_06025_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(fanout_net_42 ), .ZN(_06046_ ) );
OAI21_X1 _13893_ ( .A(_06046_ ), .B1(_06034_ ), .B2(\mylsu.araddr_tmp [3] ), .ZN(_06047_ ) );
OAI22_X1 _13894_ ( .A1(_06028_ ), .A2(_06047_ ), .B1(_03753_ ), .B2(_06037_ ), .ZN(\io_master_araddr [3] ) );
OAI221_X1 _13895_ ( .A(\IF_ID_pc [13] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01947_ ), .C2(_01948_ ), .ZN(_06048_ ) );
OR3_X1 _13896_ ( .A1(_01967_ ), .A2(\EX_LS_dest_csreg_mem [13] ), .A3(fanout_net_42 ), .ZN(_06049_ ) );
OAI211_X1 _13897_ ( .A(_06039_ ), .B(_06049_ ), .C1(\mylsu.araddr_tmp [13] ), .C2(_06034_ ), .ZN(_06050_ ) );
OAI21_X1 _13898_ ( .A(_06048_ ), .B1(\io_master_arburst [0] ), .B2(_06050_ ), .ZN(\io_master_araddr [13] ) );
OR3_X1 _13899_ ( .A1(_06025_ ), .A2(\EX_LS_dest_csreg_mem [12] ), .A3(fanout_net_42 ), .ZN(_06051_ ) );
OAI21_X1 _13900_ ( .A(_06051_ ), .B1(_06034_ ), .B2(\mylsu.araddr_tmp [12] ), .ZN(_06052_ ) );
OAI22_X1 _13901_ ( .A1(_06028_ ), .A2(_06052_ ), .B1(_01893_ ), .B2(_06037_ ), .ZN(\io_master_araddr [12] ) );
OAI221_X1 _13902_ ( .A(\IF_ID_pc [11] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01947_ ), .C2(_01948_ ), .ZN(_06053_ ) );
OR3_X1 _13903_ ( .A1(_01967_ ), .A2(\EX_LS_dest_csreg_mem [11] ), .A3(fanout_net_42 ), .ZN(_06054_ ) );
OAI211_X1 _13904_ ( .A(_06039_ ), .B(_06054_ ), .C1(\mylsu.araddr_tmp [11] ), .C2(_06034_ ), .ZN(_06055_ ) );
OAI21_X1 _13905_ ( .A(_06053_ ), .B1(\io_master_arburst [0] ), .B2(_06055_ ), .ZN(\io_master_araddr [11] ) );
NOR2_X1 _13906_ ( .A1(_01969_ ), .A2(\mylsu.araddr_tmp [10] ), .ZN(_06056_ ) );
NOR3_X1 _13907_ ( .A1(_01967_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(fanout_net_42 ), .ZN(_06057_ ) );
NOR3_X1 _13908_ ( .A1(_01956_ ), .A2(_06056_ ), .A3(_06057_ ), .ZN(_06058_ ) );
MUX2_X1 _13909_ ( .A(_06058_ ), .B(\IF_ID_pc [10] ), .S(\io_master_arburst [0] ), .Z(\io_master_araddr [10] ) );
NOR3_X1 _13910_ ( .A1(_06025_ ), .A2(_05273_ ), .A3(fanout_net_42 ), .ZN(_06059_ ) );
AOI21_X1 _13911_ ( .A(_06059_ ), .B1(_06030_ ), .B2(\mylsu.araddr_tmp [9] ), .ZN(_06060_ ) );
OAI22_X1 _13912_ ( .A1(_06028_ ), .A2(_06060_ ), .B1(_01913_ ), .B2(_06037_ ), .ZN(\io_master_araddr [9] ) );
NOR3_X1 _13913_ ( .A1(_06025_ ), .A2(_05274_ ), .A3(fanout_net_42 ), .ZN(_06061_ ) );
AOI21_X1 _13914_ ( .A(_06061_ ), .B1(_06030_ ), .B2(\mylsu.araddr_tmp [8] ), .ZN(_06062_ ) );
OAI22_X1 _13915_ ( .A1(_06028_ ), .A2(_06062_ ), .B1(_01886_ ), .B2(_06037_ ), .ZN(\io_master_araddr [8] ) );
OAI221_X1 _13916_ ( .A(\IF_ID_pc [7] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01947_ ), .C2(_01948_ ), .ZN(_06063_ ) );
OR3_X1 _13917_ ( .A1(_01967_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(fanout_net_42 ), .ZN(_06064_ ) );
OAI211_X1 _13918_ ( .A(_06039_ ), .B(_06064_ ), .C1(\mylsu.araddr_tmp [7] ), .C2(_06034_ ), .ZN(_06065_ ) );
OAI21_X1 _13919_ ( .A(_06063_ ), .B1(\io_master_arburst [0] ), .B2(_06065_ ), .ZN(\io_master_araddr [7] ) );
OAI221_X1 _13920_ ( .A(\IF_ID_pc [6] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01947_ ), .C2(_01948_ ), .ZN(_06066_ ) );
OR3_X1 _13921_ ( .A1(_01967_ ), .A2(\EX_LS_dest_csreg_mem [6] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06067_ ) );
OAI211_X1 _13922_ ( .A(_06039_ ), .B(_06067_ ), .C1(\mylsu.araddr_tmp [6] ), .C2(_06034_ ), .ZN(_06068_ ) );
OAI21_X1 _13923_ ( .A(_06066_ ), .B1(\io_master_arburst [0] ), .B2(_06068_ ), .ZN(\io_master_araddr [6] ) );
OR3_X1 _13924_ ( .A1(_01967_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06069_ ) );
OAI211_X1 _13925_ ( .A(_06039_ ), .B(_06069_ ), .C1(\mylsu.araddr_tmp [2] ), .C2(_01969_ ), .ZN(_06070_ ) );
NOR2_X1 _13926_ ( .A1(_01951_ ), .A2(_06070_ ), .ZN(_06071_ ) );
BUF_X4 _13927_ ( .A(_06071_ ), .Z(_06072_ ) );
BUF_X2 _13928_ ( .A(_06072_ ), .Z(\io_master_araddr [2] ) );
BUF_X2 _13929_ ( .A(_01966_ ), .Z(_06073_ ) );
CLKBUF_X2 _13930_ ( .A(_06073_ ), .Z(\io_master_arid [1] ) );
NOR3_X1 _13931_ ( .A1(\io_master_arburst [0] ), .A2(_02027_ ), .A3(_01956_ ), .ZN(\io_master_arsize [2] ) );
NOR3_X1 _13932_ ( .A1(\io_master_arburst [0] ), .A2(_02026_ ), .A3(_01956_ ), .ZN(\io_master_arsize [0] ) );
INV_X1 _13933_ ( .A(\EX_LS_typ [2] ), .ZN(_06074_ ) );
OAI22_X1 _13934_ ( .A1(_01949_ ), .A2(_01950_ ), .B1(_06074_ ), .B2(_01956_ ), .ZN(\io_master_arsize [1] ) );
AOI211_X1 _13935_ ( .A(_02058_ ), .B(_02060_ ), .C1(_02065_ ), .C2(_02068_ ), .ZN(io_master_arvalid ) );
AND2_X1 _13936_ ( .A1(\mylsu.state [0] ), .A2(EXU_valid_LSU ), .ZN(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ) );
AND2_X1 _13937_ ( .A1(_02045_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(_06075_ ) );
BUF_X4 _13938_ ( .A(_06075_ ), .Z(_06076_ ) );
BUF_X4 _13939_ ( .A(_06076_ ), .Z(_06077_ ) );
MUX2_X1 _13940_ ( .A(\mylsu.awaddr_tmp [31] ), .B(\EX_LS_dest_csreg_mem [31] ), .S(_06077_ ), .Z(\io_master_awaddr [31] ) );
MUX2_X1 _13941_ ( .A(\mylsu.awaddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_06077_ ), .Z(\io_master_awaddr [30] ) );
MUX2_X1 _13942_ ( .A(\mylsu.awaddr_tmp [21] ), .B(\EX_LS_dest_csreg_mem [21] ), .S(_06077_ ), .Z(\io_master_awaddr [21] ) );
MUX2_X1 _13943_ ( .A(\mylsu.awaddr_tmp [20] ), .B(\EX_LS_dest_csreg_mem [20] ), .S(_06077_ ), .Z(\io_master_awaddr [20] ) );
MUX2_X1 _13944_ ( .A(\mylsu.awaddr_tmp [19] ), .B(\EX_LS_dest_csreg_mem [19] ), .S(_06077_ ), .Z(\io_master_awaddr [19] ) );
MUX2_X1 _13945_ ( .A(\mylsu.awaddr_tmp [18] ), .B(\EX_LS_dest_csreg_mem [18] ), .S(_06077_ ), .Z(\io_master_awaddr [18] ) );
MUX2_X1 _13946_ ( .A(\mylsu.awaddr_tmp [17] ), .B(\EX_LS_dest_csreg_mem [17] ), .S(_06077_ ), .Z(\io_master_awaddr [17] ) );
MUX2_X1 _13947_ ( .A(\mylsu.awaddr_tmp [16] ), .B(\EX_LS_dest_csreg_mem [16] ), .S(_06077_ ), .Z(\io_master_awaddr [16] ) );
MUX2_X1 _13948_ ( .A(\mylsu.awaddr_tmp [15] ), .B(\EX_LS_dest_csreg_mem [15] ), .S(_06077_ ), .Z(\io_master_awaddr [15] ) );
BUF_X4 _13949_ ( .A(_06076_ ), .Z(_06078_ ) );
MUX2_X1 _13950_ ( .A(\mylsu.awaddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_06078_ ), .Z(\io_master_awaddr [14] ) );
MUX2_X1 _13951_ ( .A(\mylsu.awaddr_tmp [13] ), .B(\EX_LS_dest_csreg_mem [13] ), .S(_06078_ ), .Z(\io_master_awaddr [13] ) );
MUX2_X1 _13952_ ( .A(\mylsu.awaddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_06078_ ), .Z(\io_master_awaddr [12] ) );
MUX2_X1 _13953_ ( .A(\mylsu.awaddr_tmp [29] ), .B(\EX_LS_dest_csreg_mem [29] ), .S(_06078_ ), .Z(\io_master_awaddr [29] ) );
MUX2_X1 _13954_ ( .A(\mylsu.awaddr_tmp [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_06078_ ), .Z(\io_master_awaddr [11] ) );
MUX2_X1 _13955_ ( .A(\mylsu.awaddr_tmp [10] ), .B(\EX_LS_dest_csreg_mem [10] ), .S(_06078_ ), .Z(\io_master_awaddr [10] ) );
MUX2_X1 _13956_ ( .A(\mylsu.awaddr_tmp [9] ), .B(\EX_LS_dest_csreg_mem [9] ), .S(_06078_ ), .Z(\io_master_awaddr [9] ) );
MUX2_X1 _13957_ ( .A(\mylsu.awaddr_tmp [8] ), .B(\EX_LS_dest_csreg_mem [8] ), .S(_06078_ ), .Z(\io_master_awaddr [8] ) );
MUX2_X1 _13958_ ( .A(\mylsu.awaddr_tmp [7] ), .B(\EX_LS_dest_csreg_mem [7] ), .S(_06078_ ), .Z(\io_master_awaddr [7] ) );
MUX2_X1 _13959_ ( .A(\mylsu.awaddr_tmp [6] ), .B(\EX_LS_dest_csreg_mem [6] ), .S(_06078_ ), .Z(\io_master_awaddr [6] ) );
BUF_X4 _13960_ ( .A(_06076_ ), .Z(_06079_ ) );
MUX2_X1 _13961_ ( .A(\mylsu.awaddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_06079_ ), .Z(\io_master_awaddr [5] ) );
MUX2_X1 _13962_ ( .A(\mylsu.awaddr_tmp [4] ), .B(\EX_LS_dest_csreg_mem [4] ), .S(_06079_ ), .Z(\io_master_awaddr [4] ) );
MUX2_X1 _13963_ ( .A(\mylsu.awaddr_tmp [3] ), .B(\EX_LS_dest_csreg_mem [3] ), .S(_06079_ ), .Z(\io_master_awaddr [3] ) );
MUX2_X1 _13964_ ( .A(\mylsu.awaddr_tmp [2] ), .B(\EX_LS_dest_csreg_mem [2] ), .S(_06079_ ), .Z(\io_master_awaddr [2] ) );
MUX2_X1 _13965_ ( .A(\mylsu.awaddr_tmp [28] ), .B(\EX_LS_dest_csreg_mem [28] ), .S(_06079_ ), .Z(\io_master_awaddr [28] ) );
MUX2_X1 _13966_ ( .A(\mylsu.awaddr_tmp [1] ), .B(fanout_net_4 ), .S(_06079_ ), .Z(\io_master_awaddr [1] ) );
MUX2_X1 _13967_ ( .A(\mylsu.awaddr_tmp [0] ), .B(fanout_net_3 ), .S(_06079_ ), .Z(\io_master_awaddr [0] ) );
MUX2_X1 _13968_ ( .A(\mylsu.awaddr_tmp [27] ), .B(\EX_LS_dest_csreg_mem [27] ), .S(_06079_ ), .Z(\io_master_awaddr [27] ) );
MUX2_X1 _13969_ ( .A(\mylsu.awaddr_tmp [26] ), .B(\EX_LS_dest_csreg_mem [26] ), .S(_06079_ ), .Z(\io_master_awaddr [26] ) );
MUX2_X1 _13970_ ( .A(\mylsu.awaddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_06079_ ), .Z(\io_master_awaddr [25] ) );
MUX2_X1 _13971_ ( .A(\mylsu.awaddr_tmp [24] ), .B(\EX_LS_dest_csreg_mem [24] ), .S(_06076_ ), .Z(\io_master_awaddr [24] ) );
MUX2_X1 _13972_ ( .A(\mylsu.awaddr_tmp [23] ), .B(\EX_LS_dest_csreg_mem [23] ), .S(_06076_ ), .Z(\io_master_awaddr [23] ) );
MUX2_X1 _13973_ ( .A(\mylsu.awaddr_tmp [22] ), .B(\EX_LS_dest_csreg_mem [22] ), .S(_06076_ ), .Z(\io_master_awaddr [22] ) );
NAND4_X1 _13974_ ( .A1(_02050_ ), .A2(\EX_LS_typ [0] ), .A3(_03848_ ), .A4(_02030_ ), .ZN(\io_master_awsize [1] ) );
NOR2_X1 _13975_ ( .A1(\io_master_awsize [1] ), .A2(_02026_ ), .ZN(\io_master_awsize [0] ) );
AND3_X1 _13976_ ( .A1(_06014_ ), .A2(_02055_ ), .A3(_06076_ ), .ZN(_06080_ ) );
OR2_X1 _13977_ ( .A1(_06080_ ), .A2(\mylsu.state [4] ), .ZN(io_master_awvalid ) );
OR4_X1 _13978_ ( .A1(\mylsu.state [2] ), .A2(_06080_ ), .A3(\mylsu.state [4] ), .A4(\mylsu.state [1] ), .ZN(io_master_bready ) );
NOR3_X1 _13979_ ( .A1(_01955_ ), .A2(\mylsu.state [1] ), .A3(\mylsu.state [0] ), .ZN(_06081_ ) );
NOR2_X1 _13980_ ( .A1(\io_master_bresp [1] ), .A2(\io_master_bresp [0] ), .ZN(_06082_ ) );
AND2_X1 _13981_ ( .A1(_06082_ ), .A2(io_master_bvalid ), .ZN(_06083_ ) );
NAND2_X1 _13982_ ( .A1(\io_master_bid [1] ), .A2(\io_master_bid [0] ), .ZN(_06084_ ) );
NOR3_X1 _13983_ ( .A1(_06084_ ), .A2(\io_master_bid [3] ), .A3(\io_master_bid [2] ), .ZN(_06085_ ) );
AND2_X1 _13984_ ( .A1(_06083_ ), .A2(_06085_ ), .ZN(_06086_ ) );
INV_X1 _13985_ ( .A(_06086_ ), .ZN(_06087_ ) );
NOR2_X1 _13986_ ( .A1(_03818_ ), .A2(\io_master_rid [0] ), .ZN(_06088_ ) );
AND4_X1 _13987_ ( .A1(io_master_rlast ), .A2(_06088_ ), .A3(_03819_ ), .A4(_03820_ ), .ZN(_06089_ ) );
OAI21_X1 _13988_ ( .A(_06073_ ), .B1(_03817_ ), .B2(_06089_ ), .ZN(_06090_ ) );
AOI21_X1 _13989_ ( .A(_06090_ ), .B1(_03807_ ), .B2(_03806_ ), .ZN(_06091_ ) );
INV_X1 _13990_ ( .A(_06091_ ), .ZN(_06092_ ) );
AOI221_X4 _13991_ ( .A(_06081_ ), .B1(\mylsu.state [1] ), .B2(_06087_ ), .C1(_06092_ ), .C2(\mylsu.state [3] ), .ZN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
AOI211_X1 _13992_ ( .A(_02070_ ), .B(_02072_ ), .C1(_02065_ ), .C2(_02068_ ), .ZN(io_master_rready ) );
MUX2_X1 _13993_ ( .A(\EX_LS_result_csreg_mem [15] ), .B(\EX_LS_result_csreg_mem [7] ), .S(fanout_net_3 ), .Z(_06093_ ) );
INV_X1 _13994_ ( .A(fanout_net_4 ), .ZN(_06094_ ) );
CLKBUF_X2 _13995_ ( .A(_06094_ ), .Z(_06095_ ) );
AND2_X1 _13996_ ( .A1(_06093_ ), .A2(_06095_ ), .ZN(\io_master_wdata [15] ) );
MUX2_X1 _13997_ ( .A(\EX_LS_result_csreg_mem [14] ), .B(\EX_LS_result_csreg_mem [6] ), .S(fanout_net_3 ), .Z(_06096_ ) );
AND2_X1 _13998_ ( .A1(_06096_ ), .A2(_06095_ ), .ZN(\io_master_wdata [14] ) );
NOR3_X1 _13999_ ( .A1(_05724_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [5] ) );
NOR3_X1 _14000_ ( .A1(_05739_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [4] ) );
NOR3_X1 _14001_ ( .A1(_05755_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [3] ) );
INV_X1 _14002_ ( .A(\EX_LS_result_csreg_mem [2] ), .ZN(_06097_ ) );
NOR3_X1 _14003_ ( .A1(_06097_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [2] ) );
INV_X1 _14004_ ( .A(\EX_LS_result_csreg_mem [1] ), .ZN(_06098_ ) );
NOR3_X1 _14005_ ( .A1(_06098_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [1] ) );
INV_X1 _14006_ ( .A(\EX_LS_result_csreg_mem [0] ), .ZN(_06099_ ) );
NOR3_X1 _14007_ ( .A1(_06099_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [0] ) );
MUX2_X1 _14008_ ( .A(\EX_LS_result_csreg_mem [13] ), .B(\EX_LS_result_csreg_mem [5] ), .S(fanout_net_3 ), .Z(_06100_ ) );
AND2_X1 _14009_ ( .A1(_06100_ ), .A2(_06095_ ), .ZN(\io_master_wdata [13] ) );
MUX2_X1 _14010_ ( .A(\EX_LS_result_csreg_mem [12] ), .B(\EX_LS_result_csreg_mem [4] ), .S(fanout_net_3 ), .Z(_06101_ ) );
AND2_X1 _14011_ ( .A1(_06101_ ), .A2(_06095_ ), .ZN(\io_master_wdata [12] ) );
MUX2_X1 _14012_ ( .A(\EX_LS_result_csreg_mem [11] ), .B(\EX_LS_result_csreg_mem [3] ), .S(fanout_net_3 ), .Z(_06102_ ) );
AND2_X1 _14013_ ( .A1(_06102_ ), .A2(_06095_ ), .ZN(\io_master_wdata [11] ) );
MUX2_X1 _14014_ ( .A(\EX_LS_result_csreg_mem [10] ), .B(\EX_LS_result_csreg_mem [2] ), .S(fanout_net_3 ), .Z(_06103_ ) );
AND2_X1 _14015_ ( .A1(_06103_ ), .A2(_06095_ ), .ZN(\io_master_wdata [10] ) );
MUX2_X1 _14016_ ( .A(\EX_LS_result_csreg_mem [9] ), .B(\EX_LS_result_csreg_mem [1] ), .S(fanout_net_3 ), .Z(_06104_ ) );
AND2_X1 _14017_ ( .A1(_06104_ ), .A2(_06095_ ), .ZN(\io_master_wdata [9] ) );
MUX2_X1 _14018_ ( .A(\EX_LS_result_csreg_mem [8] ), .B(\EX_LS_result_csreg_mem [0] ), .S(fanout_net_3 ), .Z(_06105_ ) );
AND2_X1 _14019_ ( .A1(_06105_ ), .A2(_06095_ ), .ZN(\io_master_wdata [8] ) );
INV_X1 _14020_ ( .A(\EX_LS_result_csreg_mem [7] ), .ZN(_06106_ ) );
NOR3_X1 _14021_ ( .A1(_06106_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [7] ) );
NOR3_X1 _14022_ ( .A1(_05703_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [6] ) );
MUX2_X1 _14023_ ( .A(\EX_LS_result_csreg_mem [31] ), .B(\EX_LS_result_csreg_mem [23] ), .S(fanout_net_3 ), .Z(_06107_ ) );
MUX2_X1 _14024_ ( .A(_06107_ ), .B(_06093_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [31] ) );
MUX2_X1 _14025_ ( .A(\EX_LS_result_csreg_mem [30] ), .B(\EX_LS_result_csreg_mem [22] ), .S(fanout_net_3 ), .Z(_06108_ ) );
MUX2_X1 _14026_ ( .A(_06108_ ), .B(_06096_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [30] ) );
INV_X1 _14027_ ( .A(\EX_LS_result_csreg_mem [21] ), .ZN(_06109_ ) );
INV_X1 _14028_ ( .A(\EX_LS_result_csreg_mem [13] ), .ZN(_06110_ ) );
MUX2_X1 _14029_ ( .A(_06109_ ), .B(_06110_ ), .S(fanout_net_3 ), .Z(_06111_ ) );
NOR2_X1 _14030_ ( .A1(_06094_ ), .A2(fanout_net_3 ), .ZN(_06112_ ) );
INV_X1 _14031_ ( .A(_06112_ ), .ZN(_06113_ ) );
OAI22_X1 _14032_ ( .A1(_06111_ ), .A2(fanout_net_4 ), .B1(_06113_ ), .B2(_05724_ ), .ZN(\io_master_wdata [21] ) );
INV_X1 _14033_ ( .A(\EX_LS_result_csreg_mem [20] ), .ZN(_06114_ ) );
MUX2_X1 _14034_ ( .A(_06114_ ), .B(_05558_ ), .S(fanout_net_3 ), .Z(_06115_ ) );
OAI22_X1 _14035_ ( .A1(_06115_ ), .A2(fanout_net_4 ), .B1(_06113_ ), .B2(_05739_ ), .ZN(\io_master_wdata [20] ) );
INV_X1 _14036_ ( .A(fanout_net_3 ), .ZN(_06116_ ) );
OAI21_X1 _14037_ ( .A(_06094_ ), .B1(_06116_ ), .B2(\EX_LS_result_csreg_mem [11] ), .ZN(_06117_ ) );
NOR2_X1 _14038_ ( .A1(fanout_net_3 ), .A2(\EX_LS_result_csreg_mem [19] ), .ZN(_06118_ ) );
OAI22_X1 _14039_ ( .A1(_06113_ ), .A2(_05755_ ), .B1(_06117_ ), .B2(_06118_ ), .ZN(\io_master_wdata [19] ) );
INV_X1 _14040_ ( .A(\EX_LS_result_csreg_mem [18] ), .ZN(_06119_ ) );
INV_X1 _14041_ ( .A(\EX_LS_result_csreg_mem [10] ), .ZN(_06120_ ) );
MUX2_X1 _14042_ ( .A(_06119_ ), .B(_06120_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06121_ ) );
OAI22_X1 _14043_ ( .A1(_06121_ ), .A2(fanout_net_4 ), .B1(_06113_ ), .B2(_06097_ ), .ZN(\io_master_wdata [18] ) );
OAI21_X1 _14044_ ( .A(_06094_ ), .B1(_06116_ ), .B2(\EX_LS_result_csreg_mem [9] ), .ZN(_06122_ ) );
NOR2_X1 _14045_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [17] ), .ZN(_06123_ ) );
OAI22_X1 _14046_ ( .A1(_06113_ ), .A2(_06098_ ), .B1(_06122_ ), .B2(_06123_ ), .ZN(\io_master_wdata [17] ) );
INV_X1 _14047_ ( .A(\EX_LS_result_csreg_mem [16] ), .ZN(_06124_ ) );
MUX2_X1 _14048_ ( .A(_06124_ ), .B(_05653_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06125_ ) );
OAI22_X1 _14049_ ( .A1(_06125_ ), .A2(fanout_net_4 ), .B1(_06113_ ), .B2(_06099_ ), .ZN(\io_master_wdata [16] ) );
MUX2_X1 _14050_ ( .A(\EX_LS_result_csreg_mem [29] ), .B(\EX_LS_result_csreg_mem [21] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06126_ ) );
MUX2_X1 _14051_ ( .A(_06126_ ), .B(_06100_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [29] ) );
MUX2_X1 _14052_ ( .A(\EX_LS_result_csreg_mem [28] ), .B(\EX_LS_result_csreg_mem [20] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06127_ ) );
MUX2_X1 _14053_ ( .A(_06127_ ), .B(_06101_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [28] ) );
MUX2_X1 _14054_ ( .A(\EX_LS_result_csreg_mem [27] ), .B(\EX_LS_result_csreg_mem [19] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06128_ ) );
MUX2_X1 _14055_ ( .A(_06128_ ), .B(_06102_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [27] ) );
MUX2_X1 _14056_ ( .A(\EX_LS_result_csreg_mem [26] ), .B(\EX_LS_result_csreg_mem [18] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06129_ ) );
MUX2_X1 _14057_ ( .A(_06129_ ), .B(_06103_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [26] ) );
MUX2_X1 _14058_ ( .A(\EX_LS_result_csreg_mem [25] ), .B(\EX_LS_result_csreg_mem [17] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06130_ ) );
MUX2_X1 _14059_ ( .A(_06130_ ), .B(_06104_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [25] ) );
MUX2_X1 _14060_ ( .A(\EX_LS_result_csreg_mem [24] ), .B(\EX_LS_result_csreg_mem [16] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06131_ ) );
MUX2_X1 _14061_ ( .A(_06131_ ), .B(_06105_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [24] ) );
OAI21_X1 _14062_ ( .A(_06094_ ), .B1(_06116_ ), .B2(\EX_LS_result_csreg_mem [15] ), .ZN(_06132_ ) );
NOR2_X1 _14063_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [23] ), .ZN(_06133_ ) );
OAI22_X1 _14064_ ( .A1(_06113_ ), .A2(_06106_ ), .B1(_06132_ ), .B2(_06133_ ), .ZN(\io_master_wdata [23] ) );
INV_X1 _14065_ ( .A(\EX_LS_result_csreg_mem [14] ), .ZN(_06134_ ) );
MUX2_X1 _14066_ ( .A(_05919_ ), .B(_06134_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06135_ ) );
OAI22_X1 _14067_ ( .A1(_06135_ ), .A2(fanout_net_4 ), .B1(_06113_ ), .B2(_05703_ ), .ZN(\io_master_wdata [22] ) );
MUX2_X1 _14068_ ( .A(\EX_LS_typ [1] ), .B(\EX_LS_typ [0] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06136_ ) );
AND2_X1 _14069_ ( .A1(_06136_ ), .A2(_06095_ ), .ZN(\io_master_wstrb [1] ) );
AND3_X1 _14070_ ( .A1(_06116_ ), .A2(_06095_ ), .A3(\EX_LS_typ [0] ), .ZN(\io_master_wstrb [0] ) );
MUX2_X1 _14071_ ( .A(\EX_LS_typ [3] ), .B(\EX_LS_typ [2] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06137_ ) );
MUX2_X1 _14072_ ( .A(_06137_ ), .B(_06136_ ), .S(fanout_net_4 ), .Z(\io_master_wstrb [3] ) );
NAND3_X1 _14073_ ( .A1(_06094_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_typ [1] ), .ZN(_06138_ ) );
NAND3_X1 _14074_ ( .A1(_06116_ ), .A2(fanout_net_4 ), .A3(\EX_LS_typ [0] ), .ZN(_06139_ ) );
OAI211_X1 _14075_ ( .A(_06138_ ), .B(_06139_ ), .C1(_02025_ ), .C2(_06074_ ), .ZN(\io_master_wstrb [2] ) );
OR2_X1 _14076_ ( .A1(_06080_ ), .A2(\mylsu.state [2] ), .ZN(io_master_wvalid ) );
MUX2_X1 _14077_ ( .A(\LS_WB_wdata_csreg [2] ), .B(\LS_WB_wen_csreg [2] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14078_ ( .A(\LS_WB_wdata_csreg [1] ), .B(\LS_WB_wen_csreg [1] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14079_ ( .A(\LS_WB_wdata_csreg [0] ), .B(\LS_WB_wen_csreg [0] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14080_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\LS_WB_wen_csreg [3] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ) );
NOR2_X1 _14081_ ( .A1(\LS_WB_waddr_csreg [5] ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_06140_ ) );
AND2_X1 _14082_ ( .A1(\LS_WB_waddr_csreg [9] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_06141_ ) );
NOR2_X1 _14083_ ( .A1(\LS_WB_waddr_csreg [7] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_06142_ ) );
NOR2_X1 _14084_ ( .A1(\LS_WB_waddr_csreg [11] ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_06143_ ) );
AND4_X1 _14085_ ( .A1(_06140_ ), .A2(_06141_ ), .A3(_06142_ ), .A4(_06143_ ), .ZN(_06144_ ) );
AND2_X1 _14086_ ( .A1(_01547_ ), .A2(\LS_WB_wen_csreg [7] ), .ZN(_06145_ ) );
INV_X1 _14087_ ( .A(\LS_WB_waddr_csreg [0] ), .ZN(_06146_ ) );
NOR3_X1 _14088_ ( .A1(_06146_ ), .A2(\LS_WB_waddr_csreg [3] ), .A3(\LS_WB_waddr_csreg [1] ), .ZN(_06147_ ) );
AND4_X1 _14089_ ( .A1(\LS_WB_waddr_csreg [2] ), .A2(_06144_ ), .A3(_06145_ ), .A4(_06147_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ) );
NOR3_X1 _14090_ ( .A1(\LS_WB_waddr_csreg [3] ), .A2(\LS_WB_waddr_csreg [2] ), .A3(\LS_WB_waddr_csreg [7] ), .ZN(_06148_ ) );
AND3_X1 _14091_ ( .A1(_06148_ ), .A2(\LS_WB_waddr_csreg [6] ), .A3(_06140_ ), .ZN(_06149_ ) );
INV_X1 _14092_ ( .A(_06149_ ), .ZN(_06150_ ) );
NAND3_X1 _14093_ ( .A1(_06145_ ), .A2(_06143_ ), .A3(_06141_ ), .ZN(_06151_ ) );
NOR4_X1 _14094_ ( .A1(_06150_ ), .A2(\LS_WB_waddr_csreg [1] ), .A3(_06146_ ), .A4(_06151_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ) );
AND2_X1 _14095_ ( .A1(_06141_ ), .A2(_06143_ ), .ZN(_06152_ ) );
AND4_X1 _14096_ ( .A1(\LS_WB_waddr_csreg [6] ), .A2(_06152_ ), .A3(_06140_ ), .A4(_06148_ ), .ZN(_06153_ ) );
AND4_X1 _14097_ ( .A1(\LS_WB_waddr_csreg [1] ), .A2(_06153_ ), .A3(_06146_ ), .A4(_06145_ ), .ZN(_06154_ ) );
OR2_X1 _14098_ ( .A1(_06154_ ), .A2(_00093_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__B_Y_$_ORNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
AND3_X1 _14099_ ( .A1(_06145_ ), .A2(_06143_ ), .A3(_06141_ ), .ZN(_06155_ ) );
NOR4_X1 _14100_ ( .A1(\LS_WB_waddr_csreg [3] ), .A2(\LS_WB_waddr_csreg [2] ), .A3(\LS_WB_waddr_csreg [1] ), .A4(\LS_WB_waddr_csreg [0] ), .ZN(_06156_ ) );
AND4_X1 _14101_ ( .A1(_06140_ ), .A2(_06155_ ), .A3(_06142_ ), .A4(_06156_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _14102_ ( .A(_02057_ ), .ZN(_06157_ ) );
NOR2_X1 _14103_ ( .A1(_06010_ ), .A2(exception_quest_IDU ), .ZN(_06158_ ) );
NOR2_X1 _14104_ ( .A1(_06157_ ), .A2(_06158_ ), .ZN(_06159_ ) );
BUF_X4 _14105_ ( .A(_06159_ ), .Z(_06160_ ) );
MUX2_X1 _14106_ ( .A(\EX_LS_pc [21] ), .B(\ID_EX_pc [21] ), .S(_06160_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _14107_ ( .A(\EX_LS_pc [20] ), .B(\ID_EX_pc [20] ), .S(_06160_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _14108_ ( .A(\EX_LS_pc [19] ), .B(\ID_EX_pc [19] ), .S(_06160_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _14109_ ( .A(\EX_LS_pc [18] ), .B(\ID_EX_pc [18] ), .S(_06160_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _14110_ ( .A(\EX_LS_pc [17] ), .B(\ID_EX_pc [17] ), .S(_06160_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _14111_ ( .A(\EX_LS_pc [16] ), .B(\ID_EX_pc [16] ), .S(_06160_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _14112_ ( .A(\EX_LS_pc [15] ), .B(\ID_EX_pc [15] ), .S(_06160_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _14113_ ( .A(\EX_LS_pc [14] ), .B(\ID_EX_pc [14] ), .S(_06160_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _14114_ ( .A(\EX_LS_pc [13] ), .B(\ID_EX_pc [13] ), .S(_06160_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _14115_ ( .A(\EX_LS_pc [12] ), .B(\ID_EX_pc [12] ), .S(_06160_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ) );
BUF_X4 _14116_ ( .A(_06159_ ), .Z(_06161_ ) );
MUX2_X1 _14117_ ( .A(\EX_LS_pc [30] ), .B(\ID_EX_pc [30] ), .S(_06161_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14118_ ( .A(\EX_LS_pc [11] ), .B(\ID_EX_pc [11] ), .S(_06161_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _14119_ ( .A(\EX_LS_pc [10] ), .B(\ID_EX_pc [10] ), .S(_06161_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _14120_ ( .A(\EX_LS_pc [9] ), .B(\ID_EX_pc [9] ), .S(_06161_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _14121_ ( .A(\EX_LS_pc [8] ), .B(\ID_EX_pc [8] ), .S(_06161_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _14122_ ( .A(\EX_LS_pc [7] ), .B(\ID_EX_pc [7] ), .S(_06161_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _14123_ ( .A(\EX_LS_pc [6] ), .B(\ID_EX_pc [6] ), .S(_06161_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _14124_ ( .A(\EX_LS_pc [5] ), .B(\ID_EX_pc [5] ), .S(_06161_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _14125_ ( .A(\EX_LS_pc [4] ), .B(\ID_EX_pc [4] ), .S(_06161_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _14126_ ( .A(\EX_LS_pc [3] ), .B(\ID_EX_pc [3] ), .S(_06161_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ) );
BUF_X4 _14127_ ( .A(_06159_ ), .Z(_06162_ ) );
MUX2_X1 _14128_ ( .A(\EX_LS_pc [2] ), .B(\ID_EX_pc [2] ), .S(_06162_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _14129_ ( .A(\EX_LS_pc [29] ), .B(\ID_EX_pc [29] ), .S(_06162_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14130_ ( .A(\EX_LS_pc [1] ), .B(\ID_EX_pc [1] ), .S(_06162_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _14131_ ( .A(\EX_LS_pc [0] ), .B(\ID_EX_pc [0] ), .S(_06162_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _14132_ ( .A(\EX_LS_pc [28] ), .B(\ID_EX_pc [28] ), .S(_06162_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14133_ ( .A(\EX_LS_pc [27] ), .B(\ID_EX_pc [27] ), .S(_06162_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _14134_ ( .A(\EX_LS_pc [26] ), .B(\ID_EX_pc [26] ), .S(_06162_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _14135_ ( .A(\EX_LS_pc [25] ), .B(\ID_EX_pc [25] ), .S(_06162_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _14136_ ( .A(\EX_LS_pc [24] ), .B(\ID_EX_pc [24] ), .S(_06162_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _14137_ ( .A(\EX_LS_pc [23] ), .B(\ID_EX_pc [23] ), .S(_06162_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _14138_ ( .A(\EX_LS_pc [22] ), .B(\ID_EX_pc [22] ), .S(_06159_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _14139_ ( .A(\EX_LS_pc [31] ), .B(\ID_EX_pc [31] ), .S(_06159_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_D ) );
INV_X1 _14140_ ( .A(_02080_ ), .ZN(_06163_ ) );
NOR4_X1 _14141_ ( .A1(_06157_ ), .A2(exception_quest_IDU ), .A3(_06163_ ), .A4(_06158_ ), .ZN(_06164_ ) );
XOR2_X1 _14142_ ( .A(\mepc [23] ), .B(\myec.mepc_tmp [23] ), .Z(_06165_ ) );
XOR2_X1 _14143_ ( .A(\mepc [20] ), .B(\myec.mepc_tmp [20] ), .Z(_06166_ ) );
XOR2_X1 _14144_ ( .A(\mepc [22] ), .B(\myec.mepc_tmp [22] ), .Z(_06167_ ) );
XOR2_X1 _14145_ ( .A(\mepc [21] ), .B(\myec.mepc_tmp [21] ), .Z(_06168_ ) );
OR4_X1 _14146_ ( .A1(_06165_ ), .A2(_06166_ ), .A3(_06167_ ), .A4(_06168_ ), .ZN(_06169_ ) );
XOR2_X1 _14147_ ( .A(\mepc [16] ), .B(\myec.mepc_tmp [16] ), .Z(_06170_ ) );
XNOR2_X1 _14148_ ( .A(\mepc [19] ), .B(\myec.mepc_tmp [19] ), .ZN(_06171_ ) );
XNOR2_X1 _14149_ ( .A(\mepc [18] ), .B(\myec.mepc_tmp [18] ), .ZN(_06172_ ) );
NAND2_X1 _14150_ ( .A1(_06171_ ), .A2(_06172_ ), .ZN(_06173_ ) );
XOR2_X1 _14151_ ( .A(\mepc [17] ), .B(\myec.mepc_tmp [17] ), .Z(_06174_ ) );
NOR4_X1 _14152_ ( .A1(_06169_ ), .A2(_06170_ ), .A3(_06173_ ), .A4(_06174_ ), .ZN(_06175_ ) );
XNOR2_X1 _14153_ ( .A(\mepc [31] ), .B(\myec.mepc_tmp [31] ), .ZN(_06176_ ) );
XNOR2_X1 _14154_ ( .A(\mepc [30] ), .B(\myec.mepc_tmp [30] ), .ZN(_06177_ ) );
XNOR2_X1 _14155_ ( .A(\mepc [28] ), .B(\myec.mepc_tmp [28] ), .ZN(_06178_ ) );
XNOR2_X1 _14156_ ( .A(\mepc [29] ), .B(\myec.mepc_tmp [29] ), .ZN(_06179_ ) );
AND4_X1 _14157_ ( .A1(_06176_ ), .A2(_06177_ ), .A3(_06178_ ), .A4(_06179_ ), .ZN(_06180_ ) );
XNOR2_X1 _14158_ ( .A(\mepc [24] ), .B(\myec.mepc_tmp [24] ), .ZN(_06181_ ) );
XNOR2_X1 _14159_ ( .A(\mepc [26] ), .B(\myec.mepc_tmp [26] ), .ZN(_06182_ ) );
XNOR2_X1 _14160_ ( .A(\mepc [27] ), .B(\myec.mepc_tmp [27] ), .ZN(_06183_ ) );
XNOR2_X1 _14161_ ( .A(\mepc [25] ), .B(\myec.mepc_tmp [25] ), .ZN(_06184_ ) );
AND4_X1 _14162_ ( .A1(_06181_ ), .A2(_06182_ ), .A3(_06183_ ), .A4(_06184_ ), .ZN(_06185_ ) );
AND3_X1 _14163_ ( .A1(_06175_ ), .A2(_06180_ ), .A3(_06185_ ), .ZN(_06186_ ) );
XNOR2_X1 _14164_ ( .A(\mepc [2] ), .B(\myec.mepc_tmp [2] ), .ZN(_06187_ ) );
XNOR2_X1 _14165_ ( .A(\mepc [3] ), .B(\myec.mepc_tmp [3] ), .ZN(_06188_ ) );
XNOR2_X1 _14166_ ( .A(\mepc [1] ), .B(\myec.mepc_tmp [1] ), .ZN(_06189_ ) );
XNOR2_X1 _14167_ ( .A(\mepc [0] ), .B(\myec.mepc_tmp [0] ), .ZN(_06190_ ) );
NAND4_X1 _14168_ ( .A1(_06187_ ), .A2(_06188_ ), .A3(_06189_ ), .A4(_06190_ ), .ZN(_06191_ ) );
XNOR2_X1 _14169_ ( .A(\mepc [14] ), .B(\myec.mepc_tmp [14] ), .ZN(_06192_ ) );
XNOR2_X1 _14170_ ( .A(\mepc [12] ), .B(\myec.mepc_tmp [12] ), .ZN(_06193_ ) );
XNOR2_X1 _14171_ ( .A(\mepc [15] ), .B(\myec.mepc_tmp [15] ), .ZN(_06194_ ) );
XNOR2_X1 _14172_ ( .A(\mepc [13] ), .B(\myec.mepc_tmp [13] ), .ZN(_06195_ ) );
NAND4_X1 _14173_ ( .A1(_06192_ ), .A2(_06193_ ), .A3(_06194_ ), .A4(_06195_ ), .ZN(_06196_ ) );
XNOR2_X1 _14174_ ( .A(\mepc [8] ), .B(\myec.mepc_tmp [8] ), .ZN(_06197_ ) );
XNOR2_X1 _14175_ ( .A(\mepc [10] ), .B(\myec.mepc_tmp [10] ), .ZN(_06198_ ) );
XNOR2_X1 _14176_ ( .A(\mepc [11] ), .B(\myec.mepc_tmp [11] ), .ZN(_06199_ ) );
XNOR2_X1 _14177_ ( .A(\mepc [9] ), .B(\myec.mepc_tmp [9] ), .ZN(_06200_ ) );
NAND4_X1 _14178_ ( .A1(_06197_ ), .A2(_06198_ ), .A3(_06199_ ), .A4(_06200_ ), .ZN(_06201_ ) );
XNOR2_X1 _14179_ ( .A(\mepc [7] ), .B(\myec.mepc_tmp [7] ), .ZN(_06202_ ) );
XNOR2_X1 _14180_ ( .A(\mepc [6] ), .B(\myec.mepc_tmp [6] ), .ZN(_06203_ ) );
XNOR2_X1 _14181_ ( .A(\mepc [4] ), .B(\myec.mepc_tmp [4] ), .ZN(_06204_ ) );
XNOR2_X1 _14182_ ( .A(\mepc [5] ), .B(\myec.mepc_tmp [5] ), .ZN(_06205_ ) );
NAND4_X1 _14183_ ( .A1(_06202_ ), .A2(_06203_ ), .A3(_06204_ ), .A4(_06205_ ), .ZN(_06206_ ) );
NOR4_X1 _14184_ ( .A1(_06191_ ), .A2(_06196_ ), .A3(_06201_ ), .A4(_06206_ ), .ZN(_06207_ ) );
NAND3_X1 _14185_ ( .A1(_06186_ ), .A2(excp_written ), .A3(_06207_ ), .ZN(_06208_ ) );
AOI21_X1 _14186_ ( .A(_06164_ ), .B1(_06163_ ), .B2(_06208_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E ) );
NAND2_X1 _14187_ ( .A1(_05798_ ), .A2(_03003_ ), .ZN(_06209_ ) );
INV_X1 _14188_ ( .A(\ID_EX_typ [5] ), .ZN(_06210_ ) );
AND2_X2 _14189_ ( .A1(_02993_ ), .A2(_06210_ ), .ZN(_06211_ ) );
INV_X1 _14190_ ( .A(_06211_ ), .ZN(_06212_ ) );
BUF_X4 _14191_ ( .A(_06212_ ), .Z(_06213_ ) );
BUF_X4 _14192_ ( .A(_06213_ ), .Z(_06214_ ) );
OAI21_X1 _14193_ ( .A(_06209_ ), .B1(_05249_ ), .B2(_06214_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ) );
NOR4_X1 _14194_ ( .A1(_03341_ ), .A2(_03881_ ), .A3(\ID_EX_typ [5] ), .A4(\ID_EX_csr [0] ), .ZN(_06215_ ) );
XNOR2_X1 _14195_ ( .A(_04331_ ), .B(\ID_EX_imm [0] ), .ZN(_06216_ ) );
AOI21_X1 _14196_ ( .A(_06215_ ), .B1(_06216_ ), .B2(_03003_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ) );
AND2_X2 _14197_ ( .A1(_03354_ ), .A2(\ID_EX_typ [7] ), .ZN(_06217_ ) );
INV_X2 _14198_ ( .A(_06217_ ), .ZN(_06218_ ) );
BUF_X4 _14199_ ( .A(_06218_ ), .Z(_06219_ ) );
AND2_X1 _14200_ ( .A1(_05628_ ), .A2(_06219_ ), .ZN(_06220_ ) );
BUF_X4 _14201_ ( .A(_06212_ ), .Z(_06221_ ) );
MUX2_X1 _14202_ ( .A(\ID_EX_csr [10] ), .B(_06220_ ), .S(_06221_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ) );
BUF_X4 _14203_ ( .A(_06211_ ), .Z(_06222_ ) );
BUF_X4 _14204_ ( .A(_06222_ ), .Z(_06223_ ) );
AOI22_X1 _14205_ ( .A1(_05650_ ), .A2(_03003_ ), .B1(_05227_ ), .B2(_06223_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ) );
NOR2_X1 _14206_ ( .A1(_05666_ ), .A2(_02993_ ), .ZN(_06224_ ) );
BUF_X4 _14207_ ( .A(_06211_ ), .Z(_06225_ ) );
BUF_X4 _14208_ ( .A(_06225_ ), .Z(_06226_ ) );
AOI21_X1 _14209_ ( .A(_06224_ ), .B1(_05228_ ), .B2(_06226_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ) );
NAND2_X1 _14210_ ( .A1(_05688_ ), .A2(_03002_ ), .ZN(_06227_ ) );
OAI21_X1 _14211_ ( .A(_06227_ ), .B1(_05244_ ), .B2(_06214_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ) );
OR2_X1 _14212_ ( .A1(_05707_ ), .A2(_06217_ ), .ZN(_06228_ ) );
MUX2_X1 _14213_ ( .A(\ID_EX_csr [6] ), .B(_06228_ ), .S(_06221_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ) );
NAND2_X1 _14214_ ( .A1(_05730_ ), .A2(_03002_ ), .ZN(_06229_ ) );
OAI21_X1 _14215_ ( .A(_06229_ ), .B1(_05264_ ), .B2(_06214_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ) );
AND2_X1 _14216_ ( .A1(_05748_ ), .A2(_06218_ ), .ZN(_06230_ ) );
MUX2_X1 _14217_ ( .A(\ID_EX_csr [4] ), .B(_06230_ ), .S(_06221_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ) );
NAND2_X1 _14218_ ( .A1(_05764_ ), .A2(_03002_ ), .ZN(_06231_ ) );
OAI21_X1 _14219_ ( .A(_06231_ ), .B1(_05237_ ), .B2(_06214_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ) );
NAND3_X1 _14220_ ( .A1(_05781_ ), .A2(_03002_ ), .A3(_02492_ ), .ZN(_06232_ ) );
OAI21_X1 _14221_ ( .A(_06232_ ), .B1(_05238_ ), .B2(_06214_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ) );
AND2_X1 _14222_ ( .A1(_05588_ ), .A2(_06218_ ), .ZN(_06233_ ) );
MUX2_X1 _14223_ ( .A(\ID_EX_csr [11] ), .B(_06233_ ), .S(_06221_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ) );
BUF_X4 _14224_ ( .A(_04769_ ), .Z(_06234_ ) );
OAI22_X1 _14225_ ( .A1(_05954_ ), .A2(_06234_ ), .B1(_05850_ ), .B2(\ID_EX_imm [21] ), .ZN(_06235_ ) );
AOI21_X1 _14226_ ( .A(_06235_ ), .B1(_05930_ ), .B2(_04978_ ), .ZN(_06236_ ) );
NOR2_X2 _14227_ ( .A1(_04767_ ), .A2(\ID_EX_typ [2] ), .ZN(_06237_ ) );
BUF_X4 _14228_ ( .A(_06237_ ), .Z(_06238_ ) );
NAND3_X1 _14229_ ( .A1(_05951_ ), .A2(_06238_ ), .A3(_05953_ ), .ZN(_06239_ ) );
INV_X1 _14230_ ( .A(_06239_ ), .ZN(_06240_ ) );
OAI21_X1 _14231_ ( .A(_06223_ ), .B1(_06236_ ), .B2(_06240_ ), .ZN(_06241_ ) );
MUX2_X1 _14232_ ( .A(_05936_ ), .B(_04510_ ), .S(_06219_ ), .Z(_06242_ ) );
OAI21_X1 _14233_ ( .A(_06241_ ), .B1(_06226_ ), .B2(_06242_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ) );
OAI22_X1 _14234_ ( .A1(_05369_ ), .A2(_06234_ ), .B1(_05850_ ), .B2(\ID_EX_imm [20] ), .ZN(_06243_ ) );
INV_X1 _14235_ ( .A(_02294_ ), .ZN(_06244_ ) );
AOI21_X1 _14236_ ( .A(_06243_ ), .B1(_05930_ ), .B2(_06244_ ), .ZN(_06245_ ) );
BUF_X2 _14237_ ( .A(_05463_ ), .Z(_06246_ ) );
BUF_X2 _14238_ ( .A(_05466_ ), .Z(_06247_ ) );
OR3_X1 _14239_ ( .A1(_06246_ ), .A2(\EX_LS_result_csreg_mem [20] ), .A3(_06247_ ), .ZN(_06248_ ) );
INV_X1 _14240_ ( .A(_05357_ ), .ZN(_06249_ ) );
NAND4_X1 _14241_ ( .A1(_06249_ ), .A2(_05444_ ), .A3(_05362_ ), .A4(_05363_ ), .ZN(_06250_ ) );
BUF_X2 _14242_ ( .A(_05473_ ), .Z(_06251_ ) );
BUF_X2 _14243_ ( .A(_05603_ ), .Z(_06252_ ) );
OAI21_X1 _14244_ ( .A(_05361_ ), .B1(_06251_ ), .B2(_06252_ ), .ZN(_06253_ ) );
OAI211_X1 _14245_ ( .A(_06238_ ), .B(_06248_ ), .C1(_06250_ ), .C2(_06253_ ), .ZN(_06254_ ) );
INV_X1 _14246_ ( .A(_06254_ ), .ZN(_06255_ ) );
OAI21_X1 _14247_ ( .A(_06223_ ), .B1(_06245_ ), .B2(_06255_ ), .ZN(_06256_ ) );
MUX2_X1 _14248_ ( .A(_05934_ ), .B(_04487_ ), .S(_06219_ ), .Z(_06257_ ) );
OAI21_X1 _14249_ ( .A(_06256_ ), .B1(_06226_ ), .B2(_06257_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ) );
CLKBUF_X2 _14250_ ( .A(_05463_ ), .Z(_06258_ ) );
OR3_X1 _14251_ ( .A1(_06258_ ), .A2(\EX_LS_result_csreg_mem [19] ), .A3(_05603_ ), .ZN(_06259_ ) );
INV_X1 _14252_ ( .A(_05384_ ), .ZN(_06260_ ) );
NAND4_X1 _14253_ ( .A1(_06260_ ), .A2(_05414_ ), .A3(_05379_ ), .A4(_05381_ ), .ZN(_06261_ ) );
OAI21_X1 _14254_ ( .A(_05380_ ), .B1(_06246_ ), .B2(_06247_ ), .ZN(_06262_ ) );
OAI211_X1 _14255_ ( .A(_06259_ ), .B(_06237_ ), .C1(_06261_ ), .C2(_06262_ ), .ZN(_06263_ ) );
INV_X1 _14256_ ( .A(_06263_ ), .ZN(_06264_ ) );
AOI22_X1 _14257_ ( .A1(_05390_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_02371_ ), .ZN(_06265_ ) );
NAND3_X1 _14258_ ( .A1(_02349_ ), .A2(_02369_ ), .A3(_05851_ ), .ZN(_06266_ ) );
AOI211_X1 _14259_ ( .A(_06213_ ), .B(_06264_ ), .C1(_06265_ ), .C2(_06266_ ), .ZN(_06267_ ) );
MUX2_X1 _14260_ ( .A(_05399_ ), .B(_04405_ ), .S(_06219_ ), .Z(_06268_ ) );
AOI21_X1 _14261_ ( .A(_06267_ ), .B1(_06214_ ), .B2(_06268_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ) );
OR3_X1 _14262_ ( .A1(_06246_ ), .A2(\EX_LS_result_csreg_mem [18] ), .A3(_06247_ ), .ZN(_06269_ ) );
NAND4_X1 _14263_ ( .A1(_05409_ ), .A2(_05413_ ), .A3(_05411_ ), .A4(_05414_ ), .ZN(_06270_ ) );
OAI21_X1 _14264_ ( .A(_05410_ ), .B1(_06251_ ), .B2(_06252_ ), .ZN(_06271_ ) );
OAI211_X1 _14265_ ( .A(_06269_ ), .B(_06238_ ), .C1(_06270_ ), .C2(_06271_ ), .ZN(_06272_ ) );
OAI22_X1 _14266_ ( .A1(_05419_ ), .A2(_06234_ ), .B1(_05929_ ), .B2(\ID_EX_imm [18] ), .ZN(_06273_ ) );
AND3_X1 _14267_ ( .A1(_02324_ ), .A2(_05929_ ), .A3(_02345_ ), .ZN(_06274_ ) );
OAI211_X1 _14268_ ( .A(_06222_ ), .B(_06272_ ), .C1(_06273_ ), .C2(_06274_ ), .ZN(_06275_ ) );
NAND4_X1 _14269_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06276_ ) );
BUF_X4 _14270_ ( .A(_06217_ ), .Z(_06277_ ) );
OAI211_X1 _14271_ ( .A(_06221_ ), .B(_06276_ ), .C1(_04381_ ), .C2(_06277_ ), .ZN(_06278_ ) );
AND2_X1 _14272_ ( .A1(_06275_ ), .A2(_06278_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ) );
OR3_X1 _14273_ ( .A1(_06246_ ), .A2(\EX_LS_result_csreg_mem [17] ), .A3(_06247_ ), .ZN(_06279_ ) );
NAND4_X1 _14274_ ( .A1(_05444_ ), .A2(_05437_ ), .A3(_05438_ ), .A4(_05441_ ), .ZN(_06280_ ) );
OAI21_X1 _14275_ ( .A(_05440_ ), .B1(_06251_ ), .B2(_06252_ ), .ZN(_06281_ ) );
OAI211_X1 _14276_ ( .A(_06238_ ), .B(_06279_ ), .C1(_06280_ ), .C2(_06281_ ), .ZN(_06282_ ) );
OAI22_X1 _14277_ ( .A1(_05448_ ), .A2(_06234_ ), .B1(_05929_ ), .B2(\ID_EX_imm [17] ), .ZN(_06283_ ) );
AND3_X1 _14278_ ( .A1(_02374_ ), .A2(_05929_ ), .A3(_02393_ ), .ZN(_06284_ ) );
OAI211_X1 _14279_ ( .A(_06222_ ), .B(_06282_ ), .C1(_06283_ ), .C2(_06284_ ), .ZN(_06285_ ) );
NAND4_X1 _14280_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06286_ ) );
OAI211_X1 _14281_ ( .A(_06213_ ), .B(_06286_ ), .C1(_04429_ ), .C2(_06277_ ), .ZN(_06287_ ) );
AND2_X1 _14282_ ( .A1(_06285_ ), .A2(_06287_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ) );
BUF_X4 _14283_ ( .A(_06222_ ), .Z(_06288_ ) );
OAI22_X1 _14284_ ( .A1(_05476_ ), .A2(_04769_ ), .B1(_05850_ ), .B2(\ID_EX_imm [16] ), .ZN(_06289_ ) );
AOI21_X1 _14285_ ( .A(_06289_ ), .B1(_05930_ ), .B2(_04432_ ), .ZN(_06290_ ) );
INV_X1 _14286_ ( .A(_05475_ ), .ZN(_06291_ ) );
OAI211_X1 _14287_ ( .A(_06238_ ), .B(_06291_ ), .C1(_05467_ ), .C2(_05471_ ), .ZN(_06292_ ) );
INV_X1 _14288_ ( .A(_06292_ ), .ZN(_06293_ ) );
OAI21_X1 _14289_ ( .A(_06288_ ), .B1(_06290_ ), .B2(_06293_ ), .ZN(_06294_ ) );
MUX2_X1 _14290_ ( .A(_05453_ ), .B(_04459_ ), .S(_06219_ ), .Z(_06295_ ) );
OAI21_X1 _14291_ ( .A(_06294_ ), .B1(_06226_ ), .B2(_06295_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ) );
OR3_X1 _14292_ ( .A1(_06246_ ), .A2(\EX_LS_result_csreg_mem [15] ), .A3(_06247_ ), .ZN(_06296_ ) );
INV_X1 _14293_ ( .A(_05494_ ), .ZN(_06297_ ) );
NAND4_X1 _14294_ ( .A1(_06297_ ), .A2(_05414_ ), .A3(_05490_ ), .A4(_05492_ ), .ZN(_06298_ ) );
OAI21_X1 _14295_ ( .A(_05491_ ), .B1(_06251_ ), .B2(_06252_ ), .ZN(_06299_ ) );
OAI211_X1 _14296_ ( .A(_06238_ ), .B(_06296_ ), .C1(_06298_ ), .C2(_06299_ ), .ZN(_06300_ ) );
INV_X1 _14297_ ( .A(_06300_ ), .ZN(_06301_ ) );
AOI22_X1 _14298_ ( .A1(_05500_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_02695_ ), .ZN(_06302_ ) );
NAND3_X1 _14299_ ( .A1(_02674_ ), .A2(_02693_ ), .A3(_05930_ ), .ZN(_06303_ ) );
AOI211_X1 _14300_ ( .A(_06213_ ), .B(_06301_ ), .C1(_06302_ ), .C2(_06303_ ), .ZN(_06304_ ) );
AOI21_X1 _14301_ ( .A(_06217_ ), .B1(_04111_ ), .B2(_04131_ ), .ZN(_06305_ ) );
AOI211_X1 _14302_ ( .A(_06222_ ), .B(_06305_ ), .C1(\ID_EX_pc [15] ), .C2(_06277_ ), .ZN(_06306_ ) );
NOR2_X1 _14303_ ( .A1(_06304_ ), .A2(_06306_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ) );
OAI22_X1 _14304_ ( .A1(_05519_ ), .A2(_04769_ ), .B1(_05850_ ), .B2(\ID_EX_imm [14] ), .ZN(_06307_ ) );
AOI21_X1 _14305_ ( .A(_06307_ ), .B1(_05930_ ), .B2(_04134_ ), .ZN(_06308_ ) );
INV_X1 _14306_ ( .A(_05518_ ), .ZN(_06309_ ) );
OAI211_X1 _14307_ ( .A(_06238_ ), .B(_06309_ ), .C1(_05513_ ), .C2(_05516_ ), .ZN(_06310_ ) );
INV_X1 _14308_ ( .A(_06310_ ), .ZN(_06311_ ) );
OAI21_X1 _14309_ ( .A(_06288_ ), .B1(_06308_ ), .B2(_06311_ ), .ZN(_06312_ ) );
MUX2_X1 _14310_ ( .A(_05505_ ), .B(_04164_ ), .S(_06219_ ), .Z(_06313_ ) );
OAI21_X1 _14311_ ( .A(_06312_ ), .B1(_06226_ ), .B2(_06313_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ) );
OAI22_X1 _14312_ ( .A1(_05542_ ), .A2(_04769_ ), .B1(_05850_ ), .B2(\ID_EX_imm [13] ), .ZN(_06314_ ) );
INV_X1 _14313_ ( .A(_04075_ ), .ZN(_06315_ ) );
AOI21_X1 _14314_ ( .A(_06314_ ), .B1(_05929_ ), .B2(_06315_ ), .ZN(_06316_ ) );
BUF_X2 _14315_ ( .A(_06212_ ), .Z(_06317_ ) );
NAND3_X1 _14316_ ( .A1(_05539_ ), .A2(_06237_ ), .A3(_05541_ ), .ZN(_06318_ ) );
INV_X1 _14317_ ( .A(_06318_ ), .ZN(_06319_ ) );
OR3_X1 _14318_ ( .A1(_06316_ ), .A2(_06317_ ), .A3(_06319_ ), .ZN(_06320_ ) );
NAND4_X1 _14319_ ( .A1(\ID_EX_pc [13] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06321_ ) );
OAI211_X1 _14320_ ( .A(_06213_ ), .B(_06321_ ), .C1(_04074_ ), .C2(_06277_ ), .ZN(_06322_ ) );
AND2_X1 _14321_ ( .A1(_06320_ ), .A2(_06322_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ) );
OAI22_X1 _14322_ ( .A1(_05560_ ), .A2(_04769_ ), .B1(_05850_ ), .B2(\ID_EX_imm [12] ), .ZN(_06323_ ) );
AOI21_X1 _14323_ ( .A(_06323_ ), .B1(_05930_ ), .B2(_04079_ ), .ZN(_06324_ ) );
NOR3_X1 _14324_ ( .A1(_06251_ ), .A2(_06247_ ), .A3(\EX_LS_result_csreg_mem [12] ), .ZN(_06325_ ) );
INV_X1 _14325_ ( .A(_06325_ ), .ZN(_06326_ ) );
OAI211_X1 _14326_ ( .A(_05551_ ), .B(_05552_ ), .C1(_06251_ ), .C2(_06252_ ), .ZN(_06327_ ) );
NAND3_X1 _14327_ ( .A1(_05444_ ), .A2(_05554_ ), .A3(_05555_ ), .ZN(_06328_ ) );
OAI211_X1 _14328_ ( .A(_06238_ ), .B(_06326_ ), .C1(_06327_ ), .C2(_06328_ ), .ZN(_06329_ ) );
INV_X1 _14329_ ( .A(_06329_ ), .ZN(_06330_ ) );
OAI21_X1 _14330_ ( .A(_06288_ ), .B1(_06324_ ), .B2(_06330_ ), .ZN(_06331_ ) );
MUX2_X1 _14331_ ( .A(_05546_ ), .B(_04106_ ), .S(_06219_ ), .Z(_06332_ ) );
OAI21_X1 _14332_ ( .A(_06331_ ), .B1(_06226_ ), .B2(_06332_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ) );
BUF_X4 _14333_ ( .A(_06211_ ), .Z(_06333_ ) );
OR3_X1 _14334_ ( .A1(_06258_ ), .A2(\EX_LS_result_csreg_mem [30] ), .A3(_05474_ ), .ZN(_06334_ ) );
AND2_X1 _14335_ ( .A1(_05243_ ), .A2(_05254_ ), .ZN(_06335_ ) );
INV_X1 _14336_ ( .A(_05263_ ), .ZN(_06336_ ) );
NAND2_X1 _14337_ ( .A1(_06335_ ), .A2(_06336_ ), .ZN(_06337_ ) );
OAI211_X1 _14338_ ( .A(_05258_ ), .B(_05719_ ), .C1(_06246_ ), .C2(_06247_ ), .ZN(_06338_ ) );
OAI21_X1 _14339_ ( .A(_06334_ ), .B1(_06337_ ), .B2(_06338_ ), .ZN(_06339_ ) );
AOI22_X1 _14340_ ( .A1(_06339_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_02964_ ), .ZN(_06340_ ) );
INV_X1 _14341_ ( .A(_02963_ ), .ZN(_06341_ ) );
OAI211_X1 _14342_ ( .A(_06333_ ), .B(_06340_ ), .C1(_06341_ ), .C2(fanout_net_5 ), .ZN(_06342_ ) );
INV_X1 _14343_ ( .A(_06237_ ), .ZN(_06343_ ) );
OR3_X1 _14344_ ( .A1(_06339_ ), .A2(_06343_ ), .A3(_06317_ ), .ZN(_06344_ ) );
MUX2_X1 _14345_ ( .A(_03911_ ), .B(_04657_ ), .S(_06218_ ), .Z(_06345_ ) );
OAI211_X1 _14346_ ( .A(_06342_ ), .B(_06344_ ), .C1(_06226_ ), .C2(_06345_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ) );
OAI211_X1 _14347_ ( .A(_05576_ ), .B(_05577_ ), .C1(_05473_ ), .C2(_05603_ ), .ZN(_06346_ ) );
NAND3_X1 _14348_ ( .A1(_05444_ ), .A2(_05574_ ), .A3(_05575_ ), .ZN(_06347_ ) );
NOR2_X1 _14349_ ( .A1(_06346_ ), .A2(_06347_ ), .ZN(_06348_ ) );
NOR3_X1 _14350_ ( .A1(_06258_ ), .A2(_05474_ ), .A3(\EX_LS_result_csreg_mem [11] ), .ZN(_06349_ ) );
NOR2_X1 _14351_ ( .A1(_06348_ ), .A2(_06349_ ), .ZN(_06350_ ) );
OAI22_X1 _14352_ ( .A1(_06350_ ), .A2(_04769_ ), .B1(_05850_ ), .B2(\ID_EX_imm [11] ), .ZN(_06351_ ) );
AOI21_X1 _14353_ ( .A(_06351_ ), .B1(_05930_ ), .B2(_03916_ ), .ZN(_06352_ ) );
INV_X1 _14354_ ( .A(_06349_ ), .ZN(_06353_ ) );
OAI211_X1 _14355_ ( .A(_06238_ ), .B(_06353_ ), .C1(_06346_ ), .C2(_06347_ ), .ZN(_06354_ ) );
INV_X1 _14356_ ( .A(_06354_ ), .ZN(_06355_ ) );
OAI21_X1 _14357_ ( .A(_06288_ ), .B1(_06352_ ), .B2(_06355_ ), .ZN(_06356_ ) );
MUX2_X1 _14358_ ( .A(_05305_ ), .B(_03964_ ), .S(_06219_ ), .Z(_06357_ ) );
OAI21_X1 _14359_ ( .A(_06356_ ), .B1(_06226_ ), .B2(_06357_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ) );
OR3_X1 _14360_ ( .A1(_06258_ ), .A2(\EX_LS_result_csreg_mem [10] ), .A3(_05603_ ), .ZN(_06358_ ) );
AND2_X1 _14361_ ( .A1(_05616_ ), .A2(_05414_ ), .ZN(_06359_ ) );
INV_X1 _14362_ ( .A(_05612_ ), .ZN(_06360_ ) );
NAND3_X1 _14363_ ( .A1(_06359_ ), .A2(_06360_ ), .A3(_05615_ ), .ZN(_06361_ ) );
OAI21_X1 _14364_ ( .A(_05614_ ), .B1(_06246_ ), .B2(_06247_ ), .ZN(_06362_ ) );
OAI211_X1 _14365_ ( .A(_06358_ ), .B(_06237_ ), .C1(_06361_ ), .C2(_06362_ ), .ZN(_06363_ ) );
INV_X1 _14366_ ( .A(_06363_ ), .ZN(_06364_ ) );
AOI22_X1 _14367_ ( .A1(_05620_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_02743_ ), .ZN(_06365_ ) );
NAND3_X1 _14368_ ( .A1(_02721_ ), .A2(_02740_ ), .A3(_05851_ ), .ZN(_06366_ ) );
AOI211_X1 _14369_ ( .A(_06213_ ), .B(_06364_ ), .C1(_06365_ ), .C2(_06366_ ), .ZN(_06367_ ) );
MUX2_X1 _14370_ ( .A(_05306_ ), .B(_03991_ ), .S(_06219_ ), .Z(_06368_ ) );
AOI21_X1 _14371_ ( .A(_06367_ ), .B1(_06214_ ), .B2(_06368_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ) );
NOR2_X1 _14372_ ( .A1(_05643_ ), .A2(_05530_ ), .ZN(_06369_ ) );
INV_X1 _14373_ ( .A(_05639_ ), .ZN(_06370_ ) );
AND2_X1 _14374_ ( .A1(_05642_ ), .A2(_05414_ ), .ZN(_06371_ ) );
NAND4_X1 _14375_ ( .A1(_06369_ ), .A2(_06370_ ), .A3(_05641_ ), .A4(_06371_ ), .ZN(_06372_ ) );
OR3_X1 _14376_ ( .A1(_06258_ ), .A2(\EX_LS_result_csreg_mem [9] ), .A3(_05474_ ), .ZN(_06373_ ) );
NAND2_X1 _14377_ ( .A1(_06372_ ), .A2(_06373_ ), .ZN(_06374_ ) );
AOI22_X1 _14378_ ( .A1(_06374_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_02813_ ), .ZN(_06375_ ) );
OAI211_X1 _14379_ ( .A(_06375_ ), .B(_06333_ ), .C1(fanout_net_5 ), .C2(_02812_ ), .ZN(_06376_ ) );
BUF_X4 _14380_ ( .A(_06237_ ), .Z(_06377_ ) );
NAND4_X1 _14381_ ( .A1(_06372_ ), .A2(_06377_ ), .A3(_06373_ ), .A4(_06225_ ), .ZN(_06378_ ) );
MUX2_X1 _14382_ ( .A(_05630_ ), .B(_04047_ ), .S(_06218_ ), .Z(_06379_ ) );
OAI211_X1 _14383_ ( .A(_06376_ ), .B(_06378_ ), .C1(_06226_ ), .C2(_06379_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ) );
OR3_X1 _14384_ ( .A1(_05463_ ), .A2(\EX_LS_result_csreg_mem [8] ), .A3(_05466_ ), .ZN(_06380_ ) );
OAI211_X1 _14385_ ( .A(_05655_ ), .B(_05657_ ), .C1(_05473_ ), .C2(_05603_ ), .ZN(_06381_ ) );
NAND3_X1 _14386_ ( .A1(_05444_ ), .A2(_05656_ ), .A3(_05658_ ), .ZN(_06382_ ) );
OAI21_X1 _14387_ ( .A(_06380_ ), .B1(_06381_ ), .B2(_06382_ ), .ZN(_06383_ ) );
AOI221_X4 _14388_ ( .A(_06212_ ), .B1(fanout_net_5 ), .B2(_02790_ ), .C1(_06383_ ), .C2(\ID_EX_typ [2] ), .ZN(_06384_ ) );
OAI21_X1 _14389_ ( .A(_06384_ ), .B1(fanout_net_5 ), .B2(_02789_ ), .ZN(_06385_ ) );
AND2_X1 _14390_ ( .A1(_05655_ ), .A2(_05657_ ), .ZN(_06386_ ) );
AND2_X1 _14391_ ( .A1(_05656_ ), .A2(_05658_ ), .ZN(_06387_ ) );
NAND4_X1 _14392_ ( .A1(_05293_ ), .A2(_06386_ ), .A3(_06387_ ), .A4(_05444_ ), .ZN(_06388_ ) );
INV_X1 _14393_ ( .A(_05654_ ), .ZN(_06389_ ) );
NAND4_X1 _14394_ ( .A1(_06388_ ), .A2(_06377_ ), .A3(_06389_ ), .A4(_06225_ ), .ZN(_06390_ ) );
NOR2_X1 _14395_ ( .A1(_04021_ ), .A2(_06217_ ), .ZN(_06391_ ) );
AOI21_X1 _14396_ ( .A(_06391_ ), .B1(\ID_EX_pc [8] ), .B2(_06277_ ), .ZN(_06392_ ) );
BUF_X4 _14397_ ( .A(_06222_ ), .Z(_06393_ ) );
OAI211_X1 _14398_ ( .A(_06385_ ), .B(_06390_ ), .C1(_06392_ ), .C2(_06393_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ) );
NOR3_X1 _14399_ ( .A1(_06251_ ), .A2(_06252_ ), .A3(\EX_LS_result_csreg_mem [7] ), .ZN(_06394_ ) );
AND4_X1 _14400_ ( .A1(_05670_ ), .A2(_05671_ ), .A3(_05672_ ), .A4(_05673_ ), .ZN(_06395_ ) );
AOI21_X1 _14401_ ( .A(_06394_ ), .B1(_06395_ ), .B2(_05531_ ), .ZN(_06396_ ) );
AOI21_X1 _14402_ ( .A(fanout_net_5 ), .B1(_02523_ ), .B2(_02542_ ), .ZN(_06397_ ) );
AND2_X1 _14403_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [7] ), .ZN(_06398_ ) );
OAI221_X1 _14404_ ( .A(_06225_ ), .B1(_06234_ ), .B2(_06396_ ), .C1(_06397_ ), .C2(_06398_ ), .ZN(_06399_ ) );
AND2_X1 _14405_ ( .A1(_05670_ ), .A2(_05673_ ), .ZN(_06400_ ) );
AND2_X1 _14406_ ( .A1(_05671_ ), .A2(_05672_ ), .ZN(_06401_ ) );
NAND3_X1 _14407_ ( .A1(_05531_ ), .A2(_06400_ ), .A3(_06401_ ), .ZN(_06402_ ) );
OR3_X1 _14408_ ( .A1(_06251_ ), .A2(\EX_LS_result_csreg_mem [7] ), .A3(_06252_ ), .ZN(_06403_ ) );
NAND4_X1 _14409_ ( .A1(_06402_ ), .A2(_06377_ ), .A3(_06403_ ), .A4(_06225_ ), .ZN(_06404_ ) );
MUX2_X1 _14410_ ( .A(_05676_ ), .B(_04212_ ), .S(_06218_ ), .Z(_06405_ ) );
OAI211_X1 _14411_ ( .A(_06399_ ), .B(_06404_ ), .C1(_06226_ ), .C2(_06405_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ) );
OAI22_X1 _14412_ ( .A1(_05705_ ), .A2(_04769_ ), .B1(_05850_ ), .B2(\ID_EX_imm [6] ), .ZN(_06406_ ) );
AOI21_X1 _14413_ ( .A(_06406_ ), .B1(_05929_ ), .B2(_04189_ ), .ZN(_06407_ ) );
NAND3_X1 _14414_ ( .A1(_05702_ ), .A2(_06237_ ), .A3(_05704_ ), .ZN(_06408_ ) );
INV_X1 _14415_ ( .A(_06408_ ), .ZN(_06409_ ) );
OR3_X1 _14416_ ( .A1(_06407_ ), .A2(_06317_ ), .A3(_06409_ ), .ZN(_06410_ ) );
NAND4_X1 _14417_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06411_ ) );
OAI211_X1 _14418_ ( .A(_06213_ ), .B(_06411_ ), .C1(_04188_ ), .C2(_06277_ ), .ZN(_06412_ ) );
AND2_X1 _14419_ ( .A1(_06410_ ), .A2(_06412_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ) );
OAI22_X1 _14420_ ( .A1(_05726_ ), .A2(_06234_ ), .B1(_05929_ ), .B2(\ID_EX_imm [5] ), .ZN(_06413_ ) );
AOI21_X1 _14421_ ( .A(_06413_ ), .B1(_05932_ ), .B2(_04901_ ), .ZN(_06414_ ) );
NOR3_X1 _14422_ ( .A1(_06251_ ), .A2(_06252_ ), .A3(\EX_LS_result_csreg_mem [5] ), .ZN(_06415_ ) );
INV_X1 _14423_ ( .A(_06415_ ), .ZN(_06416_ ) );
NAND4_X1 _14424_ ( .A1(_05716_ ), .A2(_05720_ ), .A3(_05721_ ), .A4(_05719_ ), .ZN(_06417_ ) );
OAI21_X1 _14425_ ( .A(_05717_ ), .B1(_06251_ ), .B2(_06252_ ), .ZN(_06418_ ) );
OAI211_X1 _14426_ ( .A(_06416_ ), .B(_06377_ ), .C1(_06417_ ), .C2(_06418_ ), .ZN(_06419_ ) );
INV_X1 _14427_ ( .A(_06419_ ), .ZN(_06420_ ) );
OAI21_X1 _14428_ ( .A(_06223_ ), .B1(_06414_ ), .B2(_06420_ ), .ZN(_06421_ ) );
BUF_X4 _14429_ ( .A(_06213_ ), .Z(_06422_ ) );
NAND3_X1 _14430_ ( .A1(_03354_ ), .A2(_05709_ ), .A3(\ID_EX_typ [7] ), .ZN(_06423_ ) );
OAI211_X1 _14431_ ( .A(_06422_ ), .B(_06423_ ), .C1(_04234_ ), .C2(_06277_ ), .ZN(_06424_ ) );
NAND2_X1 _14432_ ( .A1(_06421_ ), .A2(_06424_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ) );
BUF_X4 _14433_ ( .A(_06218_ ), .Z(_06425_ ) );
NAND3_X1 _14434_ ( .A1(_04259_ ), .A2(_04279_ ), .A3(_06425_ ), .ZN(_06426_ ) );
OAI211_X1 _14435_ ( .A(_06426_ ), .B(_06221_ ), .C1(\ID_EX_pc [4] ), .C2(_06425_ ), .ZN(_06427_ ) );
INV_X1 _14436_ ( .A(_05740_ ), .ZN(_06428_ ) );
INV_X1 _14437_ ( .A(_05737_ ), .ZN(_06429_ ) );
INV_X1 _14438_ ( .A(_05695_ ), .ZN(_06430_ ) );
OAI211_X1 _14439_ ( .A(_06237_ ), .B(_06428_ ), .C1(_06429_ ), .C2(_06430_ ), .ZN(_06431_ ) );
OAI21_X1 _14440_ ( .A(_06431_ ), .B1(_05930_ ), .B2(_02612_ ), .ZN(_06432_ ) );
AOI21_X1 _14441_ ( .A(_06432_ ), .B1(_05932_ ), .B2(_02611_ ), .ZN(_06433_ ) );
BUF_X4 _14442_ ( .A(_06222_ ), .Z(_06434_ ) );
OAI21_X1 _14443_ ( .A(_06434_ ), .B1(_05741_ ), .B2(_06234_ ), .ZN(_06435_ ) );
OAI21_X1 _14444_ ( .A(_06427_ ), .B1(_06433_ ), .B2(_06435_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ) );
NAND3_X1 _14445_ ( .A1(_02495_ ), .A2(_05930_ ), .A3(_02515_ ), .ZN(_06436_ ) );
OR3_X1 _14446_ ( .A1(_06258_ ), .A2(\EX_LS_result_csreg_mem [3] ), .A3(_05474_ ), .ZN(_06437_ ) );
OAI211_X1 _14447_ ( .A(_05759_ ), .B(_05760_ ), .C1(_06246_ ), .C2(_06252_ ), .ZN(_06438_ ) );
NAND3_X1 _14448_ ( .A1(_05758_ ), .A2(_05719_ ), .A3(_05757_ ), .ZN(_06439_ ) );
OAI21_X1 _14449_ ( .A(_06437_ ), .B1(_06438_ ), .B2(_06439_ ), .ZN(_06440_ ) );
NAND2_X1 _14450_ ( .A1(_06440_ ), .A2(\ID_EX_typ [2] ), .ZN(_06441_ ) );
OR2_X1 _14451_ ( .A1(_05929_ ), .A2(\ID_EX_imm [3] ), .ZN(_06442_ ) );
NAND4_X1 _14452_ ( .A1(_06436_ ), .A2(_06333_ ), .A3(_06441_ ), .A4(_06442_ ), .ZN(_06443_ ) );
OR3_X1 _14453_ ( .A1(_06440_ ), .A2(_06343_ ), .A3(_06317_ ), .ZN(_06444_ ) );
AND3_X1 _14454_ ( .A1(_03354_ ), .A2(\ID_EX_pc [3] ), .A3(\ID_EX_typ [7] ), .ZN(_06445_ ) );
AOI21_X1 _14455_ ( .A(_06445_ ), .B1(_04328_ ), .B2(_06425_ ), .ZN(_06446_ ) );
OAI211_X1 _14456_ ( .A(_06443_ ), .B(_06444_ ), .C1(_06446_ ), .C2(_06393_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ) );
NOR2_X1 _14457_ ( .A1(_05775_ ), .A2(_05530_ ), .ZN(_06447_ ) );
NOR2_X1 _14458_ ( .A1(_05359_ ), .A2(_05776_ ), .ZN(_06448_ ) );
AND2_X1 _14459_ ( .A1(_05772_ ), .A2(_05773_ ), .ZN(_06449_ ) );
NAND3_X1 _14460_ ( .A1(_06447_ ), .A2(_06448_ ), .A3(_06449_ ), .ZN(_06450_ ) );
OR3_X1 _14461_ ( .A1(_06258_ ), .A2(\EX_LS_result_csreg_mem [2] ), .A3(_05474_ ), .ZN(_06451_ ) );
NAND2_X1 _14462_ ( .A1(_06450_ ), .A2(_06451_ ), .ZN(_06452_ ) );
AOI22_X1 _14463_ ( .A1(_06452_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_02442_ ), .ZN(_06453_ ) );
OAI211_X1 _14464_ ( .A(_06453_ ), .B(_06333_ ), .C1(_02441_ ), .C2(fanout_net_5 ), .ZN(_06454_ ) );
NAND4_X1 _14465_ ( .A1(_06450_ ), .A2(_06377_ ), .A3(_06451_ ), .A4(_06225_ ), .ZN(_06455_ ) );
AOI21_X1 _14466_ ( .A(_06217_ ), .B1(_04303_ ), .B2(_04301_ ), .ZN(_06456_ ) );
AOI21_X1 _14467_ ( .A(_06456_ ), .B1(\ID_EX_pc [2] ), .B2(_06277_ ), .ZN(_06457_ ) );
OAI211_X1 _14468_ ( .A(_06454_ ), .B(_06455_ ), .C1(_06393_ ), .C2(_06457_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ) );
OR3_X1 _14469_ ( .A1(_06258_ ), .A2(_05474_ ), .A3(\EX_LS_result_csreg_mem [29] ), .ZN(_06458_ ) );
NAND4_X1 _14470_ ( .A1(_05329_ ), .A2(_05340_ ), .A3(_05719_ ), .A4(_05335_ ), .ZN(_06459_ ) );
OAI21_X1 _14471_ ( .A(_05332_ ), .B1(_06246_ ), .B2(_06247_ ), .ZN(_06460_ ) );
OAI21_X1 _14472_ ( .A(_06458_ ), .B1(_06459_ ), .B2(_06460_ ), .ZN(_06461_ ) );
AOI22_X1 _14473_ ( .A1(_06461_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_5 ), .B2(_02935_ ), .ZN(_06462_ ) );
OAI211_X1 _14474_ ( .A(_06462_ ), .B(_06333_ ), .C1(_02934_ ), .C2(fanout_net_5 ), .ZN(_06463_ ) );
OR3_X1 _14475_ ( .A1(_06461_ ), .A2(_06343_ ), .A3(_06317_ ), .ZN(_06464_ ) );
AND3_X1 _14476_ ( .A1(_03354_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_typ [7] ), .ZN(_06465_ ) );
AOI21_X1 _14477_ ( .A(_06465_ ), .B1(_04585_ ), .B2(_06425_ ), .ZN(_06466_ ) );
OAI211_X1 _14478_ ( .A(_06463_ ), .B(_06464_ ), .C1(_06466_ ), .C2(_06393_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ) );
OR3_X1 _14479_ ( .A1(_05473_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_05603_ ), .ZN(_06467_ ) );
NAND4_X1 _14480_ ( .A1(_05787_ ), .A2(_05788_ ), .A3(_05786_ ), .A4(_05789_ ), .ZN(_06468_ ) );
OAI21_X1 _14481_ ( .A(_06467_ ), .B1(_06468_ ), .B2(_05530_ ), .ZN(_06469_ ) );
AOI22_X1 _14482_ ( .A1(_04236_ ), .A2(_05851_ ), .B1(\ID_EX_typ [2] ), .B2(_06469_ ), .ZN(_06470_ ) );
OAI211_X1 _14483_ ( .A(_06470_ ), .B(_06333_ ), .C1(_05932_ ), .C2(\ID_EX_imm [1] ), .ZN(_06471_ ) );
AND2_X1 _14484_ ( .A1(_05786_ ), .A2(_05789_ ), .ZN(_06472_ ) );
AND2_X1 _14485_ ( .A1(_05787_ ), .A2(_05788_ ), .ZN(_06473_ ) );
NAND3_X1 _14486_ ( .A1(_05531_ ), .A2(_06472_ ), .A3(_06473_ ), .ZN(_06474_ ) );
NAND4_X1 _14487_ ( .A1(_06474_ ), .A2(_06377_ ), .A3(_06467_ ), .A4(_06225_ ), .ZN(_06475_ ) );
MUX2_X1 _14488_ ( .A(_05795_ ), .B(_04256_ ), .S(_06218_ ), .Z(_06476_ ) );
OAI211_X1 _14489_ ( .A(_06471_ ), .B(_06475_ ), .C1(_06393_ ), .C2(_06476_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ) );
AOI21_X1 _14490_ ( .A(_06343_ ), .B1(_05827_ ), .B2(_05828_ ), .ZN(_06477_ ) );
AOI21_X1 _14491_ ( .A(_06477_ ), .B1(\ID_EX_typ [0] ), .B2(\ID_EX_imm [0] ), .ZN(_06478_ ) );
INV_X1 _14492_ ( .A(_04331_ ), .ZN(_06479_ ) );
OAI21_X1 _14493_ ( .A(_06478_ ), .B1(_06479_ ), .B2(\ID_EX_typ [0] ), .ZN(_06480_ ) );
OAI211_X1 _14494_ ( .A(_06480_ ), .B(_06223_ ), .C1(_06234_ ), .C2(_05830_ ), .ZN(_06481_ ) );
NAND3_X1 _14495_ ( .A1(_04351_ ), .A2(_04352_ ), .A3(_06425_ ), .ZN(_06482_ ) );
OAI211_X1 _14496_ ( .A(_06482_ ), .B(_06422_ ), .C1(\ID_EX_pc [0] ), .C2(_06425_ ), .ZN(_06483_ ) );
NAND2_X1 _14497_ ( .A1(_06481_ ), .A2(_06483_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ) );
AOI22_X1 _14498_ ( .A1(_04778_ ), .A2(_05851_ ), .B1(\ID_EX_typ [2] ), .B2(_05605_ ), .ZN(_06484_ ) );
OAI211_X1 _14499_ ( .A(_06484_ ), .B(_06333_ ), .C1(_05932_ ), .C2(\ID_EX_imm [28] ), .ZN(_06485_ ) );
NAND4_X1 _14500_ ( .A1(_05602_ ), .A2(_06377_ ), .A3(_05604_ ), .A4(_06222_ ), .ZN(_06486_ ) );
AND3_X1 _14501_ ( .A1(_03354_ ), .A2(\ID_EX_pc [28] ), .A3(\ID_EX_typ [7] ), .ZN(_06487_ ) );
AOI21_X1 _14502_ ( .A(_06487_ ), .B1(_04609_ ), .B2(_06425_ ), .ZN(_06488_ ) );
OAI211_X1 _14503_ ( .A(_06485_ ), .B(_06486_ ), .C1(_06393_ ), .C2(_06488_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ) );
AOI22_X1 _14504_ ( .A1(_05817_ ), .A2(_06238_ ), .B1(\ID_EX_typ [0] ), .B2(\ID_EX_imm [27] ), .ZN(_06489_ ) );
OAI21_X1 _14505_ ( .A(_06489_ ), .B1(\ID_EX_typ [0] ), .B2(_04708_ ), .ZN(_06490_ ) );
OAI211_X1 _14506_ ( .A(_06490_ ), .B(_06223_ ), .C1(_06234_ ), .C2(_05817_ ), .ZN(_06491_ ) );
NAND4_X1 _14507_ ( .A1(_05210_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06492_ ) );
OAI211_X1 _14508_ ( .A(_06422_ ), .B(_06492_ ), .C1(_04706_ ), .C2(_06277_ ), .ZN(_06493_ ) );
NAND2_X1 _14509_ ( .A1(_06491_ ), .A2(_06493_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ) );
OR3_X1 _14510_ ( .A1(_05473_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_05603_ ), .ZN(_06494_ ) );
NAND4_X1 _14511_ ( .A1(_05844_ ), .A2(_05845_ ), .A3(_05843_ ), .A4(_05846_ ), .ZN(_06495_ ) );
OAI21_X1 _14512_ ( .A(_06494_ ), .B1(_06495_ ), .B2(_05530_ ), .ZN(_06496_ ) );
AOI22_X1 _14513_ ( .A1(_04791_ ), .A2(_05851_ ), .B1(\ID_EX_typ [2] ), .B2(_06496_ ), .ZN(_06497_ ) );
OAI211_X1 _14514_ ( .A(_06497_ ), .B(_06333_ ), .C1(_05932_ ), .C2(\ID_EX_imm [26] ), .ZN(_06498_ ) );
AND2_X1 _14515_ ( .A1(_05843_ ), .A2(_05846_ ), .ZN(_06499_ ) );
AND2_X1 _14516_ ( .A1(_05844_ ), .A2(_05845_ ), .ZN(_06500_ ) );
NAND3_X1 _14517_ ( .A1(_05531_ ), .A2(_06499_ ), .A3(_06500_ ), .ZN(_06501_ ) );
NAND4_X1 _14518_ ( .A1(_06501_ ), .A2(_06377_ ), .A3(_06494_ ), .A4(_06222_ ), .ZN(_06502_ ) );
AND3_X1 _14519_ ( .A1(_03354_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_typ [7] ), .ZN(_06503_ ) );
AOI21_X1 _14520_ ( .A(_06503_ ), .B1(_04684_ ), .B2(_06425_ ), .ZN(_06504_ ) );
OAI211_X1 _14521_ ( .A(_06498_ ), .B(_06502_ ), .C1(_06504_ ), .C2(_06393_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ) );
OR3_X1 _14522_ ( .A1(_05473_ ), .A2(_05603_ ), .A3(\EX_LS_result_csreg_mem [25] ), .ZN(_06505_ ) );
NAND4_X1 _14523_ ( .A1(_05868_ ), .A2(_05869_ ), .A3(_05867_ ), .A4(_05870_ ), .ZN(_06506_ ) );
OAI21_X1 _14524_ ( .A(_06505_ ), .B1(_06506_ ), .B2(_05530_ ), .ZN(_06507_ ) );
AOI22_X1 _14525_ ( .A1(_02907_ ), .A2(_05851_ ), .B1(\ID_EX_typ [2] ), .B2(_06507_ ), .ZN(_06508_ ) );
OAI211_X1 _14526_ ( .A(_06508_ ), .B(_06225_ ), .C1(_05932_ ), .C2(\ID_EX_imm [25] ), .ZN(_06509_ ) );
OR3_X1 _14527_ ( .A1(_06507_ ), .A2(_06343_ ), .A3(_06317_ ), .ZN(_06510_ ) );
AND3_X1 _14528_ ( .A1(_03354_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_typ [7] ), .ZN(_06511_ ) );
AOI21_X1 _14529_ ( .A(_06511_ ), .B1(_04756_ ), .B2(_06425_ ), .ZN(_06512_ ) );
OAI211_X1 _14530_ ( .A(_06509_ ), .B(_06510_ ), .C1(_06512_ ), .C2(_06393_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ) );
OR4_X1 _14531_ ( .A1(\ID_EX_pc [24] ), .A2(_03341_ ), .A3(_03881_ ), .A4(_06210_ ), .ZN(_06513_ ) );
OAI211_X1 _14532_ ( .A(_06221_ ), .B(_06513_ ), .C1(_04733_ ), .C2(_06277_ ), .ZN(_06514_ ) );
INV_X1 _14533_ ( .A(_05889_ ), .ZN(_06515_ ) );
INV_X1 _14534_ ( .A(_05573_ ), .ZN(_06516_ ) );
INV_X1 _14535_ ( .A(_05886_ ), .ZN(_06517_ ) );
OAI211_X1 _14536_ ( .A(_06237_ ), .B(_06515_ ), .C1(_06516_ ), .C2(_06517_ ), .ZN(_06518_ ) );
OAI21_X1 _14537_ ( .A(_06518_ ), .B1(_05851_ ), .B2(_02877_ ), .ZN(_06519_ ) );
AOI21_X1 _14538_ ( .A(_06519_ ), .B1(_05932_ ), .B2(_02876_ ), .ZN(_06520_ ) );
OAI21_X1 _14539_ ( .A(_06434_ ), .B1(_05890_ ), .B2(_06234_ ), .ZN(_06521_ ) );
OAI21_X1 _14540_ ( .A(_06514_ ), .B1(_06520_ ), .B2(_06521_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ) );
OR3_X1 _14541_ ( .A1(_05473_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_05603_ ), .ZN(_06522_ ) );
NAND4_X1 _14542_ ( .A1(_05904_ ), .A2(_05905_ ), .A3(_05903_ ), .A4(_05906_ ), .ZN(_06523_ ) );
OAI21_X1 _14543_ ( .A(_06522_ ), .B1(_06523_ ), .B2(_05530_ ), .ZN(_06524_ ) );
AOI22_X1 _14544_ ( .A1(_04943_ ), .A2(_05851_ ), .B1(\ID_EX_typ [2] ), .B2(_06524_ ), .ZN(_06525_ ) );
OAI211_X1 _14545_ ( .A(_06525_ ), .B(_06434_ ), .C1(_05932_ ), .C2(\ID_EX_imm [23] ), .ZN(_06526_ ) );
AOI21_X1 _14546_ ( .A(_06217_ ), .B1(_04534_ ), .B2(_04535_ ), .ZN(_06527_ ) );
AND3_X1 _14547_ ( .A1(_03354_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_typ [7] ), .ZN(_06528_ ) );
OAI21_X1 _14548_ ( .A(_06422_ ), .B1(_06527_ ), .B2(_06528_ ), .ZN(_06529_ ) );
AND2_X1 _14549_ ( .A1(_05903_ ), .A2(_05906_ ), .ZN(_06530_ ) );
AND2_X1 _14550_ ( .A1(_05904_ ), .A2(_05905_ ), .ZN(_06531_ ) );
NAND3_X1 _14551_ ( .A1(_05531_ ), .A2(_06530_ ), .A3(_06531_ ), .ZN(_06532_ ) );
NAND4_X1 _14552_ ( .A1(_06532_ ), .A2(_06377_ ), .A3(_06522_ ), .A4(_06333_ ), .ZN(_06533_ ) );
NAND3_X1 _14553_ ( .A1(_06526_ ), .A2(_06529_ ), .A3(_06533_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ) );
OR3_X1 _14554_ ( .A1(_06258_ ), .A2(\EX_LS_result_csreg_mem [22] ), .A3(_05474_ ), .ZN(_06534_ ) );
NAND4_X1 _14555_ ( .A1(_05444_ ), .A2(_05921_ ), .A3(_05924_ ), .A4(_05922_ ), .ZN(_06535_ ) );
OAI21_X1 _14556_ ( .A(_05923_ ), .B1(_06246_ ), .B2(_06247_ ), .ZN(_06536_ ) );
OAI21_X1 _14557_ ( .A(_06534_ ), .B1(_06535_ ), .B2(_06536_ ), .ZN(_06537_ ) );
AOI22_X1 _14558_ ( .A1(_06537_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02271_ ), .ZN(_06538_ ) );
OAI211_X1 _14559_ ( .A(_06538_ ), .B(_06225_ ), .C1(\ID_EX_typ [0] ), .C2(_02270_ ), .ZN(_06539_ ) );
OR3_X1 _14560_ ( .A1(_06537_ ), .A2(_06343_ ), .A3(_06317_ ), .ZN(_06540_ ) );
MUX2_X1 _14561_ ( .A(_05912_ ), .B(_04561_ ), .S(_06219_ ), .Z(_06541_ ) );
OAI211_X1 _14562_ ( .A(_06539_ ), .B(_06540_ ), .C1(_06541_ ), .C2(_06223_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ) );
NOR3_X1 _14563_ ( .A1(_06258_ ), .A2(_05474_ ), .A3(\EX_LS_result_csreg_mem [31] ), .ZN(_06542_ ) );
INV_X1 _14564_ ( .A(_06542_ ), .ZN(_06543_ ) );
NAND4_X1 _14565_ ( .A1(_05965_ ), .A2(_05966_ ), .A3(_05967_ ), .A4(_05968_ ), .ZN(_06544_ ) );
OAI21_X1 _14566_ ( .A(_06543_ ), .B1(_06544_ ), .B2(_05530_ ), .ZN(_06545_ ) );
AOI22_X1 _14567_ ( .A1(_05007_ ), .A2(_05851_ ), .B1(\ID_EX_typ [2] ), .B2(_06545_ ), .ZN(_06546_ ) );
OAI211_X1 _14568_ ( .A(_06546_ ), .B(_06225_ ), .C1(_05932_ ), .C2(\ID_EX_imm [31] ), .ZN(_06547_ ) );
AND4_X1 _14569_ ( .A1(_05967_ ), .A2(_05965_ ), .A3(_05966_ ), .A4(_05968_ ), .ZN(_06548_ ) );
AOI21_X1 _14570_ ( .A(_06542_ ), .B1(_06548_ ), .B2(_05531_ ), .ZN(_06549_ ) );
NAND3_X1 _14571_ ( .A1(_06549_ ), .A2(_06377_ ), .A3(_06434_ ), .ZN(_06550_ ) );
AND3_X1 _14572_ ( .A1(_03354_ ), .A2(\ID_EX_pc [31] ), .A3(\ID_EX_typ [7] ), .ZN(_06551_ ) );
AOI21_X1 _14573_ ( .A(_06551_ ), .B1(_04633_ ), .B2(_06425_ ), .ZN(_06552_ ) );
OAI211_X1 _14574_ ( .A(_06547_ ), .B(_06550_ ), .C1(_06393_ ), .C2(_06552_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ) );
NOR2_X1 _14575_ ( .A1(_05947_ ), .A2(_05949_ ), .ZN(_06553_ ) );
NAND4_X1 _14576_ ( .A1(_06553_ ), .A2(_05293_ ), .A3(_05719_ ), .A4(_05946_ ), .ZN(_06554_ ) );
NAND3_X1 _14577_ ( .A1(_05840_ ), .A2(_05841_ ), .A3(_06109_ ), .ZN(_06555_ ) );
BUF_X4 _14578_ ( .A(_06222_ ), .Z(_06556_ ) );
NAND3_X1 _14579_ ( .A1(_06554_ ), .A2(_06555_ ), .A3(_06556_ ), .ZN(_06557_ ) );
NOR3_X1 _14580_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [0] ), .A3(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06558_ ) );
AND2_X1 _14581_ ( .A1(\ID_EX_typ [3] ), .A2(\ID_EX_typ [2] ), .ZN(_06559_ ) );
AND2_X2 _14582_ ( .A1(_06558_ ), .A2(_06559_ ), .ZN(_06560_ ) );
INV_X1 _14583_ ( .A(_06560_ ), .ZN(_06561_ ) );
NOR3_X1 _14584_ ( .A1(_04767_ ), .A2(\ID_EX_typ [0] ), .A3(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06562_ ) );
AND2_X1 _14585_ ( .A1(_06562_ ), .A2(_06559_ ), .ZN(_06563_ ) );
BUF_X4 _14586_ ( .A(_06563_ ), .Z(_06564_ ) );
INV_X1 _14587_ ( .A(_06564_ ), .ZN(_06565_ ) );
BUF_X4 _14588_ ( .A(_06565_ ), .Z(_06566_ ) );
OAI22_X1 _14589_ ( .A1(_05942_ ), .A2(_06561_ ), .B1(_02298_ ), .B2(_06566_ ), .ZN(_06567_ ) );
OR2_X1 _14590_ ( .A1(_05059_ ), .A2(_04462_ ), .ZN(_06568_ ) );
AND2_X1 _14591_ ( .A1(_06568_ ), .A2(_05085_ ), .ZN(_06569_ ) );
NOR2_X1 _14592_ ( .A1(_06569_ ), .A2(_04488_ ), .ZN(_06570_ ) );
XNOR2_X1 _14593_ ( .A(_04510_ ), .B(_04978_ ), .ZN(_06571_ ) );
NOR3_X1 _14594_ ( .A1(_06570_ ), .A2(_05087_ ), .A3(_06571_ ), .ZN(_06572_ ) );
AND3_X1 _14595_ ( .A1(_03913_ ), .A2(\ID_EX_typ [3] ), .A3(_04769_ ), .ZN(_06573_ ) );
AND2_X1 _14596_ ( .A1(_06573_ ), .A2(_04787_ ), .ZN(_06574_ ) );
INV_X1 _14597_ ( .A(_06574_ ), .ZN(_06575_ ) );
BUF_X4 _14598_ ( .A(_06575_ ), .Z(_06576_ ) );
NOR2_X1 _14599_ ( .A1(_06572_ ), .A2(_06576_ ), .ZN(_06577_ ) );
OAI21_X1 _14600_ ( .A(_06571_ ), .B1(_06570_ ), .B2(_05087_ ), .ZN(_06578_ ) );
AOI21_X1 _14601_ ( .A(_06567_ ), .B1(_06577_ ), .B2(_06578_ ), .ZN(_06579_ ) );
NOR2_X1 _14602_ ( .A1(_06210_ ), .A2(\ID_EX_typ [6] ), .ZN(_06580_ ) );
AND2_X1 _14603_ ( .A1(_06580_ ), .A2(_03341_ ), .ZN(_06581_ ) );
BUF_X4 _14604_ ( .A(_06581_ ), .Z(_06582_ ) );
INV_X1 _14605_ ( .A(_06582_ ), .ZN(_06583_ ) );
BUF_X4 _14606_ ( .A(_06583_ ), .Z(_06584_ ) );
OAI21_X1 _14607_ ( .A(_05928_ ), .B1(_06579_ ), .B2(_06584_ ), .ZN(_06585_ ) );
BUF_X4 _14608_ ( .A(_04765_ ), .Z(_06586_ ) );
NOR2_X1 _14609_ ( .A1(\ID_EX_typ [2] ), .A2(\ID_EX_typ [1] ), .ZN(_06587_ ) );
INV_X1 _14610_ ( .A(_06587_ ), .ZN(_06588_ ) );
NOR2_X1 _14611_ ( .A1(_06586_ ), .A2(_06588_ ), .ZN(_06589_ ) );
INV_X1 _14612_ ( .A(_06589_ ), .ZN(_06590_ ) );
INV_X1 _14613_ ( .A(_04917_ ), .ZN(_06591_ ) );
NOR2_X1 _14614_ ( .A1(_04847_ ), .A2(_04022_ ), .ZN(_06592_ ) );
AOI21_X1 _14615_ ( .A(_04918_ ), .B1(_06591_ ), .B2(_06592_ ), .ZN(_06593_ ) );
INV_X1 _14616_ ( .A(_06593_ ), .ZN(_06594_ ) );
AND2_X1 _14617_ ( .A1(_04853_ ), .A2(_04857_ ), .ZN(_06595_ ) );
AND2_X1 _14618_ ( .A1(_06594_ ), .A2(_06595_ ), .ZN(_06596_ ) );
NOR2_X1 _14619_ ( .A1(_04852_ ), .A2(_03916_ ), .ZN(_06597_ ) );
INV_X1 _14620_ ( .A(_02742_ ), .ZN(_06598_ ) );
NOR2_X1 _14621_ ( .A1(_04856_ ), .A2(_06598_ ), .ZN(_06599_ ) );
AND2_X1 _14622_ ( .A1(_04853_ ), .A2(_06599_ ), .ZN(_06600_ ) );
NOR3_X1 _14623_ ( .A1(_06596_ ), .A2(_06597_ ), .A3(_06600_ ), .ZN(_06601_ ) );
AND2_X1 _14624_ ( .A1(_04832_ ), .A2(_04837_ ), .ZN(_06602_ ) );
XNOR2_X1 _14625_ ( .A(_04824_ ), .B(_02718_ ), .ZN(_06603_ ) );
AND3_X1 _14626_ ( .A1(_06602_ ), .A2(_04821_ ), .A3(_06603_ ), .ZN(_06604_ ) );
INV_X1 _14627_ ( .A(_06604_ ), .ZN(_06605_ ) );
NOR2_X1 _14628_ ( .A1(_06601_ ), .A2(_06605_ ), .ZN(_06606_ ) );
NOR2_X1 _14629_ ( .A1(_04820_ ), .A2(_04109_ ), .ZN(_06607_ ) );
INV_X1 _14630_ ( .A(_06603_ ), .ZN(_06608_ ) );
NOR2_X1 _14631_ ( .A1(_04831_ ), .A2(_06315_ ), .ZN(_06609_ ) );
NOR2_X1 _14632_ ( .A1(_04836_ ), .A2(_04079_ ), .ZN(_06610_ ) );
AOI21_X1 _14633_ ( .A(_06609_ ), .B1(_04832_ ), .B2(_06610_ ), .ZN(_06611_ ) );
NOR3_X1 _14634_ ( .A1(_06608_ ), .A2(_06611_ ), .A3(_04931_ ), .ZN(_06612_ ) );
AND2_X1 _14635_ ( .A1(_04821_ ), .A2(_04825_ ), .ZN(_06613_ ) );
NOR4_X1 _14636_ ( .A1(_06606_ ), .A2(_06607_ ), .A3(_06612_ ), .A4(_06613_ ), .ZN(_06614_ ) );
NAND2_X1 _14637_ ( .A1(_04843_ ), .A2(_04848_ ), .ZN(_06615_ ) );
INV_X1 _14638_ ( .A(_04884_ ), .ZN(_06616_ ) );
NOR2_X1 _14639_ ( .A1(_04880_ ), .A2(_02493_ ), .ZN(_06617_ ) );
INV_X1 _14640_ ( .A(_06617_ ), .ZN(_06618_ ) );
NOR2_X1 _14641_ ( .A1(_06479_ ), .A2(_04869_ ), .ZN(_06619_ ) );
INV_X1 _14642_ ( .A(_06619_ ), .ZN(_06620_ ) );
NOR3_X2 _14643_ ( .A1(_04864_ ), .A2(_06620_ ), .A3(_04865_ ), .ZN(_06621_ ) );
NOR2_X2 _14644_ ( .A1(_06621_ ), .A2(_04864_ ), .ZN(_06622_ ) );
INV_X1 _14645_ ( .A(_04881_ ), .ZN(_06623_ ) );
OAI211_X2 _14646_ ( .A(_06616_ ), .B(_06618_ ), .C1(_06622_ ), .C2(_06623_ ), .ZN(_06624_ ) );
INV_X1 _14647_ ( .A(_04885_ ), .ZN(_06625_ ) );
AND3_X1 _14648_ ( .A1(_04895_ ), .A2(_04891_ ), .A3(_04896_ ), .ZN(_06626_ ) );
AND2_X1 _14649_ ( .A1(_04902_ ), .A2(_04907_ ), .ZN(_06627_ ) );
NAND4_X2 _14650_ ( .A1(_06624_ ), .A2(_06625_ ), .A3(_06626_ ), .A4(_06627_ ), .ZN(_06628_ ) );
INV_X1 _14651_ ( .A(_02543_ ), .ZN(_06629_ ) );
NOR2_X1 _14652_ ( .A1(_06629_ ), .A2(_04890_ ), .ZN(_06630_ ) );
AOI21_X1 _14653_ ( .A(_02543_ ), .B1(_04888_ ), .B2(_04889_ ), .ZN(_06631_ ) );
NOR4_X1 _14654_ ( .A1(_04894_ ), .A2(_04189_ ), .A3(_06630_ ), .A4(_06631_ ), .ZN(_06632_ ) );
AND2_X1 _14655_ ( .A1(_04900_ ), .A2(_02589_ ), .ZN(_06633_ ) );
NOR2_X1 _14656_ ( .A1(_04906_ ), .A2(_04258_ ), .ZN(_06634_ ) );
AOI21_X1 _14657_ ( .A(_06633_ ), .B1(_04902_ ), .B2(_06634_ ), .ZN(_06635_ ) );
INV_X1 _14658_ ( .A(_06635_ ), .ZN(_06636_ ) );
AOI211_X1 _14659_ ( .A(_06630_ ), .B(_06632_ ), .C1(_06636_ ), .C2(_06626_ ), .ZN(_06637_ ) );
AOI21_X2 _14660_ ( .A(_06615_ ), .B1(_06628_ ), .B2(_06637_ ), .ZN(_06638_ ) );
NAND3_X1 _14661_ ( .A1(_06638_ ), .A2(_06604_ ), .A3(_06595_ ), .ZN(_06639_ ) );
AND2_X1 _14662_ ( .A1(_06614_ ), .A2(_06639_ ), .ZN(_06640_ ) );
INV_X2 _14663_ ( .A(_06640_ ), .ZN(_06641_ ) );
AND2_X1 _14664_ ( .A1(_04968_ ), .A2(_04972_ ), .ZN(_06642_ ) );
NAND4_X1 _14665_ ( .A1(_06641_ ), .A2(_04960_ ), .A3(_04964_ ), .A4(_06642_ ), .ZN(_06643_ ) );
NOR2_X1 _14666_ ( .A1(_04967_ ), .A2(_04430_ ), .ZN(_06644_ ) );
NOR2_X1 _14667_ ( .A1(_04971_ ), .A2(_04432_ ), .ZN(_06645_ ) );
AOI21_X1 _14668_ ( .A(_06644_ ), .B1(_04968_ ), .B2(_06645_ ), .ZN(_06646_ ) );
INV_X1 _14669_ ( .A(_06646_ ), .ZN(_06647_ ) );
AND3_X1 _14670_ ( .A1(_06647_ ), .A2(_04960_ ), .A3(_04964_ ), .ZN(_06648_ ) );
OR2_X1 _14671_ ( .A1(_04959_ ), .A2(_04383_ ), .ZN(_06649_ ) );
NOR2_X1 _14672_ ( .A1(_04963_ ), .A2(_04357_ ), .ZN(_06650_ ) );
INV_X1 _14673_ ( .A(_06650_ ), .ZN(_06651_ ) );
AND3_X1 _14674_ ( .A1(_04957_ ), .A2(_04383_ ), .A3(_04958_ ), .ZN(_06652_ ) );
OAI21_X1 _14675_ ( .A(_06649_ ), .B1(_06651_ ), .B2(_06652_ ), .ZN(_06653_ ) );
NOR2_X1 _14676_ ( .A1(_06648_ ), .A2(_06653_ ), .ZN(_06654_ ) );
AND2_X2 _14677_ ( .A1(_06643_ ), .A2(_06654_ ), .ZN(_06655_ ) );
INV_X2 _14678_ ( .A(_06655_ ), .ZN(_06656_ ) );
NAND2_X1 _14679_ ( .A1(_06656_ ), .A2(_04955_ ), .ZN(_06657_ ) );
NOR2_X1 _14680_ ( .A1(_04954_ ), .A2(_06244_ ), .ZN(_06658_ ) );
INV_X1 _14681_ ( .A(_06658_ ), .ZN(_06659_ ) );
NAND2_X1 _14682_ ( .A1(_06657_ ), .A2(_06659_ ), .ZN(_06660_ ) );
AOI21_X1 _14683_ ( .A(_06590_ ), .B1(_06660_ ), .B2(_04951_ ), .ZN(_06661_ ) );
OAI21_X1 _14684_ ( .A(_06661_ ), .B1(_04951_ ), .B2(_06660_ ), .ZN(_06662_ ) );
INV_X1 _14685_ ( .A(_04869_ ), .ZN(_06663_ ) );
BUF_X4 _14686_ ( .A(_06663_ ), .Z(_06664_ ) );
NAND3_X1 _14687_ ( .A1(_06664_ ), .A2(_02961_ ), .A3(_02962_ ), .ZN(_06665_ ) );
BUF_X4 _14688_ ( .A(_04869_ ), .Z(_06666_ ) );
NAND2_X1 _14689_ ( .A1(_02940_ ), .A2(_06666_ ), .ZN(_06667_ ) );
NAND2_X1 _14690_ ( .A1(_06665_ ), .A2(_06667_ ), .ZN(_06668_ ) );
BUF_X4 _14691_ ( .A(_04872_ ), .Z(_06669_ ) );
NAND2_X1 _14692_ ( .A1(_06668_ ), .A2(_06669_ ), .ZN(_06670_ ) );
BUF_X4 _14693_ ( .A(_04872_ ), .Z(_06671_ ) );
BUF_X4 _14694_ ( .A(_06666_ ), .Z(_06672_ ) );
AND2_X1 _14695_ ( .A1(_02990_ ), .A2(_06672_ ), .ZN(_06673_ ) );
OAI21_X1 _14696_ ( .A(_06670_ ), .B1(_06671_ ), .B2(_06673_ ), .ZN(_06674_ ) );
INV_X2 _14697_ ( .A(_04880_ ), .ZN(_06675_ ) );
BUF_X4 _14698_ ( .A(_06675_ ), .Z(_06676_ ) );
BUF_X2 _14699_ ( .A(_06676_ ), .Z(_06677_ ) );
NOR2_X1 _14700_ ( .A1(_06674_ ), .A2(_06677_ ), .ZN(_06678_ ) );
NOR2_X1 _14701_ ( .A1(_06666_ ), .A2(_02196_ ), .ZN(_06679_ ) );
INV_X1 _14702_ ( .A(_06679_ ), .ZN(_06680_ ) );
OAI211_X1 _14703_ ( .A(_06671_ ), .B(_06680_ ), .C1(_02899_ ), .C2(_06664_ ), .ZN(_06681_ ) );
BUF_X2 _14704_ ( .A(_06675_ ), .Z(_06682_ ) );
NOR2_X1 _14705_ ( .A1(_06666_ ), .A2(_02167_ ), .ZN(_06683_ ) );
INV_X1 _14706_ ( .A(_06683_ ), .ZN(_06684_ ) );
BUF_X4 _14707_ ( .A(_04867_ ), .Z(_06685_ ) );
BUF_X4 _14708_ ( .A(_04868_ ), .Z(_06686_ ) );
AOI21_X1 _14709_ ( .A(_04707_ ), .B1(_06685_ ), .B2(_06686_ ), .ZN(_06687_ ) );
INV_X1 _14710_ ( .A(_06687_ ), .ZN(_06688_ ) );
BUF_X4 _14711_ ( .A(_04861_ ), .Z(_06689_ ) );
BUF_X4 _14712_ ( .A(_04863_ ), .Z(_06690_ ) );
NAND4_X1 _14713_ ( .A1(_06684_ ), .A2(_06688_ ), .A3(_06689_ ), .A4(_06690_ ), .ZN(_06691_ ) );
AND3_X1 _14714_ ( .A1(_06681_ ), .A2(_06682_ ), .A3(_06691_ ), .ZN(_06692_ ) );
BUF_X4 _14715_ ( .A(_06676_ ), .Z(_06693_ ) );
AOI21_X1 _14716_ ( .A(_04511_ ), .B1(_06685_ ), .B2(_06686_ ), .ZN(_06694_ ) );
NOR2_X1 _14717_ ( .A1(_06666_ ), .A2(_02270_ ), .ZN(_06695_ ) );
OAI21_X1 _14718_ ( .A(_06669_ ), .B1(_06694_ ), .B2(_06695_ ), .ZN(_06696_ ) );
NOR2_X1 _14719_ ( .A1(_06666_ ), .A2(_02876_ ), .ZN(_06697_ ) );
AOI21_X1 _14720_ ( .A(_02247_ ), .B1(_06685_ ), .B2(_06686_ ), .ZN(_06698_ ) );
OAI211_X1 _14721_ ( .A(_04861_ ), .B(_04863_ ), .C1(_06697_ ), .C2(_06698_ ), .ZN(_06699_ ) );
AOI21_X1 _14722_ ( .A(_06693_ ), .B1(_06696_ ), .B2(_06699_ ), .ZN(_06700_ ) );
NOR2_X1 _14723_ ( .A1(_06692_ ), .A2(_06700_ ), .ZN(_06701_ ) );
INV_X1 _14724_ ( .A(_04876_ ), .ZN(_06702_ ) );
BUF_X4 _14725_ ( .A(_06702_ ), .Z(_06703_ ) );
BUF_X4 _14726_ ( .A(_06703_ ), .Z(_06704_ ) );
MUX2_X1 _14727_ ( .A(_06678_ ), .B(_06701_ ), .S(_06704_ ), .Z(_06705_ ) );
BUF_X2 _14728_ ( .A(_04906_ ), .Z(_06706_ ) );
BUF_X2 _14729_ ( .A(_06706_ ), .Z(_06707_ ) );
BUF_X2 _14730_ ( .A(_06707_ ), .Z(_06708_ ) );
AND2_X2 _14731_ ( .A1(_04768_ ), .A2(\ID_EX_typ [2] ), .ZN(_06709_ ) );
BUF_X2 _14732_ ( .A(_06709_ ), .Z(_06710_ ) );
BUF_X2 _14733_ ( .A(_06710_ ), .Z(_06711_ ) );
NAND3_X1 _14734_ ( .A1(_06705_ ), .A2(_06708_ ), .A3(_06711_ ), .ZN(_06712_ ) );
BUF_X2 _14735_ ( .A(_04771_ ), .Z(_06713_ ) );
OAI211_X1 _14736_ ( .A(_06662_ ), .B(_06712_ ), .C1(_04979_ ), .C2(_06713_ ), .ZN(_06714_ ) );
AND2_X1 _14737_ ( .A1(_05024_ ), .A2(\ID_EX_typ [2] ), .ZN(_06715_ ) );
BUF_X4 _14738_ ( .A(_06715_ ), .Z(_06716_ ) );
INV_X1 _14739_ ( .A(_06716_ ), .ZN(_06717_ ) );
BUF_X4 _14740_ ( .A(_06717_ ), .Z(_06718_ ) );
OR2_X1 _14741_ ( .A1(_04894_ ), .A2(_04890_ ), .ZN(_06719_ ) );
AND2_X1 _14742_ ( .A1(_04872_ ), .A2(_04869_ ), .ZN(_06720_ ) );
AND2_X1 _14743_ ( .A1(_06720_ ), .A2(_04880_ ), .ZN(_06721_ ) );
AND2_X4 _14744_ ( .A1(_06721_ ), .A2(_06702_ ), .ZN(_06722_ ) );
AOI221_X4 _14745_ ( .A(_06719_ ), .B1(_04898_ ), .B2(_04899_ ), .C1(_06722_ ), .C2(_06706_ ), .ZN(_06723_ ) );
AND3_X1 _14746_ ( .A1(_04892_ ), .A2(_04890_ ), .A3(_04893_ ), .ZN(_06724_ ) );
NAND4_X1 _14747_ ( .A1(_06722_ ), .A2(_04900_ ), .A3(_04906_ ), .A4(_06724_ ), .ZN(_06725_ ) );
NAND4_X1 _14748_ ( .A1(_04894_ ), .A2(_04890_ ), .A3(_04898_ ), .A4(_04899_ ), .ZN(_06726_ ) );
NAND2_X1 _14749_ ( .A1(_06725_ ), .A2(_06726_ ), .ZN(_06727_ ) );
OAI21_X1 _14750_ ( .A(_02990_ ), .B1(_06723_ ), .B2(_06727_ ), .ZN(_06728_ ) );
AND3_X1 _14751_ ( .A1(_04847_ ), .A2(_04841_ ), .A3(_04840_ ), .ZN(_06729_ ) );
AND2_X1 _14752_ ( .A1(_06727_ ), .A2(_06729_ ), .ZN(_06730_ ) );
INV_X1 _14753_ ( .A(_06730_ ), .ZN(_06731_ ) );
OR3_X1 _14754_ ( .A1(_06727_ ), .A2(_04842_ ), .A3(_04847_ ), .ZN(_06732_ ) );
OR3_X1 _14755_ ( .A1(_06730_ ), .A2(_04852_ ), .A3(_04856_ ), .ZN(_06733_ ) );
NAND3_X1 _14756_ ( .A1(_06727_ ), .A2(_04856_ ), .A3(_06729_ ), .ZN(_06734_ ) );
NOR2_X2 _14757_ ( .A1(_06734_ ), .A2(_04924_ ), .ZN(_06735_ ) );
INV_X1 _14758_ ( .A(_06735_ ), .ZN(_06736_ ) );
AOI221_X2 _14759_ ( .A(_06728_ ), .B1(_06731_ ), .B2(_06732_ ), .C1(_06733_ ), .C2(_06736_ ), .ZN(_06737_ ) );
AND3_X1 _14760_ ( .A1(_04824_ ), .A2(_04831_ ), .A3(_04836_ ), .ZN(_06738_ ) );
NOR4_X1 _14761_ ( .A1(_04783_ ), .A2(_05018_ ), .A3(_04777_ ), .A4(_05012_ ), .ZN(_06739_ ) );
AOI22_X1 _14762_ ( .A1(_04796_ ), .A2(_04797_ ), .B1(_04788_ ), .B2(_04789_ ), .ZN(_06740_ ) );
AND4_X1 _14763_ ( .A1(_04806_ ), .A2(_06739_ ), .A3(_04813_ ), .A4(_06740_ ), .ZN(_06741_ ) );
AND3_X1 _14764_ ( .A1(_04963_ ), .A2(_04957_ ), .A3(_04958_ ), .ZN(_06742_ ) );
AND3_X1 _14765_ ( .A1(_06742_ ), .A2(_04967_ ), .A3(_04971_ ), .ZN(_06743_ ) );
AND4_X1 _14766_ ( .A1(_04942_ ), .A2(_04938_ ), .A3(_04950_ ), .A4(_04954_ ), .ZN(_06744_ ) );
NAND3_X1 _14767_ ( .A1(_06741_ ), .A2(_06743_ ), .A3(_06744_ ), .ZN(_06745_ ) );
NAND4_X1 _14768_ ( .A1(_06735_ ), .A2(_04820_ ), .A3(_06738_ ), .A4(_06745_ ), .ZN(_06746_ ) );
NAND2_X1 _14769_ ( .A1(_06737_ ), .A2(_06746_ ), .ZN(_06747_ ) );
NAND3_X1 _14770_ ( .A1(_06735_ ), .A2(_04820_ ), .A3(_06738_ ), .ZN(_06748_ ) );
NOR4_X1 _14771_ ( .A1(_04938_ ), .A2(_04942_ ), .A3(_04950_ ), .A4(_04954_ ), .ZN(_06749_ ) );
AOI22_X1 _14772_ ( .A1(_04965_ ), .A2(_04966_ ), .B1(_04969_ ), .B2(_04970_ ), .ZN(_06750_ ) );
NAND4_X1 _14773_ ( .A1(_06749_ ), .A2(_04989_ ), .A3(_04991_ ), .A4(_06750_ ), .ZN(_06751_ ) );
OR4_X1 _14774_ ( .A1(_04820_ ), .A2(_04824_ ), .A3(_04831_ ), .A4(_04836_ ), .ZN(_06752_ ) );
NOR2_X1 _14775_ ( .A1(_06751_ ), .A2(_06752_ ), .ZN(_06753_ ) );
INV_X1 _14776_ ( .A(_04783_ ), .ZN(_06754_ ) );
NOR4_X1 _14777_ ( .A1(_06754_ ), .A2(_05019_ ), .A3(_04806_ ), .A4(_04813_ ), .ZN(_06755_ ) );
AND4_X1 _14778_ ( .A1(_04796_ ), .A2(_06755_ ), .A3(_04797_ ), .A4(_05012_ ), .ZN(_06756_ ) );
AND4_X1 _14779_ ( .A1(_04999_ ), .A2(_06753_ ), .A3(_05018_ ), .A4(_06756_ ), .ZN(_06757_ ) );
OAI21_X1 _14780_ ( .A(_06757_ ), .B1(_06734_ ), .B2(_04924_ ), .ZN(_06758_ ) );
AND2_X2 _14781_ ( .A1(_06748_ ), .A2(_06758_ ), .ZN(_06759_ ) );
NOR2_X4 _14782_ ( .A1(_06747_ ), .A2(_06759_ ), .ZN(_06760_ ) );
AND2_X1 _14783_ ( .A1(_06722_ ), .A2(_06706_ ), .ZN(_06761_ ) );
XNOR2_X1 _14784_ ( .A(_06761_ ), .B(_04900_ ), .ZN(_06762_ ) );
AND2_X2 _14785_ ( .A1(_06760_ ), .A2(_06762_ ), .ZN(_06763_ ) );
XNOR2_X1 _14786_ ( .A(_06722_ ), .B(_06706_ ), .ZN(_06764_ ) );
NOR2_X1 _14787_ ( .A1(_06764_ ), .A2(_04900_ ), .ZN(_06765_ ) );
BUF_X2 _14788_ ( .A(_06764_ ), .Z(_06766_ ) );
BUF_X4 _14789_ ( .A(_06669_ ), .Z(_06767_ ) );
BUF_X4 _14790_ ( .A(_06672_ ), .Z(_06768_ ) );
XNOR2_X1 _14791_ ( .A(_06767_ ), .B(_06768_ ), .ZN(_06769_ ) );
NOR2_X1 _14792_ ( .A1(_06769_ ), .A2(_06693_ ), .ZN(_06770_ ) );
XNOR2_X1 _14793_ ( .A(_06721_ ), .B(_04876_ ), .ZN(_06771_ ) );
NOR4_X1 _14794_ ( .A1(_06747_ ), .A2(_06770_ ), .A3(_06771_ ), .A4(_06759_ ), .ZN(_06772_ ) );
OAI22_X1 _14795_ ( .A1(_06763_ ), .A2(_06765_ ), .B1(_06766_ ), .B2(_06772_ ), .ZN(_06773_ ) );
NAND2_X1 _14796_ ( .A1(_06705_ ), .A2(_06708_ ), .ZN(_06774_ ) );
AOI21_X1 _14797_ ( .A(_06718_ ), .B1(_06773_ ), .B2(_06774_ ), .ZN(_06775_ ) );
INV_X1 _14798_ ( .A(_05099_ ), .ZN(_06776_ ) );
INV_X1 _14799_ ( .A(_04872_ ), .ZN(_06777_ ) );
BUF_X4 _14800_ ( .A(_06685_ ), .Z(_06778_ ) );
BUF_X4 _14801_ ( .A(_06686_ ), .Z(_06779_ ) );
AOI21_X1 _14802_ ( .A(_04075_ ), .B1(_06778_ ), .B2(_06779_ ), .ZN(_06780_ ) );
NOR2_X1 _14803_ ( .A1(_06672_ ), .A2(_02647_ ), .ZN(_06781_ ) );
OR3_X1 _14804_ ( .A1(_06777_ ), .A2(_06780_ ), .A3(_06781_ ), .ZN(_06782_ ) );
BUF_X4 _14805_ ( .A(_06666_ ), .Z(_06783_ ) );
NOR2_X1 _14806_ ( .A1(_06783_ ), .A2(_02742_ ), .ZN(_06784_ ) );
INV_X1 _14807_ ( .A(_06784_ ), .ZN(_06785_ ) );
AOI21_X1 _14808_ ( .A(_02765_ ), .B1(_06778_ ), .B2(_06779_ ), .ZN(_06786_ ) );
INV_X1 _14809_ ( .A(_06786_ ), .ZN(_06787_ ) );
NAND4_X1 _14810_ ( .A1(_06785_ ), .A2(_06787_ ), .A3(_06689_ ), .A4(_06690_ ), .ZN(_06788_ ) );
AOI21_X1 _14811_ ( .A(_06675_ ), .B1(_06782_ ), .B2(_06788_ ), .ZN(_06789_ ) );
BUF_X4 _14812_ ( .A(_04880_ ), .Z(_06790_ ) );
BUF_X4 _14813_ ( .A(_06790_ ), .Z(_06791_ ) );
BUF_X4 _14814_ ( .A(_06685_ ), .Z(_06792_ ) );
BUF_X4 _14815_ ( .A(_06686_ ), .Z(_06793_ ) );
AOI21_X1 _14816_ ( .A(_02543_ ), .B1(_06792_ ), .B2(_06793_ ), .ZN(_06794_ ) );
INV_X1 _14817_ ( .A(_06794_ ), .ZN(_06795_ ) );
OAI211_X1 _14818_ ( .A(_06777_ ), .B(_06795_ ), .C1(_02565_ ), .C2(_06768_ ), .ZN(_06796_ ) );
BUF_X4 _14819_ ( .A(_06669_ ), .Z(_06797_ ) );
NOR2_X1 _14820_ ( .A1(_06783_ ), .A2(_02789_ ), .ZN(_06798_ ) );
INV_X1 _14821_ ( .A(_06798_ ), .ZN(_06799_ ) );
AOI21_X1 _14822_ ( .A(_02812_ ), .B1(_06792_ ), .B2(_06793_ ), .ZN(_06800_ ) );
INV_X1 _14823_ ( .A(_06800_ ), .ZN(_06801_ ) );
NAND3_X1 _14824_ ( .A1(_06797_ ), .A2(_06799_ ), .A3(_06801_ ), .ZN(_06802_ ) );
AOI21_X1 _14825_ ( .A(_06791_ ), .B1(_06796_ ), .B2(_06802_ ), .ZN(_06803_ ) );
OR3_X1 _14826_ ( .A1(_06789_ ), .A2(_06703_ ), .A3(_06803_ ), .ZN(_06804_ ) );
BUF_X4 _14827_ ( .A(_06791_ ), .Z(_06805_ ) );
AOI21_X1 _14828_ ( .A(_02394_ ), .B1(_06778_ ), .B2(_06779_ ), .ZN(_06806_ ) );
NOR2_X1 _14829_ ( .A1(_06672_ ), .A2(_02417_ ), .ZN(_06807_ ) );
OR3_X1 _14830_ ( .A1(_06777_ ), .A2(_06806_ ), .A3(_06807_ ), .ZN(_06808_ ) );
AOI21_X1 _14831_ ( .A(_02694_ ), .B1(_06792_ ), .B2(_06793_ ), .ZN(_06809_ ) );
INV_X1 _14832_ ( .A(_06809_ ), .ZN(_06810_ ) );
OAI211_X1 _14833_ ( .A(_06777_ ), .B(_06810_ ), .C1(_02718_ ), .C2(_06768_ ), .ZN(_06811_ ) );
AOI21_X1 _14834_ ( .A(_06805_ ), .B1(_06808_ ), .B2(_06811_ ), .ZN(_06812_ ) );
BUF_X4 _14835_ ( .A(_04876_ ), .Z(_06813_ ) );
BUF_X2 _14836_ ( .A(_06813_ ), .Z(_06814_ ) );
BUF_X4 _14837_ ( .A(_06671_ ), .Z(_06815_ ) );
NOR2_X1 _14838_ ( .A1(_06666_ ), .A2(_02294_ ), .ZN(_06816_ ) );
OAI21_X1 _14839_ ( .A(_06815_ ), .B1(_06694_ ), .B2(_06816_ ), .ZN(_06817_ ) );
BUF_X2 _14840_ ( .A(_06790_ ), .Z(_06818_ ) );
BUF_X4 _14841_ ( .A(_04861_ ), .Z(_06819_ ) );
BUF_X4 _14842_ ( .A(_06690_ ), .Z(_06820_ ) );
NOR2_X1 _14843_ ( .A1(_06672_ ), .A2(_02346_ ), .ZN(_06821_ ) );
AOI21_X1 _14844_ ( .A(_02370_ ), .B1(_06685_ ), .B2(_06686_ ), .ZN(_06822_ ) );
OAI211_X1 _14845_ ( .A(_06819_ ), .B(_06820_ ), .C1(_06821_ ), .C2(_06822_ ), .ZN(_06823_ ) );
AND3_X1 _14846_ ( .A1(_06817_ ), .A2(_06818_ ), .A3(_06823_ ), .ZN(_06824_ ) );
OR3_X1 _14847_ ( .A1(_06812_ ), .A2(_06814_ ), .A3(_06824_ ), .ZN(_06825_ ) );
NAND3_X1 _14848_ ( .A1(_06804_ ), .A2(_06825_ ), .A3(_06707_ ), .ZN(_06826_ ) );
AOI21_X1 _14849_ ( .A(_02589_ ), .B1(_06792_ ), .B2(_06793_ ), .ZN(_06827_ ) );
NOR2_X1 _14850_ ( .A1(_06783_ ), .A2(_02611_ ), .ZN(_06828_ ) );
OAI21_X1 _14851_ ( .A(_06671_ ), .B1(_06827_ ), .B2(_06828_ ), .ZN(_06829_ ) );
NOR2_X1 _14852_ ( .A1(_06783_ ), .A2(_02441_ ), .ZN(_06830_ ) );
AOI21_X1 _14853_ ( .A(_02516_ ), .B1(_06792_ ), .B2(_06793_ ), .ZN(_06831_ ) );
OAI211_X1 _14854_ ( .A(_06689_ ), .B(_06690_ ), .C1(_06830_ ), .C2(_06831_ ), .ZN(_06832_ ) );
NAND3_X1 _14855_ ( .A1(_06829_ ), .A2(_06791_ ), .A3(_06832_ ), .ZN(_06833_ ) );
AOI21_X1 _14856_ ( .A(_02464_ ), .B1(_06792_ ), .B2(_06793_ ), .ZN(_06834_ ) );
NOR2_X1 _14857_ ( .A1(_04870_ ), .A2(_06834_ ), .ZN(_06835_ ) );
NAND3_X1 _14858_ ( .A1(_06835_ ), .A2(_06675_ ), .A3(_06767_ ), .ZN(_06836_ ) );
AND2_X1 _14859_ ( .A1(_06833_ ), .A2(_06836_ ), .ZN(_06837_ ) );
BUF_X2 _14860_ ( .A(_06706_ ), .Z(_06838_ ) );
BUF_X2 _14861_ ( .A(_06813_ ), .Z(_06839_ ) );
OR3_X1 _14862_ ( .A1(_06837_ ), .A2(_06838_ ), .A3(_06839_ ), .ZN(_06840_ ) );
AOI21_X1 _14863_ ( .A(_06776_ ), .B1(_06826_ ), .B2(_06840_ ), .ZN(_06841_ ) );
NOR3_X1 _14864_ ( .A1(_04979_ ), .A2(_04980_ ), .A3(_05026_ ), .ZN(_06842_ ) );
BUF_X2 _14865_ ( .A(_04766_ ), .Z(_06843_ ) );
NOR3_X1 _14866_ ( .A1(_04950_ ), .A2(_04978_ ), .A3(_06843_ ), .ZN(_06844_ ) );
OR3_X1 _14867_ ( .A1(_06841_ ), .A2(_06842_ ), .A3(_06844_ ), .ZN(_06845_ ) );
OR3_X1 _14868_ ( .A1(_06714_ ), .A2(_06775_ ), .A3(_06845_ ), .ZN(_06846_ ) );
OAI21_X1 _14869_ ( .A(_06559_ ), .B1(_06562_ ), .B2(_06558_ ), .ZN(_06847_ ) );
NOR2_X1 _14870_ ( .A1(_05318_ ), .A2(\ID_EX_typ [2] ), .ZN(_06848_ ) );
OAI211_X1 _14871_ ( .A(_06848_ ), .B(_04767_ ), .C1(_04787_ ), .C2(_03877_ ), .ZN(_06849_ ) );
AND2_X1 _14872_ ( .A1(_06847_ ), .A2(_06849_ ), .ZN(_06850_ ) );
NOR2_X1 _14873_ ( .A1(_06850_ ), .A2(_06583_ ), .ZN(_06851_ ) );
INV_X2 _14874_ ( .A(_06851_ ), .ZN(_06852_ ) );
BUF_X4 _14875_ ( .A(_06852_ ), .Z(_06853_ ) );
AOI21_X1 _14876_ ( .A(_06585_ ), .B1(_06846_ ), .B2(_06853_ ), .ZN(_06854_ ) );
BUF_X4 _14877_ ( .A(_06317_ ), .Z(_06855_ ) );
OAI21_X1 _14878_ ( .A(_06855_ ), .B1(_05937_ ), .B2(_05407_ ), .ZN(_06856_ ) );
OAI21_X1 _14879_ ( .A(_06557_ ), .B1(_06854_ ), .B2(_06856_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_10_D ) );
OAI21_X1 _14880_ ( .A(_06288_ ), .B1(_05365_ ), .B2(_05368_ ), .ZN(_06857_ ) );
BUF_X4 _14881_ ( .A(_06574_ ), .Z(_06858_ ) );
OAI21_X1 _14882_ ( .A(_06858_ ), .B1(_06569_ ), .B2(_04488_ ), .ZN(_06859_ ) );
AOI21_X1 _14883_ ( .A(_06859_ ), .B1(_04488_ ), .B2(_06569_ ), .ZN(_06860_ ) );
BUF_X2 _14884_ ( .A(_06561_ ), .Z(_06861_ ) );
OAI22_X1 _14885_ ( .A1(_05355_ ), .A2(_06861_ ), .B1(_02295_ ), .B2(_06566_ ), .ZN(_06862_ ) );
OAI21_X1 _14886_ ( .A(_06582_ ), .B1(_06860_ ), .B2(_06862_ ), .ZN(_06863_ ) );
NAND2_X1 _14887_ ( .A1(_06863_ ), .A2(_05347_ ), .ZN(_06864_ ) );
BUF_X4 _14888_ ( .A(_06716_ ), .Z(_06865_ ) );
INV_X1 _14889_ ( .A(_06771_ ), .ZN(_06866_ ) );
BUF_X2 _14890_ ( .A(_06866_ ), .Z(_06867_ ) );
BUF_X4 _14891_ ( .A(_06805_ ), .Z(_06868_ ) );
OAI21_X1 _14892_ ( .A(_06868_ ), .B1(_06777_ ), .B2(_06664_ ), .ZN(_06869_ ) );
AND3_X1 _14893_ ( .A1(_06760_ ), .A2(_06867_ ), .A3(_06869_ ), .ZN(_06870_ ) );
INV_X1 _14894_ ( .A(_06870_ ), .ZN(_06871_ ) );
INV_X1 _14895_ ( .A(_06766_ ), .ZN(_06872_ ) );
INV_X1 _14896_ ( .A(_06763_ ), .ZN(_06873_ ) );
INV_X1 _14897_ ( .A(_06765_ ), .ZN(_06874_ ) );
AOI22_X1 _14898_ ( .A1(_06871_ ), .A2(_06872_ ), .B1(_06873_ ), .B2(_06874_ ), .ZN(_06875_ ) );
INV_X1 _14899_ ( .A(_06706_ ), .ZN(_06876_ ) );
BUF_X2 _14900_ ( .A(_06876_ ), .Z(_06877_ ) );
AOI21_X1 _14901_ ( .A(_02876_ ), .B1(_06778_ ), .B2(_06779_ ), .ZN(_06878_ ) );
NOR2_X1 _14902_ ( .A1(_06672_ ), .A2(_02899_ ), .ZN(_06879_ ) );
AOI211_X1 _14903_ ( .A(_06878_ ), .B(_06879_ ), .C1(_06689_ ), .C2(_06690_ ), .ZN(_06880_ ) );
AOI21_X1 _14904_ ( .A(_02196_ ), .B1(_06778_ ), .B2(_06779_ ), .ZN(_06881_ ) );
NOR2_X1 _14905_ ( .A1(_06783_ ), .A2(_04707_ ), .ZN(_06882_ ) );
NOR3_X1 _14906_ ( .A1(_06671_ ), .A2(_06881_ ), .A3(_06882_ ), .ZN(_06883_ ) );
NOR3_X1 _14907_ ( .A1(_06880_ ), .A2(_06883_ ), .A3(_06818_ ), .ZN(_06884_ ) );
AOI21_X1 _14908_ ( .A(_02294_ ), .B1(_06778_ ), .B2(_06779_ ), .ZN(_06885_ ) );
NOR2_X1 _14909_ ( .A1(_06672_ ), .A2(_04511_ ), .ZN(_06886_ ) );
OAI21_X1 _14910_ ( .A(_06767_ ), .B1(_06885_ ), .B2(_06886_ ), .ZN(_06887_ ) );
BUF_X4 _14911_ ( .A(_04861_ ), .Z(_06888_ ) );
BUF_X4 _14912_ ( .A(_04863_ ), .Z(_06889_ ) );
NOR2_X1 _14913_ ( .A1(_06783_ ), .A2(_02247_ ), .ZN(_06890_ ) );
AOI21_X1 _14914_ ( .A(_02270_ ), .B1(_06685_ ), .B2(_06686_ ), .ZN(_06891_ ) );
OAI211_X1 _14915_ ( .A(_06888_ ), .B(_06889_ ), .C1(_06890_ ), .C2(_06891_ ), .ZN(_06892_ ) );
AOI21_X1 _14916_ ( .A(_06676_ ), .B1(_06887_ ), .B2(_06892_ ), .ZN(_06893_ ) );
OR3_X1 _14917_ ( .A1(_06884_ ), .A2(_06839_ ), .A3(_06893_ ), .ZN(_06894_ ) );
AND3_X1 _14918_ ( .A1(_06666_ ), .A2(_02961_ ), .A3(_02962_ ), .ZN(_06895_ ) );
AOI21_X1 _14919_ ( .A(_06895_ ), .B1(_05007_ ), .B2(_06664_ ), .ZN(_06896_ ) );
NOR2_X1 _14920_ ( .A1(_06783_ ), .A2(_02934_ ), .ZN(_06897_ ) );
AOI21_X1 _14921_ ( .A(_02167_ ), .B1(_06778_ ), .B2(_06779_ ), .ZN(_06898_ ) );
NOR2_X1 _14922_ ( .A1(_06897_ ), .A2(_06898_ ), .ZN(_06899_ ) );
MUX2_X1 _14923_ ( .A(_06896_ ), .B(_06899_ ), .S(_06797_ ), .Z(_06900_ ) );
BUF_X2 _14924_ ( .A(_06814_ ), .Z(_06901_ ) );
NAND3_X1 _14925_ ( .A1(_06900_ ), .A2(_06901_ ), .A3(_06868_ ), .ZN(_06902_ ) );
AOI21_X1 _14926_ ( .A(_06877_ ), .B1(_06894_ ), .B2(_06902_ ), .ZN(_06903_ ) );
OAI21_X1 _14927_ ( .A(_06865_ ), .B1(_06875_ ), .B2(_06903_ ), .ZN(_06904_ ) );
BUF_X2 _14928_ ( .A(_06590_ ), .Z(_06905_ ) );
AOI21_X1 _14929_ ( .A(_06905_ ), .B1(_06656_ ), .B2(_04955_ ), .ZN(_06906_ ) );
OAI21_X1 _14930_ ( .A(_06906_ ), .B1(_04955_ ), .B2(_06656_ ), .ZN(_06907_ ) );
NOR2_X1 _14931_ ( .A1(_06783_ ), .A2(_02694_ ), .ZN(_06908_ ) );
INV_X1 _14932_ ( .A(_06908_ ), .ZN(_06909_ ) );
OAI211_X1 _14933_ ( .A(_06797_ ), .B(_06909_ ), .C1(_02417_ ), .C2(_06664_ ), .ZN(_06910_ ) );
NOR2_X1 _14934_ ( .A1(_06783_ ), .A2(_04075_ ), .ZN(_06911_ ) );
INV_X1 _14935_ ( .A(_06911_ ), .ZN(_06912_ ) );
AOI21_X1 _14936_ ( .A(_02718_ ), .B1(_06778_ ), .B2(_06779_ ), .ZN(_06913_ ) );
INV_X1 _14937_ ( .A(_06913_ ), .ZN(_06914_ ) );
NAND4_X1 _14938_ ( .A1(_06912_ ), .A2(_06914_ ), .A3(_06689_ ), .A4(_06690_ ), .ZN(_06915_ ) );
AND3_X1 _14939_ ( .A1(_06910_ ), .A2(_06676_ ), .A3(_06915_ ), .ZN(_06916_ ) );
NOR2_X1 _14940_ ( .A1(_06672_ ), .A2(_02370_ ), .ZN(_06917_ ) );
OAI21_X1 _14941_ ( .A(_06797_ ), .B1(_06885_ ), .B2(_06917_ ), .ZN(_06918_ ) );
NOR2_X1 _14942_ ( .A1(_06672_ ), .A2(_02394_ ), .ZN(_06919_ ) );
AOI21_X1 _14943_ ( .A(_02346_ ), .B1(_06778_ ), .B2(_06779_ ), .ZN(_06920_ ) );
OAI211_X1 _14944_ ( .A(_06888_ ), .B(_06889_ ), .C1(_06919_ ), .C2(_06920_ ), .ZN(_06921_ ) );
AOI21_X1 _14945_ ( .A(_06676_ ), .B1(_06918_ ), .B2(_06921_ ), .ZN(_06922_ ) );
OR3_X1 _14946_ ( .A1(_06916_ ), .A2(_06813_ ), .A3(_06922_ ), .ZN(_06923_ ) );
NOR2_X1 _14947_ ( .A1(_06666_ ), .A2(_02812_ ), .ZN(_06924_ ) );
AOI21_X1 _14948_ ( .A(_02742_ ), .B1(_06685_ ), .B2(_06686_ ), .ZN(_06925_ ) );
NOR2_X1 _14949_ ( .A1(_06924_ ), .A2(_06925_ ), .ZN(_06926_ ) );
NAND3_X1 _14950_ ( .A1(_06926_ ), .A2(_06819_ ), .A3(_06820_ ), .ZN(_06927_ ) );
NOR2_X1 _14951_ ( .A1(_06768_ ), .A2(_02765_ ), .ZN(_06928_ ) );
INV_X1 _14952_ ( .A(_06928_ ), .ZN(_06929_ ) );
AOI21_X1 _14953_ ( .A(_02647_ ), .B1(_06792_ ), .B2(_06793_ ), .ZN(_06930_ ) );
INV_X1 _14954_ ( .A(_06930_ ), .ZN(_06931_ ) );
NAND3_X1 _14955_ ( .A1(_06815_ ), .A2(_06929_ ), .A3(_06931_ ), .ZN(_06932_ ) );
AOI21_X1 _14956_ ( .A(_06682_ ), .B1(_06927_ ), .B2(_06932_ ), .ZN(_06933_ ) );
AOI21_X1 _14957_ ( .A(_02789_ ), .B1(_06685_ ), .B2(_06686_ ), .ZN(_06934_ ) );
NOR2_X1 _14958_ ( .A1(_06672_ ), .A2(_02543_ ), .ZN(_06935_ ) );
OAI21_X1 _14959_ ( .A(_06815_ ), .B1(_06934_ ), .B2(_06935_ ), .ZN(_06936_ ) );
NOR2_X1 _14960_ ( .A1(_06768_ ), .A2(_02589_ ), .ZN(_06937_ ) );
AOI21_X1 _14961_ ( .A(_02565_ ), .B1(_06792_ ), .B2(_06793_ ), .ZN(_06938_ ) );
OAI211_X1 _14962_ ( .A(_06819_ ), .B(_06820_ ), .C1(_06937_ ), .C2(_06938_ ), .ZN(_06939_ ) );
AND3_X1 _14963_ ( .A1(_06936_ ), .A2(_06682_ ), .A3(_06939_ ), .ZN(_06940_ ) );
OAI21_X1 _14964_ ( .A(_06814_ ), .B1(_06933_ ), .B2(_06940_ ), .ZN(_06941_ ) );
AOI21_X1 _14965_ ( .A(_06876_ ), .B1(_06923_ ), .B2(_06941_ ), .ZN(_06942_ ) );
BUF_X2 _14966_ ( .A(_06706_ ), .Z(_06943_ ) );
AOI21_X1 _14967_ ( .A(_02611_ ), .B1(_06792_ ), .B2(_06793_ ), .ZN(_06944_ ) );
NOR2_X1 _14968_ ( .A1(_06783_ ), .A2(_02516_ ), .ZN(_06945_ ) );
AOI211_X1 _14969_ ( .A(_06944_ ), .B(_06945_ ), .C1(_06888_ ), .C2(_06889_ ), .ZN(_06946_ ) );
AOI21_X1 _14970_ ( .A(_02441_ ), .B1(_06792_ ), .B2(_06793_ ), .ZN(_06947_ ) );
NOR2_X1 _14971_ ( .A1(_06768_ ), .A2(_02464_ ), .ZN(_06948_ ) );
NOR3_X1 _14972_ ( .A1(_06797_ ), .A2(_06947_ ), .A3(_06948_ ), .ZN(_06949_ ) );
OAI21_X1 _14973_ ( .A(_06818_ ), .B1(_06946_ ), .B2(_06949_ ), .ZN(_06950_ ) );
BUF_X4 _14974_ ( .A(_06797_ ), .Z(_06951_ ) );
AND2_X1 _14975_ ( .A1(_04331_ ), .A2(_06768_ ), .ZN(_06952_ ) );
NAND3_X1 _14976_ ( .A1(_06951_ ), .A2(_06676_ ), .A3(_06952_ ), .ZN(_06953_ ) );
AOI211_X1 _14977_ ( .A(_06943_ ), .B(_06814_ ), .C1(_06950_ ), .C2(_06953_ ), .ZN(_06954_ ) );
OAI21_X1 _14978_ ( .A(_05099_ ), .B1(_06942_ ), .B2(_06954_ ), .ZN(_06955_ ) );
NAND3_X1 _14979_ ( .A1(_04952_ ), .A2(_06244_ ), .A3(_04953_ ), .ZN(_06956_ ) );
NAND3_X1 _14980_ ( .A1(_06659_ ), .A2(_06956_ ), .A3(_05025_ ), .ZN(_06957_ ) );
OAI211_X1 _14981_ ( .A(_06955_ ), .B(_06957_ ), .C1(_06659_ ), .C2(_06843_ ), .ZN(_06958_ ) );
BUF_X4 _14982_ ( .A(_04770_ ), .Z(_06959_ ) );
AOI221_X4 _14983_ ( .A(_06958_ ), .B1(_06956_ ), .B2(_06959_ ), .C1(_06711_ ), .C2(_06903_ ), .ZN(_06960_ ) );
NAND3_X1 _14984_ ( .A1(_06904_ ), .A2(_06907_ ), .A3(_06960_ ), .ZN(_06961_ ) );
AOI21_X1 _14985_ ( .A(_06864_ ), .B1(_06961_ ), .B2(_06853_ ), .ZN(_06962_ ) );
OAI21_X1 _14986_ ( .A(_06855_ ), .B1(_05350_ ), .B2(_05407_ ), .ZN(_06963_ ) );
OAI21_X1 _14987_ ( .A(_06857_ ), .B1(_06962_ ), .B2(_06963_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_11_D ) );
OAI21_X1 _14988_ ( .A(_06288_ ), .B1(_05388_ ), .B2(_05389_ ), .ZN(_06964_ ) );
OAI22_X1 _14989_ ( .A1(_05396_ ), .A2(_06561_ ), .B1(_02371_ ), .B2(_06566_ ), .ZN(_06965_ ) );
AND2_X1 _14990_ ( .A1(_04381_ ), .A2(_02346_ ), .ZN(_06966_ ) );
INV_X1 _14991_ ( .A(_04460_ ), .ZN(_06967_ ) );
AOI21_X1 _14992_ ( .A(_06967_ ), .B1(_05043_ ), .B2(_05058_ ), .ZN(_06968_ ) );
NOR2_X1 _14993_ ( .A1(_06968_ ), .A2(_05077_ ), .ZN(_06969_ ) );
NOR2_X1 _14994_ ( .A1(_04429_ ), .A2(_02394_ ), .ZN(_06970_ ) );
OAI21_X1 _14995_ ( .A(_05080_ ), .B1(_06969_ ), .B2(_06970_ ), .ZN(_06971_ ) );
AOI21_X1 _14996_ ( .A(_06966_ ), .B1(_06971_ ), .B2(_04382_ ), .ZN(_06972_ ) );
XNOR2_X1 _14997_ ( .A(_06972_ ), .B(_04406_ ), .ZN(_06973_ ) );
BUF_X4 _14998_ ( .A(_06574_ ), .Z(_06974_ ) );
AOI21_X1 _14999_ ( .A(_06965_ ), .B1(_06973_ ), .B2(_06974_ ), .ZN(_06975_ ) );
OAI21_X1 _15000_ ( .A(_05928_ ), .B1(_06975_ ), .B2(_06584_ ), .ZN(_06976_ ) );
AND2_X4 _15001_ ( .A1(_06763_ ), .A2(_06764_ ), .ZN(_06977_ ) );
NAND2_X1 _15002_ ( .A1(_06668_ ), .A2(_06777_ ), .ZN(_06978_ ) );
OAI21_X1 _15003_ ( .A(_06669_ ), .B1(_06687_ ), .B2(_06683_ ), .ZN(_06979_ ) );
NAND3_X1 _15004_ ( .A1(_06978_ ), .A2(_06790_ ), .A3(_06979_ ), .ZN(_06980_ ) );
NAND3_X1 _15005_ ( .A1(_06671_ ), .A2(_06675_ ), .A3(_06673_ ), .ZN(_06981_ ) );
NAND2_X1 _15006_ ( .A1(_06980_ ), .A2(_06981_ ), .ZN(_06982_ ) );
NAND2_X1 _15007_ ( .A1(_06982_ ), .A2(_04876_ ), .ZN(_06983_ ) );
OAI21_X1 _15008_ ( .A(_06669_ ), .B1(_06822_ ), .B2(_06816_ ), .ZN(_06984_ ) );
OAI211_X1 _15009_ ( .A(_04861_ ), .B(_04863_ ), .C1(_06695_ ), .C2(_06694_ ), .ZN(_06985_ ) );
NAND2_X1 _15010_ ( .A1(_06984_ ), .A2(_06985_ ), .ZN(_06986_ ) );
NAND2_X1 _15011_ ( .A1(_06986_ ), .A2(_06790_ ), .ZN(_06987_ ) );
OAI21_X1 _15012_ ( .A(_04872_ ), .B1(_06698_ ), .B2(_06697_ ), .ZN(_06988_ ) );
AOI21_X1 _15013_ ( .A(_02899_ ), .B1(_06685_ ), .B2(_06686_ ), .ZN(_06989_ ) );
OAI211_X1 _15014_ ( .A(_04861_ ), .B(_04863_ ), .C1(_06679_ ), .C2(_06989_ ), .ZN(_06990_ ) );
NAND2_X1 _15015_ ( .A1(_06988_ ), .A2(_06990_ ), .ZN(_06991_ ) );
NAND2_X1 _15016_ ( .A1(_06991_ ), .A2(_06675_ ), .ZN(_06992_ ) );
NAND2_X1 _15017_ ( .A1(_06987_ ), .A2(_06992_ ), .ZN(_06993_ ) );
OAI21_X1 _15018_ ( .A(_06983_ ), .B1(_06813_ ), .B2(_06993_ ), .ZN(_06994_ ) );
AND2_X1 _15019_ ( .A1(_06994_ ), .A2(_06706_ ), .ZN(_06995_ ) );
XNOR2_X1 _15020_ ( .A(_06720_ ), .B(_06790_ ), .ZN(_06996_ ) );
AND4_X1 _15021_ ( .A1(_06866_ ), .A2(_06760_ ), .A3(_06996_ ), .A4(_06762_ ), .ZN(_06997_ ) );
OR3_X1 _15022_ ( .A1(_06977_ ), .A2(_06995_ ), .A3(_06997_ ), .ZN(_06998_ ) );
AND2_X1 _15023_ ( .A1(_06998_ ), .A2(_06716_ ), .ZN(_06999_ ) );
BUF_X4 _15024_ ( .A(_06707_ ), .Z(_07000_ ) );
BUF_X2 _15025_ ( .A(_06704_ ), .Z(_07001_ ) );
NOR2_X1 _15026_ ( .A1(_06768_ ), .A2(_02565_ ), .ZN(_07002_ ) );
OAI21_X1 _15027_ ( .A(_06951_ ), .B1(_06794_ ), .B2(_07002_ ), .ZN(_07003_ ) );
BUF_X4 _15028_ ( .A(_06888_ ), .Z(_07004_ ) );
BUF_X4 _15029_ ( .A(_06889_ ), .Z(_07005_ ) );
OAI211_X1 _15030_ ( .A(_07004_ ), .B(_07005_ ), .C1(_06828_ ), .C2(_06827_ ), .ZN(_07006_ ) );
NAND2_X1 _15031_ ( .A1(_07003_ ), .A2(_07006_ ), .ZN(_07007_ ) );
BUF_X4 _15032_ ( .A(_06693_ ), .Z(_07008_ ) );
NAND2_X1 _15033_ ( .A1(_07007_ ), .A2(_07008_ ), .ZN(_07009_ ) );
NAND4_X1 _15034_ ( .A1(_06799_ ), .A2(_06801_ ), .A3(_07004_ ), .A4(_07005_ ), .ZN(_07010_ ) );
BUF_X2 _15035_ ( .A(_06767_ ), .Z(_07011_ ) );
NAND3_X1 _15036_ ( .A1(_07011_ ), .A2(_06785_ ), .A3(_06787_ ), .ZN(_07012_ ) );
BUF_X4 _15037_ ( .A(_06791_ ), .Z(_07013_ ) );
BUF_X4 _15038_ ( .A(_07013_ ), .Z(_07014_ ) );
NAND3_X1 _15039_ ( .A1(_07010_ ), .A2(_07012_ ), .A3(_07014_ ), .ZN(_07015_ ) );
AOI21_X1 _15040_ ( .A(_07001_ ), .B1(_07009_ ), .B2(_07015_ ), .ZN(_07016_ ) );
BUF_X4 _15041_ ( .A(_06951_ ), .Z(_07017_ ) );
NOR2_X1 _15042_ ( .A1(_06768_ ), .A2(_02718_ ), .ZN(_07018_ ) );
OAI21_X1 _15043_ ( .A(_07017_ ), .B1(_06809_ ), .B2(_07018_ ), .ZN(_07019_ ) );
OAI211_X1 _15044_ ( .A(_07004_ ), .B(_07005_ ), .C1(_06780_ ), .C2(_06781_ ), .ZN(_07020_ ) );
NAND3_X1 _15045_ ( .A1(_07019_ ), .A2(_07020_ ), .A3(_06677_ ), .ZN(_07021_ ) );
OAI21_X1 _15046_ ( .A(_07011_ ), .B1(_06822_ ), .B2(_06821_ ), .ZN(_07022_ ) );
OAI211_X1 _15047_ ( .A(_07004_ ), .B(_07005_ ), .C1(_06807_ ), .C2(_06806_ ), .ZN(_07023_ ) );
NAND3_X1 _15048_ ( .A1(_07022_ ), .A2(_07014_ ), .A3(_07023_ ), .ZN(_07024_ ) );
BUF_X2 _15049_ ( .A(_06703_ ), .Z(_07025_ ) );
AND3_X1 _15050_ ( .A1(_07021_ ), .A2(_07024_ ), .A3(_07025_ ), .ZN(_07026_ ) );
OAI21_X1 _15051_ ( .A(_07000_ ), .B1(_07016_ ), .B2(_07026_ ), .ZN(_07027_ ) );
OAI21_X1 _15052_ ( .A(_06951_ ), .B1(_06831_ ), .B2(_06830_ ), .ZN(_07028_ ) );
OAI21_X1 _15053_ ( .A(_07028_ ), .B1(_07011_ ), .B2(_06835_ ), .ZN(_07029_ ) );
INV_X1 _15054_ ( .A(_07029_ ), .ZN(_07030_ ) );
NAND3_X1 _15055_ ( .A1(_07030_ ), .A2(_07025_ ), .A3(_06868_ ), .ZN(_07031_ ) );
BUF_X2 _15056_ ( .A(_06877_ ), .Z(_07032_ ) );
AOI21_X1 _15057_ ( .A(_06776_ ), .B1(_07031_ ), .B2(_07032_ ), .ZN(_07033_ ) );
AOI221_X1 _15058_ ( .A(_06999_ ), .B1(_06710_ ), .B2(_06995_ ), .C1(_07027_ ), .C2(_07033_ ), .ZN(_07034_ ) );
AND2_X1 _15059_ ( .A1(_06641_ ), .A2(_06642_ ), .ZN(_07035_ ) );
OAI21_X1 _15060_ ( .A(_04964_ ), .B1(_07035_ ), .B2(_06647_ ), .ZN(_07036_ ) );
NAND2_X1 _15061_ ( .A1(_07036_ ), .A2(_06651_ ), .ZN(_07037_ ) );
AOI21_X1 _15062_ ( .A(_06905_ ), .B1(_07037_ ), .B2(_04960_ ), .ZN(_07038_ ) );
OAI21_X1 _15063_ ( .A(_07038_ ), .B1(_04960_ ), .B2(_07037_ ), .ZN(_07039_ ) );
OAI22_X1 _15064_ ( .A1(_06649_ ), .A2(_06843_ ), .B1(_06652_ ), .B2(_06713_ ), .ZN(_07040_ ) );
BUF_X4 _15065_ ( .A(_05025_ ), .Z(_07041_ ) );
BUF_X4 _15066_ ( .A(_07041_ ), .Z(_07042_ ) );
AOI21_X1 _15067_ ( .A(_07040_ ), .B1(_04960_ ), .B2(_07042_ ), .ZN(_07043_ ) );
NAND3_X1 _15068_ ( .A1(_07034_ ), .A2(_07039_ ), .A3(_07043_ ), .ZN(_07044_ ) );
AOI21_X1 _15069_ ( .A(_06976_ ), .B1(_07044_ ), .B2(_06853_ ), .ZN(_07045_ ) );
NAND2_X1 _15070_ ( .A1(_05400_ ), .A2(_05610_ ), .ZN(_07046_ ) );
NAND2_X1 _15071_ ( .A1(_07046_ ), .A2(_06214_ ), .ZN(_07047_ ) );
OAI21_X1 _15072_ ( .A(_06964_ ), .B1(_07045_ ), .B2(_07047_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_12_D ) );
OAI21_X1 _15073_ ( .A(_06288_ ), .B1(_05416_ ), .B2(_05417_ ), .ZN(_07048_ ) );
NAND2_X1 _15074_ ( .A1(_05424_ ), .A2(_03892_ ), .ZN(_07049_ ) );
NAND3_X1 _15075_ ( .A1(_06896_ ), .A2(_06693_ ), .A3(_07011_ ), .ZN(_07050_ ) );
OAI21_X1 _15076_ ( .A(_06797_ ), .B1(_06881_ ), .B2(_06882_ ), .ZN(_07051_ ) );
OAI211_X1 _15077_ ( .A(_06689_ ), .B(_06690_ ), .C1(_06897_ ), .C2(_06898_ ), .ZN(_07052_ ) );
NAND3_X1 _15078_ ( .A1(_07051_ ), .A2(_07013_ ), .A3(_07052_ ), .ZN(_07053_ ) );
AND2_X1 _15079_ ( .A1(_07050_ ), .A2(_07053_ ), .ZN(_07054_ ) );
NOR2_X1 _15080_ ( .A1(_06917_ ), .A2(_06920_ ), .ZN(_07055_ ) );
AND2_X1 _15081_ ( .A1(_07055_ ), .A2(_06815_ ), .ZN(_07056_ ) );
NOR3_X1 _15082_ ( .A1(_06815_ ), .A2(_06885_ ), .A3(_06886_ ), .ZN(_07057_ ) );
OAI21_X1 _15083_ ( .A(_06805_ ), .B1(_07056_ ), .B2(_07057_ ), .ZN(_07058_ ) );
OAI21_X1 _15084_ ( .A(_06797_ ), .B1(_06891_ ), .B2(_06890_ ), .ZN(_07059_ ) );
OAI211_X1 _15085_ ( .A(_06689_ ), .B(_06690_ ), .C1(_06879_ ), .C2(_06878_ ), .ZN(_07060_ ) );
NAND3_X1 _15086_ ( .A1(_07059_ ), .A2(_06693_ ), .A3(_07060_ ), .ZN(_07061_ ) );
AND2_X1 _15087_ ( .A1(_07058_ ), .A2(_07061_ ), .ZN(_07062_ ) );
BUF_X2 _15088_ ( .A(_06703_ ), .Z(_07063_ ) );
MUX2_X1 _15089_ ( .A(_07054_ ), .B(_07062_ ), .S(_07063_ ), .Z(_07064_ ) );
INV_X1 _15090_ ( .A(_06709_ ), .ZN(_07065_ ) );
OR3_X1 _15091_ ( .A1(_07064_ ), .A2(_07032_ ), .A3(_07065_ ), .ZN(_07066_ ) );
OR3_X1 _15092_ ( .A1(_07035_ ), .A2(_04964_ ), .A3(_06647_ ), .ZN(_07067_ ) );
AND3_X1 _15093_ ( .A1(_07067_ ), .A2(_06589_ ), .A3(_07036_ ), .ZN(_07068_ ) );
OAI21_X1 _15094_ ( .A(_06767_ ), .B1(_06947_ ), .B2(_06948_ ), .ZN(_07069_ ) );
OAI211_X1 _15095_ ( .A(_06888_ ), .B(_06889_ ), .C1(_06664_ ), .C2(_06479_ ), .ZN(_07070_ ) );
AND3_X1 _15096_ ( .A1(_07069_ ), .A2(_06805_ ), .A3(_07070_ ), .ZN(_07071_ ) );
AND2_X1 _15097_ ( .A1(_07071_ ), .A2(_07063_ ), .ZN(_07072_ ) );
OAI21_X1 _15098_ ( .A(_05099_ ), .B1(_07072_ ), .B2(_06707_ ), .ZN(_07073_ ) );
AND2_X1 _15099_ ( .A1(_06926_ ), .A2(_06669_ ), .ZN(_07074_ ) );
NOR3_X1 _15100_ ( .A1(_06669_ ), .A2(_06934_ ), .A3(_06935_ ), .ZN(_07075_ ) );
OAI21_X1 _15101_ ( .A(_06805_ ), .B1(_07074_ ), .B2(_07075_ ), .ZN(_07076_ ) );
OAI21_X1 _15102_ ( .A(_06767_ ), .B1(_06938_ ), .B2(_06937_ ), .ZN(_07077_ ) );
OAI211_X1 _15103_ ( .A(_06888_ ), .B(_06889_ ), .C1(_06945_ ), .C2(_06944_ ), .ZN(_07078_ ) );
NAND3_X1 _15104_ ( .A1(_07077_ ), .A2(_06677_ ), .A3(_07078_ ), .ZN(_07079_ ) );
AND2_X1 _15105_ ( .A1(_07076_ ), .A2(_07079_ ), .ZN(_07080_ ) );
NAND4_X1 _15106_ ( .A1(_06929_ ), .A2(_06931_ ), .A3(_06888_ ), .A4(_06889_ ), .ZN(_07081_ ) );
NAND3_X1 _15107_ ( .A1(_06767_ ), .A2(_06912_ ), .A3(_06914_ ), .ZN(_07082_ ) );
AND2_X1 _15108_ ( .A1(_07081_ ), .A2(_07082_ ), .ZN(_07083_ ) );
AOI211_X1 _15109_ ( .A(_06920_ ), .B(_06919_ ), .C1(_06689_ ), .C2(_04863_ ), .ZN(_07084_ ) );
AOI21_X1 _15110_ ( .A(_02417_ ), .B1(_06778_ ), .B2(_06779_ ), .ZN(_07085_ ) );
NOR3_X1 _15111_ ( .A1(_06671_ ), .A2(_07085_ ), .A3(_06908_ ), .ZN(_07086_ ) );
NOR2_X1 _15112_ ( .A1(_07084_ ), .A2(_07086_ ), .ZN(_07087_ ) );
MUX2_X1 _15113_ ( .A(_07083_ ), .B(_07087_ ), .S(_06805_ ), .Z(_07088_ ) );
MUX2_X1 _15114_ ( .A(_07080_ ), .B(_07088_ ), .S(_07063_ ), .Z(_07089_ ) );
AOI21_X1 _15115_ ( .A(_07073_ ), .B1(_07089_ ), .B2(_07000_ ), .ZN(_07090_ ) );
NOR2_X1 _15116_ ( .A1(_07068_ ), .A2(_07090_ ), .ZN(_07091_ ) );
BUF_X4 _15117_ ( .A(_06586_ ), .Z(_07092_ ) );
NAND3_X1 _15118_ ( .A1(_04991_ ), .A2(_02346_ ), .A3(_07092_ ), .ZN(_07093_ ) );
NAND3_X1 _15119_ ( .A1(_04961_ ), .A2(_04357_ ), .A3(_04962_ ), .ZN(_07094_ ) );
AOI22_X1 _15120_ ( .A1(_04964_ ), .A2(_07042_ ), .B1(_07094_ ), .B2(_06959_ ), .ZN(_07095_ ) );
AND4_X1 _15121_ ( .A1(_07066_ ), .A2(_07091_ ), .A3(_07093_ ), .A4(_07095_ ), .ZN(_07096_ ) );
BUF_X4 _15122_ ( .A(_06760_ ), .Z(_07097_ ) );
AND2_X1 _15123_ ( .A1(_04872_ ), .A2(_06663_ ), .ZN(_07098_ ) );
INV_X1 _15124_ ( .A(_07098_ ), .ZN(_07099_ ) );
NAND4_X1 _15125_ ( .A1(_07097_ ), .A2(_07099_ ), .A3(_06867_ ), .A4(_06996_ ), .ZN(_07100_ ) );
AOI22_X1 _15126_ ( .A1(_06873_ ), .A2(_06874_ ), .B1(_06872_ ), .B2(_07100_ ), .ZN(_07101_ ) );
NOR2_X1 _15127_ ( .A1(_07064_ ), .A2(_07032_ ), .ZN(_07102_ ) );
OAI21_X1 _15128_ ( .A(_06865_ ), .B1(_07101_ ), .B2(_07102_ ), .ZN(_07103_ ) );
AOI21_X1 _15129_ ( .A(_06851_ ), .B1(_07096_ ), .B2(_07103_ ), .ZN(_07104_ ) );
XNOR2_X1 _15130_ ( .A(_06971_ ), .B(_04382_ ), .ZN(_07105_ ) );
NOR2_X1 _15131_ ( .A1(_07105_ ), .A2(_06576_ ), .ZN(_07106_ ) );
OAI22_X1 _15132_ ( .A1(_05422_ ), .A2(_06861_ ), .B1(_02347_ ), .B2(_06566_ ), .ZN(_07107_ ) );
OAI21_X1 _15133_ ( .A(_06582_ ), .B1(_07106_ ), .B2(_07107_ ), .ZN(_07108_ ) );
NAND2_X1 _15134_ ( .A1(_07108_ ), .A2(_05347_ ), .ZN(_07109_ ) );
OAI21_X1 _15135_ ( .A(_07049_ ), .B1(_07104_ ), .B2(_07109_ ), .ZN(_07110_ ) );
OAI21_X1 _15136_ ( .A(_07048_ ), .B1(_07110_ ), .B2(_06393_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_13_D ) );
NAND3_X1 _15137_ ( .A1(_05445_ ), .A2(_05447_ ), .A3(_06556_ ), .ZN(_07111_ ) );
OAI22_X1 _15138_ ( .A1(_05433_ ), .A2(_06561_ ), .B1(_02395_ ), .B2(_06565_ ), .ZN(_07112_ ) );
XNOR2_X1 _15139_ ( .A(_06969_ ), .B(_04431_ ), .ZN(_07113_ ) );
AOI21_X1 _15140_ ( .A(_07112_ ), .B1(_07113_ ), .B2(_06974_ ), .ZN(_07114_ ) );
OAI21_X1 _15141_ ( .A(_05928_ ), .B1(_07114_ ), .B2(_06584_ ), .ZN(_07115_ ) );
AND3_X1 _15142_ ( .A1(_06760_ ), .A2(_06867_ ), .A3(_06996_ ), .ZN(_07116_ ) );
NAND2_X1 _15143_ ( .A1(_07116_ ), .A2(_06769_ ), .ZN(_07117_ ) );
AOI22_X1 _15144_ ( .A1(_07117_ ), .A2(_06872_ ), .B1(_06873_ ), .B2(_06874_ ), .ZN(_07118_ ) );
NAND2_X1 _15145_ ( .A1(_06674_ ), .A2(_06676_ ), .ZN(_07119_ ) );
NAND3_X1 _15146_ ( .A1(_06681_ ), .A2(_06790_ ), .A3(_06691_ ), .ZN(_07120_ ) );
NAND3_X1 _15147_ ( .A1(_07119_ ), .A2(_06813_ ), .A3(_07120_ ), .ZN(_07121_ ) );
OAI21_X1 _15148_ ( .A(_06669_ ), .B1(_06806_ ), .B2(_06821_ ), .ZN(_07122_ ) );
OAI211_X1 _15149_ ( .A(_04861_ ), .B(_04863_ ), .C1(_06816_ ), .C2(_06822_ ), .ZN(_07123_ ) );
AOI21_X1 _15150_ ( .A(_06675_ ), .B1(_07122_ ), .B2(_07123_ ), .ZN(_07124_ ) );
AOI21_X1 _15151_ ( .A(_06790_ ), .B1(_06696_ ), .B2(_06699_ ), .ZN(_07125_ ) );
OR2_X1 _15152_ ( .A1(_07124_ ), .A2(_07125_ ), .ZN(_07126_ ) );
OAI21_X1 _15153_ ( .A(_07121_ ), .B1(_06813_ ), .B2(_07126_ ), .ZN(_07127_ ) );
AND2_X1 _15154_ ( .A1(_07127_ ), .A2(_06708_ ), .ZN(_07128_ ) );
OAI21_X1 _15155_ ( .A(_06865_ ), .B1(_07118_ ), .B2(_07128_ ), .ZN(_07129_ ) );
NAND2_X1 _15156_ ( .A1(_06641_ ), .A2(_04972_ ), .ZN(_07130_ ) );
INV_X1 _15157_ ( .A(_06645_ ), .ZN(_07131_ ) );
NAND2_X1 _15158_ ( .A1(_07130_ ), .A2(_07131_ ), .ZN(_07132_ ) );
AOI21_X1 _15159_ ( .A(_06905_ ), .B1(_07132_ ), .B2(_04968_ ), .ZN(_07133_ ) );
OAI21_X1 _15160_ ( .A(_07133_ ), .B1(_04968_ ), .B2(_07132_ ), .ZN(_07134_ ) );
BUF_X4 _15161_ ( .A(_06813_ ), .Z(_07135_ ) );
AND3_X1 _15162_ ( .A1(_06796_ ), .A2(_06802_ ), .A3(_06791_ ), .ZN(_07136_ ) );
AOI21_X1 _15163_ ( .A(_06791_ ), .B1(_06829_ ), .B2(_06832_ ), .ZN(_07137_ ) );
OAI21_X1 _15164_ ( .A(_07135_ ), .B1(_07136_ ), .B2(_07137_ ), .ZN(_07138_ ) );
NAND3_X1 _15165_ ( .A1(_06808_ ), .A2(_06791_ ), .A3(_06811_ ), .ZN(_07139_ ) );
NAND3_X1 _15166_ ( .A1(_06782_ ), .A2(_06676_ ), .A3(_06788_ ), .ZN(_07140_ ) );
AND2_X1 _15167_ ( .A1(_07139_ ), .A2(_07140_ ), .ZN(_07141_ ) );
OAI211_X1 _15168_ ( .A(_06943_ ), .B(_07138_ ), .C1(_07141_ ), .C2(_07135_ ), .ZN(_07142_ ) );
AND3_X1 _15169_ ( .A1(_06835_ ), .A2(_07013_ ), .A3(_07011_ ), .ZN(_07143_ ) );
NAND3_X1 _15170_ ( .A1(_07143_ ), .A2(_06876_ ), .A3(_06703_ ), .ZN(_07144_ ) );
AOI21_X1 _15171_ ( .A(_06776_ ), .B1(_07142_ ), .B2(_07144_ ), .ZN(_07145_ ) );
AOI21_X1 _15172_ ( .A(_04771_ ), .B1(_04967_ ), .B2(_04430_ ), .ZN(_07146_ ) );
AND3_X1 _15173_ ( .A1(_07127_ ), .A2(_06943_ ), .A3(_06709_ ), .ZN(_07147_ ) );
OR3_X1 _15174_ ( .A1(_07145_ ), .A2(_07146_ ), .A3(_07147_ ), .ZN(_07148_ ) );
AOI221_X4 _15175_ ( .A(_07148_ ), .B1(_06644_ ), .B2(_07092_ ), .C1(_04968_ ), .C2(_07042_ ), .ZN(_07149_ ) );
NAND3_X1 _15176_ ( .A1(_07129_ ), .A2(_07134_ ), .A3(_07149_ ), .ZN(_07150_ ) );
AOI21_X1 _15177_ ( .A(_07115_ ), .B1(_07150_ ), .B2(_06853_ ), .ZN(_07151_ ) );
NAND2_X1 _15178_ ( .A1(_05430_ ), .A2(_05610_ ), .ZN(_07152_ ) );
NAND2_X1 _15179_ ( .A1(_07152_ ), .A2(_06422_ ), .ZN(_07153_ ) );
OAI21_X1 _15180_ ( .A(_07111_ ), .B1(_07151_ ), .B2(_07153_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_14_D ) );
AND2_X1 _15181_ ( .A1(_05459_ ), .A2(_05460_ ), .ZN(_07154_ ) );
AND2_X1 _15182_ ( .A1(_05468_ ), .A2(_05470_ ), .ZN(_07155_ ) );
NAND4_X1 _15183_ ( .A1(_05293_ ), .A2(_07154_ ), .A3(_07155_ ), .A4(_05444_ ), .ZN(_07156_ ) );
NAND3_X1 _15184_ ( .A1(_05840_ ), .A2(_05841_ ), .A3(_06124_ ), .ZN(_07157_ ) );
NAND3_X1 _15185_ ( .A1(_07156_ ), .A2(_07157_ ), .A3(_06556_ ), .ZN(_07158_ ) );
OAI21_X1 _15186_ ( .A(_06858_ ), .B1(_05059_ ), .B2(_06967_ ), .ZN(_07159_ ) );
AOI21_X1 _15187_ ( .A(_07159_ ), .B1(_06967_ ), .B2(_05059_ ), .ZN(_07160_ ) );
OAI22_X1 _15188_ ( .A1(_05457_ ), .A2(_06861_ ), .B1(_02418_ ), .B2(_06566_ ), .ZN(_07161_ ) );
OAI21_X1 _15189_ ( .A(_06582_ ), .B1(_07160_ ), .B2(_07161_ ), .ZN(_07162_ ) );
NAND2_X1 _15190_ ( .A1(_07162_ ), .A2(_05347_ ), .ZN(_07163_ ) );
INV_X1 _15191_ ( .A(_06722_ ), .ZN(_07164_ ) );
AOI21_X1 _15192_ ( .A(_06873_ ), .B1(_06708_ ), .B2(_07164_ ), .ZN(_07165_ ) );
OR3_X1 _15193_ ( .A1(_06777_ ), .A2(_07085_ ), .A3(_06919_ ), .ZN(_07166_ ) );
NAND3_X1 _15194_ ( .A1(_07055_ ), .A2(_06819_ ), .A3(_06820_ ), .ZN(_07167_ ) );
AND3_X1 _15195_ ( .A1(_07166_ ), .A2(_06818_ ), .A3(_07167_ ), .ZN(_07168_ ) );
AOI21_X1 _15196_ ( .A(_06818_ ), .B1(_06887_ ), .B2(_06892_ ), .ZN(_07169_ ) );
OR3_X1 _15197_ ( .A1(_07168_ ), .A2(_07135_ ), .A3(_07169_ ), .ZN(_07170_ ) );
OR3_X1 _15198_ ( .A1(_06880_ ), .A2(_06883_ ), .A3(_06675_ ), .ZN(_07171_ ) );
OAI21_X1 _15199_ ( .A(_07171_ ), .B1(_06900_ ), .B2(_07013_ ), .ZN(_07172_ ) );
OAI21_X1 _15200_ ( .A(_07170_ ), .B1(_07172_ ), .B2(_07063_ ), .ZN(_07173_ ) );
BUF_X2 _15201_ ( .A(_06943_ ), .Z(_07174_ ) );
AND2_X1 _15202_ ( .A1(_07173_ ), .A2(_07174_ ), .ZN(_07175_ ) );
OAI21_X1 _15203_ ( .A(_06865_ ), .B1(_07165_ ), .B2(_07175_ ), .ZN(_07176_ ) );
AOI21_X1 _15204_ ( .A(_06905_ ), .B1(_06641_ ), .B2(_04972_ ), .ZN(_07177_ ) );
OAI21_X1 _15205_ ( .A(_07177_ ), .B1(_04972_ ), .B2(_06641_ ), .ZN(_07178_ ) );
NAND3_X1 _15206_ ( .A1(_06927_ ), .A2(_06682_ ), .A3(_06932_ ), .ZN(_07179_ ) );
NAND3_X1 _15207_ ( .A1(_06910_ ), .A2(_06818_ ), .A3(_06915_ ), .ZN(_07180_ ) );
AOI21_X1 _15208_ ( .A(_07135_ ), .B1(_07179_ ), .B2(_07180_ ), .ZN(_07181_ ) );
OAI21_X1 _15209_ ( .A(_06682_ ), .B1(_06946_ ), .B2(_06949_ ), .ZN(_07182_ ) );
NAND3_X1 _15210_ ( .A1(_06936_ ), .A2(_07013_ ), .A3(_06939_ ), .ZN(_07183_ ) );
AND2_X1 _15211_ ( .A1(_07182_ ), .A2(_07183_ ), .ZN(_07184_ ) );
AOI211_X1 _15212_ ( .A(_06876_ ), .B(_07181_ ), .C1(_07184_ ), .C2(_06839_ ), .ZN(_07185_ ) );
AND3_X1 _15213_ ( .A1(_07011_ ), .A2(_07013_ ), .A3(_06952_ ), .ZN(_07186_ ) );
AND3_X1 _15214_ ( .A1(_07186_ ), .A2(_06876_ ), .A3(_06703_ ), .ZN(_07187_ ) );
OAI21_X1 _15215_ ( .A(_05099_ ), .B1(_07185_ ), .B2(_07187_ ), .ZN(_07188_ ) );
NAND3_X1 _15216_ ( .A1(_04969_ ), .A2(_04432_ ), .A3(_04970_ ), .ZN(_07189_ ) );
NAND3_X1 _15217_ ( .A1(_07131_ ), .A2(_07189_ ), .A3(_05025_ ), .ZN(_07190_ ) );
OAI211_X1 _15218_ ( .A(_07188_ ), .B(_07190_ ), .C1(_07131_ ), .C2(_06843_ ), .ZN(_07191_ ) );
AOI221_X4 _15219_ ( .A(_07191_ ), .B1(_07189_ ), .B2(_06959_ ), .C1(_06711_ ), .C2(_07175_ ), .ZN(_07192_ ) );
NAND3_X1 _15220_ ( .A1(_07176_ ), .A2(_07178_ ), .A3(_07192_ ), .ZN(_07193_ ) );
AOI21_X1 _15221_ ( .A(_07163_ ), .B1(_07193_ ), .B2(_06853_ ), .ZN(_07194_ ) );
OAI21_X1 _15222_ ( .A(_06855_ ), .B1(_05454_ ), .B2(_05407_ ), .ZN(_07195_ ) );
OAI21_X1 _15223_ ( .A(_07158_ ), .B1(_07194_ ), .B2(_07195_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_15_D ) );
OAI21_X1 _15224_ ( .A(_06288_ ), .B1(_05498_ ), .B2(_05499_ ), .ZN(_07196_ ) );
BUF_X4 _15225_ ( .A(_06583_ ), .Z(_07197_ ) );
OAI21_X1 _15226_ ( .A(_05056_ ), .B1(_05041_ ), .B2(_04050_ ), .ZN(_07198_ ) );
AND2_X1 _15227_ ( .A1(_07198_ ), .A2(_04108_ ), .ZN(_07199_ ) );
OAI21_X1 _15228_ ( .A(_04165_ ), .B1(_07199_ ), .B2(_05047_ ), .ZN(_07200_ ) );
NAND2_X1 _15229_ ( .A1(_04164_ ), .A2(_02718_ ), .ZN(_07201_ ) );
AND2_X1 _15230_ ( .A1(_07200_ ), .A2(_07201_ ), .ZN(_07202_ ) );
XNOR2_X1 _15231_ ( .A(_07202_ ), .B(_04133_ ), .ZN(_07203_ ) );
NAND2_X1 _15232_ ( .A1(_07203_ ), .A2(_06974_ ), .ZN(_07204_ ) );
BUF_X2 _15233_ ( .A(_06560_ ), .Z(_07205_ ) );
BUF_X4 _15234_ ( .A(_06564_ ), .Z(_07206_ ) );
AOI22_X1 _15235_ ( .A1(_05485_ ), .A2(_07205_ ), .B1(\ID_EX_imm [15] ), .B2(_07206_ ), .ZN(_07207_ ) );
AOI21_X1 _15236_ ( .A(_07197_ ), .B1(_07204_ ), .B2(_07207_ ), .ZN(_07208_ ) );
OR2_X1 _15237_ ( .A1(_07208_ ), .A2(_03892_ ), .ZN(_07209_ ) );
AND2_X1 _15238_ ( .A1(_04831_ ), .A2(_06315_ ), .ZN(_07210_ ) );
AND2_X1 _15239_ ( .A1(_06638_ ), .A2(_06595_ ), .ZN(_07211_ ) );
INV_X1 _15240_ ( .A(_07211_ ), .ZN(_07212_ ) );
AOI21_X1 _15241_ ( .A(_04838_ ), .B1(_07212_ ), .B2(_06601_ ), .ZN(_07213_ ) );
INV_X1 _15242_ ( .A(_07213_ ), .ZN(_07214_ ) );
INV_X1 _15243_ ( .A(_06610_ ), .ZN(_07215_ ) );
AOI21_X1 _15244_ ( .A(_07210_ ), .B1(_07214_ ), .B2(_07215_ ), .ZN(_07216_ ) );
NOR2_X1 _15245_ ( .A1(_07216_ ), .A2(_06609_ ), .ZN(_07217_ ) );
NOR2_X1 _15246_ ( .A1(_07217_ ), .A2(_06608_ ), .ZN(_07218_ ) );
INV_X1 _15247_ ( .A(_07218_ ), .ZN(_07219_ ) );
NAND3_X1 _15248_ ( .A1(_07219_ ), .A2(_04931_ ), .A3(_04826_ ), .ZN(_07220_ ) );
BUF_X2 _15249_ ( .A(_06589_ ), .Z(_07221_ ) );
OAI21_X1 _15250_ ( .A(_04821_ ), .B1(_07218_ ), .B2(_04825_ ), .ZN(_07222_ ) );
NAND3_X1 _15251_ ( .A1(_07220_ ), .A2(_07221_ ), .A3(_07222_ ), .ZN(_07223_ ) );
NAND4_X1 _15252_ ( .A1(_07097_ ), .A2(_06865_ ), .A3(_06766_ ), .A4(_06762_ ), .ZN(_07224_ ) );
AOI21_X1 _15253_ ( .A(_06818_ ), .B1(_06978_ ), .B2(_06979_ ), .ZN(_07225_ ) );
AOI21_X1 _15254_ ( .A(_06676_ ), .B1(_06988_ ), .B2(_06990_ ), .ZN(_07226_ ) );
OR3_X1 _15255_ ( .A1(_07225_ ), .A2(_07063_ ), .A3(_07226_ ), .ZN(_07227_ ) );
BUF_X4 _15256_ ( .A(_07135_ ), .Z(_07228_ ) );
BUF_X2 _15257_ ( .A(_07228_ ), .Z(_07229_ ) );
OAI21_X1 _15258_ ( .A(_06767_ ), .B1(_06809_ ), .B2(_06807_ ), .ZN(_07230_ ) );
OAI211_X1 _15259_ ( .A(_06888_ ), .B(_06889_ ), .C1(_06821_ ), .C2(_06806_ ), .ZN(_07231_ ) );
NAND2_X1 _15260_ ( .A1(_07230_ ), .A2(_07231_ ), .ZN(_07232_ ) );
MUX2_X1 _15261_ ( .A(_07232_ ), .B(_06986_ ), .S(_06682_ ), .Z(_07233_ ) );
OAI211_X1 _15262_ ( .A(_07227_ ), .B(_07000_ ), .C1(_07229_ ), .C2(_07233_ ), .ZN(_07234_ ) );
NAND3_X1 _15263_ ( .A1(_07017_ ), .A2(_07014_ ), .A3(_06673_ ), .ZN(_07235_ ) );
OAI21_X1 _15264_ ( .A(_07032_ ), .B1(_07235_ ), .B2(_07229_ ), .ZN(_07236_ ) );
AND2_X1 _15265_ ( .A1(\ID_EX_typ [2] ), .A2(\ID_EX_typ [1] ), .ZN(_07237_ ) );
NAND3_X1 _15266_ ( .A1(_07234_ ), .A2(_07236_ ), .A3(_07237_ ), .ZN(_07238_ ) );
OR3_X1 _15267_ ( .A1(_04820_ ), .A2(_04109_ ), .A3(_06843_ ), .ZN(_07239_ ) );
AOI21_X1 _15268_ ( .A(_06713_ ), .B1(_04820_ ), .B2(_04109_ ), .ZN(_07240_ ) );
AOI21_X1 _15269_ ( .A(_07240_ ), .B1(_04821_ ), .B2(_07042_ ), .ZN(_07241_ ) );
MUX2_X1 _15270_ ( .A(_07007_ ), .B(_07029_ ), .S(_06677_ ), .Z(_07242_ ) );
NAND2_X1 _15271_ ( .A1(_07242_ ), .A2(_07229_ ), .ZN(_07243_ ) );
AND3_X1 _15272_ ( .A1(_07010_ ), .A2(_07012_ ), .A3(_06677_ ), .ZN(_07244_ ) );
AOI21_X1 _15273_ ( .A(_07008_ ), .B1(_07019_ ), .B2(_07020_ ), .ZN(_07245_ ) );
OAI21_X1 _15274_ ( .A(_07001_ ), .B1(_07244_ ), .B2(_07245_ ), .ZN(_07246_ ) );
AND2_X1 _15275_ ( .A1(_06706_ ), .A2(_05099_ ), .ZN(_07247_ ) );
BUF_X2 _15276_ ( .A(_07247_ ), .Z(_07248_ ) );
NAND3_X1 _15277_ ( .A1(_07243_ ), .A2(_07246_ ), .A3(_07248_ ), .ZN(_07249_ ) );
AND4_X1 _15278_ ( .A1(_07238_ ), .A2(_07239_ ), .A3(_07241_ ), .A4(_07249_ ), .ZN(_07250_ ) );
NAND3_X1 _15279_ ( .A1(_07223_ ), .A2(_07224_ ), .A3(_07250_ ), .ZN(_07251_ ) );
AOI21_X1 _15280_ ( .A(_07209_ ), .B1(_07251_ ), .B2(_06853_ ), .ZN(_07252_ ) );
NAND2_X1 _15281_ ( .A1(_05488_ ), .A2(_05610_ ), .ZN(_07253_ ) );
NAND2_X1 _15282_ ( .A1(_07253_ ), .A2(_06422_ ), .ZN(_07254_ ) );
OAI21_X1 _15283_ ( .A(_07196_ ), .B1(_07252_ ), .B2(_07254_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_16_D ) );
AND2_X1 _15284_ ( .A1(_05511_ ), .A2(_05512_ ), .ZN(_07255_ ) );
AND2_X1 _15285_ ( .A1(_05514_ ), .A2(_05515_ ), .ZN(_07256_ ) );
NAND4_X1 _15286_ ( .A1(_05293_ ), .A2(_07255_ ), .A3(_07256_ ), .A4(_05444_ ), .ZN(_07257_ ) );
NAND3_X1 _15287_ ( .A1(_05840_ ), .A2(_05841_ ), .A3(_06134_ ), .ZN(_07258_ ) );
NAND3_X1 _15288_ ( .A1(_07257_ ), .A2(_07258_ ), .A3(_06556_ ), .ZN(_07259_ ) );
OR3_X1 _15289_ ( .A1(_07199_ ), .A2(_04165_ ), .A3(_05047_ ), .ZN(_07260_ ) );
NAND3_X1 _15290_ ( .A1(_07260_ ), .A2(_06858_ ), .A3(_07200_ ), .ZN(_07261_ ) );
AOI22_X1 _15291_ ( .A1(_05508_ ), .A2(_07205_ ), .B1(\ID_EX_imm [14] ), .B2(_07206_ ), .ZN(_07262_ ) );
AOI21_X1 _15292_ ( .A(_07197_ ), .B1(_07261_ ), .B2(_07262_ ), .ZN(_07263_ ) );
OR2_X1 _15293_ ( .A1(_07263_ ), .A2(_05609_ ), .ZN(_07264_ ) );
AND2_X1 _15294_ ( .A1(_07098_ ), .A2(_04880_ ), .ZN(_07265_ ) );
AND2_X1 _15295_ ( .A1(_06771_ ), .A2(_07265_ ), .ZN(_07266_ ) );
OR3_X1 _15296_ ( .A1(_06873_ ), .A2(_06872_ ), .A3(_07266_ ), .ZN(_07267_ ) );
AOI21_X1 _15297_ ( .A(_06675_ ), .B1(_07059_ ), .B2(_07060_ ), .ZN(_07268_ ) );
AOI21_X1 _15298_ ( .A(_06790_ ), .B1(_07051_ ), .B2(_07052_ ), .ZN(_07269_ ) );
NOR2_X1 _15299_ ( .A1(_07268_ ), .A2(_07269_ ), .ZN(_07270_ ) );
OAI21_X1 _15300_ ( .A(_06693_ ), .B1(_07056_ ), .B2(_07057_ ), .ZN(_07271_ ) );
OAI21_X1 _15301_ ( .A(_06951_ ), .B1(_06913_ ), .B2(_06908_ ), .ZN(_07272_ ) );
OAI211_X1 _15302_ ( .A(_07004_ ), .B(_07005_ ), .C1(_06919_ ), .C2(_07085_ ), .ZN(_07273_ ) );
NAND3_X1 _15303_ ( .A1(_07272_ ), .A2(_07013_ ), .A3(_07273_ ), .ZN(_07274_ ) );
NAND2_X1 _15304_ ( .A1(_07271_ ), .A2(_07274_ ), .ZN(_07275_ ) );
MUX2_X1 _15305_ ( .A(_07270_ ), .B(_07275_ ), .S(_06704_ ), .Z(_07276_ ) );
AND2_X1 _15306_ ( .A1(_07276_ ), .A2(_07174_ ), .ZN(_07277_ ) );
AND3_X1 _15307_ ( .A1(_06896_ ), .A2(_04880_ ), .A3(_06669_ ), .ZN(_07278_ ) );
AND3_X1 _15308_ ( .A1(_07278_ ), .A2(_06877_ ), .A3(_07025_ ), .ZN(_07279_ ) );
NOR2_X1 _15309_ ( .A1(_07277_ ), .A2(_07279_ ), .ZN(_07280_ ) );
AOI21_X1 _15310_ ( .A(_06718_ ), .B1(_07267_ ), .B2(_07280_ ), .ZN(_07281_ ) );
OAI21_X1 _15311_ ( .A(_06589_ ), .B1(_07217_ ), .B2(_06608_ ), .ZN(_07282_ ) );
AOI21_X1 _15312_ ( .A(_07282_ ), .B1(_06608_ ), .B2(_07217_ ), .ZN(_07283_ ) );
OAI21_X1 _15313_ ( .A(_06710_ ), .B1(_07277_ ), .B2(_07279_ ), .ZN(_07284_ ) );
OR3_X1 _15314_ ( .A1(_04824_ ), .A2(_04134_ ), .A3(_06843_ ), .ZN(_07285_ ) );
AOI22_X1 _15315_ ( .A1(_06603_ ), .A2(_07041_ ), .B1(_04827_ ), .B2(_04770_ ), .ZN(_07286_ ) );
OR3_X1 _15316_ ( .A1(_07074_ ), .A2(_07075_ ), .A3(_06790_ ), .ZN(_07287_ ) );
NAND3_X1 _15317_ ( .A1(_07081_ ), .A2(_07082_ ), .A3(_06791_ ), .ZN(_07288_ ) );
AND3_X1 _15318_ ( .A1(_07287_ ), .A2(_06702_ ), .A3(_07288_ ), .ZN(_07289_ ) );
NAND3_X1 _15319_ ( .A1(_07069_ ), .A2(_06676_ ), .A3(_07070_ ), .ZN(_07290_ ) );
NAND3_X1 _15320_ ( .A1(_07077_ ), .A2(_06818_ ), .A3(_07078_ ), .ZN(_07291_ ) );
AOI21_X1 _15321_ ( .A(_06702_ ), .B1(_07290_ ), .B2(_07291_ ), .ZN(_07292_ ) );
OAI21_X1 _15322_ ( .A(_07248_ ), .B1(_07289_ ), .B2(_07292_ ), .ZN(_07293_ ) );
NAND4_X1 _15323_ ( .A1(_07284_ ), .A2(_07285_ ), .A3(_07286_ ), .A4(_07293_ ), .ZN(_07294_ ) );
OR3_X1 _15324_ ( .A1(_07281_ ), .A2(_07283_ ), .A3(_07294_ ), .ZN(_07295_ ) );
AOI21_X1 _15325_ ( .A(_07264_ ), .B1(_07295_ ), .B2(_06853_ ), .ZN(_07296_ ) );
OAI21_X1 _15326_ ( .A(_06855_ ), .B1(_05506_ ), .B2(_05407_ ), .ZN(_07297_ ) );
OAI21_X1 _15327_ ( .A(_07259_ ), .B1(_07296_ ), .B2(_07297_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_17_D ) );
NOR2_X1 _15328_ ( .A1(_05535_ ), .A2(_05537_ ), .ZN(_07298_ ) );
NAND4_X1 _15329_ ( .A1(_07298_ ), .A2(_05293_ ), .A3(_05719_ ), .A4(_05534_ ), .ZN(_07299_ ) );
NAND3_X1 _15330_ ( .A1(_05840_ ), .A2(_05841_ ), .A3(_06110_ ), .ZN(_07300_ ) );
NAND3_X1 _15331_ ( .A1(_07299_ ), .A2(_07300_ ), .A3(_06434_ ), .ZN(_07301_ ) );
AND2_X1 _15332_ ( .A1(_04106_ ), .A2(_02647_ ), .ZN(_07302_ ) );
AOI21_X1 _15333_ ( .A(_07302_ ), .B1(_07198_ ), .B2(_04107_ ), .ZN(_07303_ ) );
XNOR2_X1 _15334_ ( .A(_07303_ ), .B(_04078_ ), .ZN(_07304_ ) );
NAND2_X1 _15335_ ( .A1(_07304_ ), .A2(_06974_ ), .ZN(_07305_ ) );
AOI22_X1 _15336_ ( .A1(_05525_ ), .A2(_07205_ ), .B1(\ID_EX_imm [13] ), .B2(_07206_ ), .ZN(_07306_ ) );
AOI21_X1 _15337_ ( .A(_07197_ ), .B1(_07305_ ), .B2(_07306_ ), .ZN(_07307_ ) );
OR2_X1 _15338_ ( .A1(_07307_ ), .A2(_05609_ ), .ZN(_07308_ ) );
AND2_X1 _15339_ ( .A1(_06771_ ), .A2(_06770_ ), .ZN(_07309_ ) );
INV_X1 _15340_ ( .A(_07309_ ), .ZN(_07310_ ) );
NAND4_X1 _15341_ ( .A1(_07097_ ), .A2(_06766_ ), .A3(_06762_ ), .A4(_07310_ ), .ZN(_07311_ ) );
NAND3_X1 _15342_ ( .A1(_07122_ ), .A2(_06693_ ), .A3(_07123_ ), .ZN(_07312_ ) );
OAI21_X1 _15343_ ( .A(_06951_ ), .B1(_06780_ ), .B2(_07018_ ), .ZN(_07313_ ) );
OAI211_X1 _15344_ ( .A(_06819_ ), .B(_06820_ ), .C1(_06807_ ), .C2(_06809_ ), .ZN(_07314_ ) );
NAND3_X1 _15345_ ( .A1(_07313_ ), .A2(_06805_ ), .A3(_07314_ ), .ZN(_07315_ ) );
NAND3_X1 _15346_ ( .A1(_07312_ ), .A2(_07315_ ), .A3(_06703_ ), .ZN(_07316_ ) );
OAI211_X1 _15347_ ( .A(_06838_ ), .B(_07316_ ), .C1(_06701_ ), .C2(_06704_ ), .ZN(_07317_ ) );
NAND3_X1 _15348_ ( .A1(_06678_ ), .A2(_06877_ ), .A3(_07063_ ), .ZN(_07318_ ) );
AND2_X1 _15349_ ( .A1(_07317_ ), .A2(_07318_ ), .ZN(_07319_ ) );
AOI21_X1 _15350_ ( .A(_06718_ ), .B1(_07311_ ), .B2(_07319_ ), .ZN(_07320_ ) );
NAND3_X1 _15351_ ( .A1(_07214_ ), .A2(_04832_ ), .A3(_07215_ ), .ZN(_07321_ ) );
OAI21_X1 _15352_ ( .A(_04833_ ), .B1(_07213_ ), .B2(_06610_ ), .ZN(_07322_ ) );
AOI21_X1 _15353_ ( .A(_06590_ ), .B1(_07321_ ), .B2(_07322_ ), .ZN(_07323_ ) );
OAI21_X1 _15354_ ( .A(_06702_ ), .B1(_06789_ ), .B2(_06803_ ), .ZN(_07324_ ) );
OAI21_X1 _15355_ ( .A(_07324_ ), .B1(_06837_ ), .B2(_06703_ ), .ZN(_07325_ ) );
AND2_X1 _15356_ ( .A1(_07325_ ), .A2(_07247_ ), .ZN(_07326_ ) );
AOI221_X4 _15357_ ( .A(_07326_ ), .B1(_06609_ ), .B2(_06586_ ), .C1(_04832_ ), .C2(_07041_ ), .ZN(_07327_ ) );
OR2_X1 _15358_ ( .A1(_07319_ ), .A2(_07065_ ), .ZN(_07328_ ) );
OR2_X1 _15359_ ( .A1(_07210_ ), .A2(_06713_ ), .ZN(_07329_ ) );
NAND3_X1 _15360_ ( .A1(_07327_ ), .A2(_07328_ ), .A3(_07329_ ), .ZN(_07330_ ) );
OR3_X1 _15361_ ( .A1(_07320_ ), .A2(_07323_ ), .A3(_07330_ ), .ZN(_07331_ ) );
AOI21_X1 _15362_ ( .A(_07308_ ), .B1(_07331_ ), .B2(_06853_ ), .ZN(_07332_ ) );
NAND2_X1 _15363_ ( .A1(_05528_ ), .A2(_05610_ ), .ZN(_07333_ ) );
NAND2_X1 _15364_ ( .A1(_07333_ ), .A2(_06422_ ), .ZN(_07334_ ) );
OAI21_X1 _15365_ ( .A(_07301_ ), .B1(_07332_ ), .B2(_07334_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_18_D ) );
NAND3_X1 _15366_ ( .A1(_05557_ ), .A2(_05559_ ), .A3(_06434_ ), .ZN(_07335_ ) );
AOI21_X1 _15367_ ( .A(_06576_ ), .B1(_07198_ ), .B2(_04107_ ), .ZN(_07336_ ) );
OAI21_X1 _15368_ ( .A(_07336_ ), .B1(_04107_ ), .B2(_07198_ ), .ZN(_07337_ ) );
AOI22_X1 _15369_ ( .A1(_05548_ ), .A2(_07205_ ), .B1(\ID_EX_imm [12] ), .B2(_07206_ ), .ZN(_07338_ ) );
AOI21_X1 _15370_ ( .A(_07197_ ), .B1(_07337_ ), .B2(_07338_ ), .ZN(_07339_ ) );
OR2_X1 _15371_ ( .A1(_07339_ ), .A2(_05609_ ), .ZN(_07340_ ) );
NOR3_X1 _15372_ ( .A1(_06720_ ), .A2(_06901_ ), .A3(_07008_ ), .ZN(_07341_ ) );
INV_X1 _15373_ ( .A(_07341_ ), .ZN(_07342_ ) );
NAND4_X1 _15374_ ( .A1(_07097_ ), .A2(_06766_ ), .A3(_06762_ ), .A4(_07342_ ), .ZN(_07343_ ) );
OR3_X1 _15375_ ( .A1(_06884_ ), .A2(_06702_ ), .A3(_06893_ ), .ZN(_07344_ ) );
NAND3_X1 _15376_ ( .A1(_07166_ ), .A2(_06677_ ), .A3(_07167_ ), .ZN(_07345_ ) );
NAND4_X1 _15377_ ( .A1(_06909_ ), .A2(_06914_ ), .A3(_06819_ ), .A4(_06820_ ), .ZN(_07346_ ) );
NAND3_X1 _15378_ ( .A1(_06767_ ), .A2(_06912_ ), .A3(_06931_ ), .ZN(_07347_ ) );
NAND3_X1 _15379_ ( .A1(_07346_ ), .A2(_07347_ ), .A3(_06805_ ), .ZN(_07348_ ) );
NAND2_X1 _15380_ ( .A1(_07345_ ), .A2(_07348_ ), .ZN(_07349_ ) );
OAI211_X1 _15381_ ( .A(_07344_ ), .B(_06838_ ), .C1(_07349_ ), .C2(_06839_ ), .ZN(_07350_ ) );
AND3_X1 _15382_ ( .A1(_06900_ ), .A2(_06702_ ), .A3(_07013_ ), .ZN(_07351_ ) );
OR2_X1 _15383_ ( .A1(_07351_ ), .A2(_06943_ ), .ZN(_07352_ ) );
NAND2_X1 _15384_ ( .A1(_07350_ ), .A2(_07352_ ), .ZN(_07353_ ) );
AOI21_X1 _15385_ ( .A(_06718_ ), .B1(_07343_ ), .B2(_07353_ ), .ZN(_07354_ ) );
AND3_X1 _15386_ ( .A1(_07212_ ), .A2(_04838_ ), .A3(_06601_ ), .ZN(_07355_ ) );
NOR3_X1 _15387_ ( .A1(_07355_ ), .A2(_07213_ ), .A3(_06590_ ), .ZN(_07356_ ) );
NOR2_X1 _15388_ ( .A1(_06933_ ), .A2(_06940_ ), .ZN(_07357_ ) );
NOR2_X1 _15389_ ( .A1(_07357_ ), .A2(_06839_ ), .ZN(_07358_ ) );
AOI21_X1 _15390_ ( .A(_06704_ ), .B1(_06950_ ), .B2(_06953_ ), .ZN(_07359_ ) );
OAI21_X1 _15391_ ( .A(_07248_ ), .B1(_07358_ ), .B2(_07359_ ), .ZN(_07360_ ) );
OAI221_X1 _15392_ ( .A(_07360_ ), .B1(_07215_ ), .B2(_04766_ ), .C1(_04838_ ), .C2(_05026_ ), .ZN(_07361_ ) );
AND3_X1 _15393_ ( .A1(_07350_ ), .A2(_06709_ ), .A3(_07352_ ), .ZN(_07362_ ) );
AOI21_X1 _15394_ ( .A(_04771_ ), .B1(_04836_ ), .B2(_04079_ ), .ZN(_07363_ ) );
OR3_X1 _15395_ ( .A1(_07361_ ), .A2(_07362_ ), .A3(_07363_ ), .ZN(_07364_ ) );
OR3_X1 _15396_ ( .A1(_07354_ ), .A2(_07356_ ), .A3(_07364_ ), .ZN(_07365_ ) );
AOI21_X1 _15397_ ( .A(_07340_ ), .B1(_07365_ ), .B2(_06853_ ), .ZN(_07366_ ) );
OAI21_X1 _15398_ ( .A(_06855_ ), .B1(_05547_ ), .B2(_05407_ ), .ZN(_07367_ ) );
OAI21_X1 _15399_ ( .A(_07335_ ), .B1(_07366_ ), .B2(_07367_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_19_D ) );
AND2_X1 _15400_ ( .A1(_05222_ ), .A2(_07205_ ), .ZN(_07368_ ) );
AOI211_X1 _15401_ ( .A(_04563_ ), .B(_04462_ ), .C1(_05043_ ), .C2(_05058_ ), .ZN(_07369_ ) );
OAI211_X1 _15402_ ( .A(_04711_ ), .B(_04760_ ), .C1(_07369_ ), .C2(_05096_ ), .ZN(_07370_ ) );
AND2_X1 _15403_ ( .A1(_07370_ ), .A2(_05074_ ), .ZN(_07371_ ) );
INV_X1 _15404_ ( .A(_04610_ ), .ZN(_07372_ ) );
NOR4_X1 _15405_ ( .A1(_07371_ ), .A2(_07372_ ), .A3(_04586_ ), .A4(_04587_ ), .ZN(_07373_ ) );
OR2_X1 _15406_ ( .A1(_07373_ ), .A2(_05064_ ), .ZN(_07374_ ) );
AOI21_X1 _15407_ ( .A(_06575_ ), .B1(_07374_ ), .B2(_04658_ ), .ZN(_07375_ ) );
OAI21_X1 _15408_ ( .A(_07375_ ), .B1(_04658_ ), .B2(_07374_ ), .ZN(_07376_ ) );
OAI21_X1 _15409_ ( .A(_07376_ ), .B1(_02964_ ), .B2(_06566_ ), .ZN(_07377_ ) );
OAI21_X1 _15410_ ( .A(_06582_ ), .B1(_07368_ ), .B2(_07377_ ), .ZN(_07378_ ) );
AND2_X1 _15411_ ( .A1(_07278_ ), .A2(_06702_ ), .ZN(_07379_ ) );
AND2_X1 _15412_ ( .A1(_07379_ ), .A2(_06706_ ), .ZN(_07380_ ) );
NOR4_X1 _15413_ ( .A1(_06747_ ), .A2(_06759_ ), .A3(_06874_ ), .A4(_07266_ ), .ZN(_07381_ ) );
AOI211_X1 _15414_ ( .A(_07380_ ), .B(_07381_ ), .C1(_06763_ ), .C2(_06764_ ), .ZN(_07382_ ) );
NOR2_X1 _15415_ ( .A1(_07382_ ), .A2(_06717_ ), .ZN(_07383_ ) );
OR3_X1 _15416_ ( .A1(_07289_ ), .A2(_06943_ ), .A3(_07292_ ), .ZN(_07384_ ) );
OAI21_X1 _15417_ ( .A(_06671_ ), .B1(_06881_ ), .B2(_06879_ ), .ZN(_07385_ ) );
OAI211_X1 _15418_ ( .A(_04861_ ), .B(_06690_ ), .C1(_06890_ ), .C2(_06878_ ), .ZN(_07386_ ) );
NAND2_X1 _15419_ ( .A1(_07385_ ), .A2(_07386_ ), .ZN(_07387_ ) );
OAI21_X1 _15420_ ( .A(_06671_ ), .B1(_06895_ ), .B2(_06897_ ), .ZN(_07388_ ) );
NOR2_X1 _15421_ ( .A1(_06882_ ), .A2(_06898_ ), .ZN(_07389_ ) );
OAI21_X1 _15422_ ( .A(_07388_ ), .B1(_06797_ ), .B2(_07389_ ), .ZN(_07390_ ) );
MUX2_X1 _15423_ ( .A(_07387_ ), .B(_07390_ ), .S(_06791_ ), .Z(_07391_ ) );
OAI21_X1 _15424_ ( .A(_06675_ ), .B1(_07084_ ), .B2(_07086_ ), .ZN(_07392_ ) );
AOI211_X1 _15425_ ( .A(_06891_ ), .B(_06886_ ), .C1(_06689_ ), .C2(_04863_ ), .ZN(_07393_ ) );
NOR3_X1 _15426_ ( .A1(_06671_ ), .A2(_06885_ ), .A3(_06917_ ), .ZN(_07394_ ) );
OAI21_X1 _15427_ ( .A(_06790_ ), .B1(_07393_ ), .B2(_07394_ ), .ZN(_07395_ ) );
AND2_X1 _15428_ ( .A1(_07392_ ), .A2(_07395_ ), .ZN(_07396_ ) );
MUX2_X1 _15429_ ( .A(_07391_ ), .B(_07396_ ), .S(_06813_ ), .Z(_07397_ ) );
AOI21_X1 _15430_ ( .A(_06776_ ), .B1(_07397_ ), .B2(_06838_ ), .ZN(_07398_ ) );
AOI221_X4 _15431_ ( .A(_07383_ ), .B1(_06709_ ), .B2(_07380_ ), .C1(_07384_ ), .C2(_07398_ ), .ZN(_07399_ ) );
NAND2_X1 _15432_ ( .A1(_05013_ ), .A2(_07042_ ), .ZN(_07400_ ) );
NAND3_X1 _15433_ ( .A1(_06341_ ), .A2(_05012_ ), .A3(_07092_ ), .ZN(_07401_ ) );
OAI21_X1 _15434_ ( .A(_06959_ ), .B1(_06341_ ), .B2(_05012_ ), .ZN(_07402_ ) );
NAND4_X1 _15435_ ( .A1(_07399_ ), .A2(_07400_ ), .A3(_07401_ ), .A4(_07402_ ), .ZN(_07403_ ) );
AND2_X1 _15436_ ( .A1(_04951_ ), .A2(_04955_ ), .ZN(_07404_ ) );
NAND4_X1 _15437_ ( .A1(_06656_ ), .A2(_04946_ ), .A3(_04939_ ), .A4(_07404_ ), .ZN(_07405_ ) );
INV_X1 _15438_ ( .A(_04939_ ), .ZN(_07406_ ) );
AOI21_X1 _15439_ ( .A(_04980_ ), .B1(_04951_ ), .B2(_06658_ ), .ZN(_07407_ ) );
INV_X1 _15440_ ( .A(_04946_ ), .ZN(_07408_ ) );
NOR3_X1 _15441_ ( .A1(_07406_ ), .A2(_07407_ ), .A3(_07408_ ), .ZN(_07409_ ) );
NOR4_X1 _15442_ ( .A1(_04944_ ), .A2(_04938_ ), .A3(_04538_ ), .A4(_04945_ ), .ZN(_07410_ ) );
NOR3_X1 _15443_ ( .A1(_07409_ ), .A2(_04944_ ), .A3(_07410_ ), .ZN(_07411_ ) );
AND2_X2 _15444_ ( .A1(_07405_ ), .A2(_07411_ ), .ZN(_07412_ ) );
INV_X2 _15445_ ( .A(_07412_ ), .ZN(_07413_ ) );
NAND3_X4 _15446_ ( .A1(_07413_ ), .A2(_04810_ ), .A3(_04816_ ), .ZN(_07414_ ) );
INV_X1 _15447_ ( .A(_04815_ ), .ZN(_07415_ ) );
AOI21_X1 _15448_ ( .A(_04814_ ), .B1(_04808_ ), .B2(_07415_ ), .ZN(_07416_ ) );
AOI211_X2 _15449_ ( .A(_04802_ ), .B(_04795_ ), .C1(_07414_ ), .C2(_07416_ ), .ZN(_07417_ ) );
AOI21_X1 _15450_ ( .A(_04799_ ), .B1(_04801_ ), .B2(_04792_ ), .ZN(_07418_ ) );
INV_X1 _15451_ ( .A(_07418_ ), .ZN(_07419_ ) );
NOR2_X1 _15452_ ( .A1(_07417_ ), .A2(_07419_ ), .ZN(_07420_ ) );
NOR4_X1 _15453_ ( .A1(_07420_ ), .A2(_04784_ ), .A3(_04785_ ), .A4(_04780_ ), .ZN(_07421_ ) );
INV_X1 _15454_ ( .A(_07421_ ), .ZN(_07422_ ) );
INV_X1 _15455_ ( .A(_04785_ ), .ZN(_07423_ ) );
AND2_X1 _15456_ ( .A1(_04777_ ), .A2(_02167_ ), .ZN(_07424_ ) );
OAI21_X1 _15457_ ( .A(_07423_ ), .B1(_04784_ ), .B2(_07424_ ), .ZN(_07425_ ) );
AND2_X1 _15458_ ( .A1(_07422_ ), .A2(_07425_ ), .ZN(_07426_ ) );
XNOR2_X1 _15459_ ( .A(_07426_ ), .B(_05013_ ), .ZN(_07427_ ) );
AOI21_X1 _15460_ ( .A(_07403_ ), .B1(_07427_ ), .B2(_07221_ ), .ZN(_07428_ ) );
OAI211_X1 _15461_ ( .A(_05347_ ), .B(_07378_ ), .C1(_07428_ ), .C2(_06851_ ), .ZN(_07429_ ) );
NAND2_X1 _15462_ ( .A1(_03912_ ), .A2(_05610_ ), .ZN(_07430_ ) );
NAND3_X1 _15463_ ( .A1(_07429_ ), .A2(_06214_ ), .A3(_07430_ ), .ZN(_07431_ ) );
OR2_X1 _15464_ ( .A1(_05294_ ), .A2(_06221_ ), .ZN(_07432_ ) );
NAND2_X1 _15465_ ( .A1(_07431_ ), .A2(_07432_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_1_D ) );
INV_X1 _15466_ ( .A(_05581_ ), .ZN(_07433_ ) );
INV_X1 _15467_ ( .A(_05578_ ), .ZN(_07434_ ) );
OAI211_X1 _15468_ ( .A(_07433_ ), .B(_06434_ ), .C1(_06516_ ), .C2(_07434_ ), .ZN(_07435_ ) );
NAND3_X1 _15469_ ( .A1(_05042_ ), .A2(_04023_ ), .A3(_04048_ ), .ZN(_07436_ ) );
OAI21_X1 _15470_ ( .A(_07436_ ), .B1(_05051_ ), .B2(_05050_ ), .ZN(_07437_ ) );
AND2_X1 _15471_ ( .A1(_07437_ ), .A2(_03992_ ), .ZN(_07438_ ) );
AOI21_X1 _15472_ ( .A(_07438_ ), .B1(_02742_ ), .B2(_03991_ ), .ZN(_07439_ ) );
XNOR2_X1 _15473_ ( .A(_07439_ ), .B(_03965_ ), .ZN(_07440_ ) );
NAND2_X1 _15474_ ( .A1(_07440_ ), .A2(_06974_ ), .ZN(_07441_ ) );
AOI22_X1 _15475_ ( .A1(_05568_ ), .A2(_07205_ ), .B1(\ID_EX_imm [11] ), .B2(_07206_ ), .ZN(_07442_ ) );
AOI21_X1 _15476_ ( .A(_07197_ ), .B1(_07441_ ), .B2(_07442_ ), .ZN(_07443_ ) );
OR2_X1 _15477_ ( .A1(_07443_ ), .A2(_05609_ ), .ZN(_07444_ ) );
AND2_X1 _15478_ ( .A1(_06762_ ), .A2(_06764_ ), .ZN(_07445_ ) );
OAI211_X1 _15479_ ( .A(_07097_ ), .B(_07445_ ), .C1(_06867_ ), .C2(_06996_ ), .ZN(_07446_ ) );
OAI21_X1 _15480_ ( .A(_06815_ ), .B1(_06786_ ), .B2(_06781_ ), .ZN(_07447_ ) );
OAI211_X1 _15481_ ( .A(_06819_ ), .B(_06820_ ), .C1(_06780_ ), .C2(_07018_ ), .ZN(_07448_ ) );
AOI21_X1 _15482_ ( .A(_06677_ ), .B1(_07447_ ), .B2(_07448_ ), .ZN(_07449_ ) );
AOI21_X1 _15483_ ( .A(_06805_ ), .B1(_07230_ ), .B2(_07231_ ), .ZN(_07450_ ) );
OR3_X1 _15484_ ( .A1(_07449_ ), .A2(_07450_ ), .A3(_06839_ ), .ZN(_07451_ ) );
OAI211_X1 _15485_ ( .A(_07451_ ), .B(_07000_ ), .C1(_07001_ ), .C2(_06993_ ), .ZN(_07452_ ) );
AOI21_X1 _15486_ ( .A(_06839_ ), .B1(_06980_ ), .B2(_06981_ ), .ZN(_07453_ ) );
OR2_X1 _15487_ ( .A1(_07453_ ), .A2(_06707_ ), .ZN(_07454_ ) );
NAND2_X1 _15488_ ( .A1(_07452_ ), .A2(_07454_ ), .ZN(_07455_ ) );
AOI21_X1 _15489_ ( .A(_06718_ ), .B1(_07446_ ), .B2(_07455_ ), .ZN(_07456_ ) );
INV_X1 _15490_ ( .A(_07247_ ), .ZN(_07457_ ) );
NAND3_X1 _15491_ ( .A1(_07030_ ), .A2(_06901_ ), .A3(_06868_ ), .ZN(_07458_ ) );
NAND3_X1 _15492_ ( .A1(_07009_ ), .A2(_07025_ ), .A3(_07015_ ), .ZN(_07459_ ) );
AOI21_X1 _15493_ ( .A(_07457_ ), .B1(_07458_ ), .B2(_07459_ ), .ZN(_07460_ ) );
AOI21_X1 _15494_ ( .A(_04771_ ), .B1(_04852_ ), .B2(_03916_ ), .ZN(_07461_ ) );
NAND3_X1 _15495_ ( .A1(_04924_ ), .A2(_02765_ ), .A3(_06586_ ), .ZN(_07462_ ) );
OAI21_X1 _15496_ ( .A(_07462_ ), .B1(_04922_ ), .B2(_05026_ ), .ZN(_07463_ ) );
OR3_X1 _15497_ ( .A1(_07460_ ), .A2(_07461_ ), .A3(_07463_ ), .ZN(_07464_ ) );
OAI21_X1 _15498_ ( .A(_04857_ ), .B1(_06638_ ), .B2(_06594_ ), .ZN(_07465_ ) );
INV_X1 _15499_ ( .A(_06599_ ), .ZN(_07466_ ) );
NAND2_X1 _15500_ ( .A1(_07465_ ), .A2(_07466_ ), .ZN(_07467_ ) );
AOI21_X1 _15501_ ( .A(_06590_ ), .B1(_07467_ ), .B2(_04853_ ), .ZN(_07468_ ) );
OAI21_X1 _15502_ ( .A(_07468_ ), .B1(_04853_ ), .B2(_07467_ ), .ZN(_07469_ ) );
OAI21_X1 _15503_ ( .A(_07469_ ), .B1(_07065_ ), .B2(_07455_ ), .ZN(_07470_ ) );
OR3_X1 _15504_ ( .A1(_07456_ ), .A2(_07464_ ), .A3(_07470_ ), .ZN(_07471_ ) );
AOI21_X1 _15505_ ( .A(_07444_ ), .B1(_07471_ ), .B2(_06853_ ), .ZN(_07472_ ) );
NAND2_X1 _15506_ ( .A1(_05570_ ), .A2(_03892_ ), .ZN(_07473_ ) );
NAND2_X1 _15507_ ( .A1(_07473_ ), .A2(_06422_ ), .ZN(_07474_ ) );
OAI21_X1 _15508_ ( .A(_07435_ ), .B1(_07472_ ), .B2(_07474_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_20_D ) );
OAI21_X1 _15509_ ( .A(_06288_ ), .B1(_05618_ ), .B2(_05619_ ), .ZN(_07475_ ) );
AOI21_X1 _15510_ ( .A(_06576_ ), .B1(_07437_ ), .B2(_03992_ ), .ZN(_07476_ ) );
OAI21_X1 _15511_ ( .A(_07476_ ), .B1(_03992_ ), .B2(_07437_ ), .ZN(_07477_ ) );
AOI22_X1 _15512_ ( .A1(_05624_ ), .A2(_07205_ ), .B1(\ID_EX_imm [10] ), .B2(_06564_ ), .ZN(_07478_ ) );
AOI21_X1 _15513_ ( .A(_07197_ ), .B1(_07477_ ), .B2(_07478_ ), .ZN(_07479_ ) );
OR2_X1 _15514_ ( .A1(_07479_ ), .A2(_05609_ ), .ZN(_07480_ ) );
AND2_X1 _15515_ ( .A1(_06760_ ), .A2(_06867_ ), .ZN(_07481_ ) );
INV_X1 _15516_ ( .A(_06996_ ), .ZN(_07482_ ) );
NOR4_X1 _15517_ ( .A1(_06747_ ), .A2(_07098_ ), .A3(_06759_ ), .A4(_07482_ ), .ZN(_07483_ ) );
OAI21_X1 _15518_ ( .A(_07445_ ), .B1(_07481_ ), .B2(_07483_ ), .ZN(_07484_ ) );
NAND3_X1 _15519_ ( .A1(_07058_ ), .A2(_07135_ ), .A3(_07061_ ), .ZN(_07485_ ) );
OAI211_X1 _15520_ ( .A(_06815_ ), .B(_06929_ ), .C1(_02742_ ), .C2(_06664_ ), .ZN(_07486_ ) );
NAND4_X1 _15521_ ( .A1(_06912_ ), .A2(_06931_ ), .A3(_06819_ ), .A4(_06820_ ), .ZN(_07487_ ) );
AND3_X1 _15522_ ( .A1(_07486_ ), .A2(_06818_ ), .A3(_07487_ ), .ZN(_07488_ ) );
AOI21_X1 _15523_ ( .A(_07013_ ), .B1(_07272_ ), .B2(_07273_ ), .ZN(_07489_ ) );
NOR2_X1 _15524_ ( .A1(_07488_ ), .A2(_07489_ ), .ZN(_07490_ ) );
OAI211_X1 _15525_ ( .A(_07485_ ), .B(_06943_ ), .C1(_07490_ ), .C2(_06839_ ), .ZN(_07491_ ) );
AOI21_X1 _15526_ ( .A(_07135_ ), .B1(_07050_ ), .B2(_07053_ ), .ZN(_07492_ ) );
NAND2_X1 _15527_ ( .A1(_07492_ ), .A2(_06876_ ), .ZN(_07493_ ) );
AND2_X1 _15528_ ( .A1(_07491_ ), .A2(_07493_ ), .ZN(_07494_ ) );
AOI21_X1 _15529_ ( .A(_06718_ ), .B1(_07484_ ), .B2(_07494_ ), .ZN(_07495_ ) );
AOI21_X1 _15530_ ( .A(_06713_ ), .B1(_04856_ ), .B2(_06598_ ), .ZN(_07496_ ) );
OR3_X1 _15531_ ( .A1(_06638_ ), .A2(_04857_ ), .A3(_06594_ ), .ZN(_07497_ ) );
NAND3_X1 _15532_ ( .A1(_07497_ ), .A2(_06589_ ), .A3(_07465_ ), .ZN(_07498_ ) );
OR2_X1 _15533_ ( .A1(_07494_ ), .A2(_07065_ ), .ZN(_07499_ ) );
OR2_X1 _15534_ ( .A1(_07071_ ), .A2(_07025_ ), .ZN(_07500_ ) );
NAND3_X1 _15535_ ( .A1(_07076_ ), .A2(_07001_ ), .A3(_07079_ ), .ZN(_07501_ ) );
NAND3_X1 _15536_ ( .A1(_07500_ ), .A2(_07501_ ), .A3(_07248_ ), .ZN(_07502_ ) );
AOI22_X1 _15537_ ( .A1(_04857_ ), .A2(_07041_ ), .B1(_06599_ ), .B2(_06586_ ), .ZN(_07503_ ) );
NAND4_X1 _15538_ ( .A1(_07498_ ), .A2(_07499_ ), .A3(_07502_ ), .A4(_07503_ ), .ZN(_07504_ ) );
OR3_X1 _15539_ ( .A1(_07495_ ), .A2(_07496_ ), .A3(_07504_ ), .ZN(_07505_ ) );
BUF_X4 _15540_ ( .A(_06852_ ), .Z(_07506_ ) );
AOI21_X1 _15541_ ( .A(_07480_ ), .B1(_07505_ ), .B2(_07506_ ), .ZN(_07507_ ) );
OAI21_X1 _15542_ ( .A(_06855_ ), .B1(_05622_ ), .B2(_05407_ ), .ZN(_07508_ ) );
OAI21_X1 _15543_ ( .A(_07475_ ), .B1(_07507_ ), .B2(_07508_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_21_D ) );
NAND2_X1 _15544_ ( .A1(_05646_ ), .A2(_06223_ ), .ZN(_07509_ ) );
AOI21_X1 _15545_ ( .A(_05049_ ), .B1(_05042_ ), .B2(_04023_ ), .ZN(_07510_ ) );
XNOR2_X1 _15546_ ( .A(_07510_ ), .B(_04048_ ), .ZN(_07511_ ) );
NAND2_X1 _15547_ ( .A1(_07511_ ), .A2(_06858_ ), .ZN(_07512_ ) );
AOI22_X1 _15548_ ( .A1(_05634_ ), .A2(_07205_ ), .B1(\ID_EX_imm [9] ), .B2(_06564_ ), .ZN(_07513_ ) );
AOI21_X1 _15549_ ( .A(_07197_ ), .B1(_07512_ ), .B2(_07513_ ), .ZN(_07514_ ) );
OR2_X1 _15550_ ( .A1(_07514_ ), .A2(_05609_ ), .ZN(_07515_ ) );
INV_X1 _15551_ ( .A(_06769_ ), .ZN(_07516_ ) );
NOR4_X1 _15552_ ( .A1(_06747_ ), .A2(_07516_ ), .A3(_06759_ ), .A4(_07482_ ), .ZN(_07517_ ) );
OAI21_X1 _15553_ ( .A(_07445_ ), .B1(_07481_ ), .B2(_07517_ ), .ZN(_07518_ ) );
OAI21_X1 _15554_ ( .A(_06814_ ), .B1(_07124_ ), .B2(_07125_ ), .ZN(_07519_ ) );
OAI21_X1 _15555_ ( .A(_06951_ ), .B1(_06800_ ), .B2(_06784_ ), .ZN(_07520_ ) );
OAI211_X1 _15556_ ( .A(_07004_ ), .B(_07005_ ), .C1(_06781_ ), .C2(_06786_ ), .ZN(_07521_ ) );
AOI21_X1 _15557_ ( .A(_06693_ ), .B1(_07520_ ), .B2(_07521_ ), .ZN(_07522_ ) );
AOI21_X1 _15558_ ( .A(_07013_ ), .B1(_07313_ ), .B2(_07314_ ), .ZN(_07523_ ) );
NOR2_X1 _15559_ ( .A1(_07522_ ), .A2(_07523_ ), .ZN(_07524_ ) );
OAI211_X1 _15560_ ( .A(_07519_ ), .B(_06838_ ), .C1(_07524_ ), .C2(_06839_ ), .ZN(_07525_ ) );
NAND4_X1 _15561_ ( .A1(_07119_ ), .A2(_06876_ ), .A3(_06704_ ), .A4(_07120_ ), .ZN(_07526_ ) );
AND2_X1 _15562_ ( .A1(_07525_ ), .A2(_07526_ ), .ZN(_07527_ ) );
AOI21_X1 _15563_ ( .A(_06717_ ), .B1(_07518_ ), .B2(_07527_ ), .ZN(_07528_ ) );
AOI21_X1 _15564_ ( .A(_07065_ ), .B1(_07525_ ), .B2(_07526_ ), .ZN(_07529_ ) );
OR3_X1 _15565_ ( .A1(_07136_ ), .A2(_06814_ ), .A3(_07137_ ), .ZN(_07530_ ) );
NAND4_X1 _15566_ ( .A1(_06835_ ), .A2(_07228_ ), .A3(_07014_ ), .A4(_07017_ ), .ZN(_07531_ ) );
AOI21_X1 _15567_ ( .A(_07457_ ), .B1(_07530_ ), .B2(_07531_ ), .ZN(_07532_ ) );
OR3_X1 _15568_ ( .A1(_07528_ ), .A2(_07529_ ), .A3(_07532_ ), .ZN(_07533_ ) );
AOI21_X1 _15569_ ( .A(_04849_ ), .B1(_06628_ ), .B2(_06637_ ), .ZN(_07534_ ) );
OR3_X1 _15570_ ( .A1(_07534_ ), .A2(_04843_ ), .A3(_06592_ ), .ZN(_07535_ ) );
OAI21_X1 _15571_ ( .A(_04843_ ), .B1(_07534_ ), .B2(_06592_ ), .ZN(_07536_ ) );
AND3_X1 _15572_ ( .A1(_07535_ ), .A2(_07221_ ), .A3(_07536_ ), .ZN(_07537_ ) );
AOI22_X1 _15573_ ( .A1(_06591_ ), .A2(_06959_ ), .B1(_04918_ ), .B2(_06586_ ), .ZN(_07538_ ) );
OAI21_X1 _15574_ ( .A(_07538_ ), .B1(_04844_ ), .B2(_05026_ ), .ZN(_07539_ ) );
OR3_X1 _15575_ ( .A1(_07533_ ), .A2(_07537_ ), .A3(_07539_ ), .ZN(_07540_ ) );
AOI21_X1 _15576_ ( .A(_07515_ ), .B1(_07540_ ), .B2(_07506_ ), .ZN(_07541_ ) );
BUF_X4 _15577_ ( .A(_05324_ ), .Z(_07542_ ) );
OAI21_X1 _15578_ ( .A(_06855_ ), .B1(_05631_ ), .B2(_07542_ ), .ZN(_07543_ ) );
OAI21_X1 _15579_ ( .A(_07509_ ), .B1(_07541_ ), .B2(_07543_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_22_D ) );
AOI21_X1 _15580_ ( .A(_06576_ ), .B1(_05042_ ), .B2(_04023_ ), .ZN(_07544_ ) );
OAI21_X1 _15581_ ( .A(_07544_ ), .B1(_04023_ ), .B2(_05042_ ), .ZN(_07545_ ) );
AOI22_X1 _15582_ ( .A1(_05663_ ), .A2(_07205_ ), .B1(\ID_EX_imm [8] ), .B2(_07206_ ), .ZN(_07546_ ) );
AOI21_X1 _15583_ ( .A(_07197_ ), .B1(_07545_ ), .B2(_07546_ ), .ZN(_07547_ ) );
NOR2_X1 _15584_ ( .A1(_07547_ ), .A2(_03892_ ), .ZN(_07548_ ) );
OAI211_X1 _15585_ ( .A(_06763_ ), .B(_06766_ ), .C1(_07229_ ), .C2(_06721_ ), .ZN(_07549_ ) );
OR3_X1 _15586_ ( .A1(_07172_ ), .A2(_06943_ ), .A3(_07135_ ), .ZN(_07550_ ) );
OAI21_X1 _15587_ ( .A(_06767_ ), .B1(_06934_ ), .B2(_06924_ ), .ZN(_07551_ ) );
OAI211_X1 _15588_ ( .A(_06888_ ), .B(_06889_ ), .C1(_06928_ ), .C2(_06925_ ), .ZN(_07552_ ) );
AND3_X1 _15589_ ( .A1(_07551_ ), .A2(_06791_ ), .A3(_07552_ ), .ZN(_07553_ ) );
AOI21_X1 _15590_ ( .A(_06818_ ), .B1(_07346_ ), .B2(_07347_ ), .ZN(_07554_ ) );
OR3_X1 _15591_ ( .A1(_07553_ ), .A2(_07554_ ), .A3(_07135_ ), .ZN(_07555_ ) );
OAI21_X1 _15592_ ( .A(_06814_ ), .B1(_07168_ ), .B2(_07169_ ), .ZN(_07556_ ) );
NAND3_X1 _15593_ ( .A1(_07555_ ), .A2(_06838_ ), .A3(_07556_ ), .ZN(_07557_ ) );
AND2_X1 _15594_ ( .A1(_07550_ ), .A2(_07557_ ), .ZN(_07558_ ) );
AOI21_X1 _15595_ ( .A(_06718_ ), .B1(_07549_ ), .B2(_07558_ ), .ZN(_07559_ ) );
AOI21_X1 _15596_ ( .A(_07065_ ), .B1(_07550_ ), .B2(_07557_ ), .ZN(_07560_ ) );
NAND3_X1 _15597_ ( .A1(_07182_ ), .A2(_07025_ ), .A3(_07183_ ), .ZN(_07561_ ) );
OR2_X1 _15598_ ( .A1(_07186_ ), .A2(_06704_ ), .ZN(_07562_ ) );
AND3_X1 _15599_ ( .A1(_07561_ ), .A2(_07248_ ), .A3(_07562_ ), .ZN(_07563_ ) );
OR3_X1 _15600_ ( .A1(_07559_ ), .A2(_07560_ ), .A3(_07563_ ), .ZN(_07564_ ) );
AND3_X1 _15601_ ( .A1(_06628_ ), .A2(_06637_ ), .A3(_04849_ ), .ZN(_07565_ ) );
NOR3_X1 _15602_ ( .A1(_07565_ ), .A2(_07534_ ), .A3(_06905_ ), .ZN(_07566_ ) );
AND2_X1 _15603_ ( .A1(_04848_ ), .A2(_07041_ ), .ZN(_07567_ ) );
NOR3_X1 _15604_ ( .A1(_04847_ ), .A2(_04022_ ), .A3(_06843_ ), .ZN(_07568_ ) );
AOI21_X1 _15605_ ( .A(_04771_ ), .B1(_04847_ ), .B2(_04022_ ), .ZN(_07569_ ) );
OR3_X1 _15606_ ( .A1(_07567_ ), .A2(_07568_ ), .A3(_07569_ ), .ZN(_07570_ ) );
NOR3_X1 _15607_ ( .A1(_07564_ ), .A2(_07566_ ), .A3(_07570_ ), .ZN(_07571_ ) );
OAI21_X1 _15608_ ( .A(_07548_ ), .B1(_07571_ ), .B2(_06851_ ), .ZN(_07572_ ) );
NAND2_X1 _15609_ ( .A1(_05661_ ), .A2(_05610_ ), .ZN(_07573_ ) );
NAND3_X1 _15610_ ( .A1(_07572_ ), .A2(_06214_ ), .A3(_07573_ ), .ZN(_07574_ ) );
NAND3_X1 _15611_ ( .A1(_06388_ ), .A2(_06389_ ), .A3(_06223_ ), .ZN(_07575_ ) );
NAND2_X1 _15612_ ( .A1(_07574_ ), .A2(_07575_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_23_D ) );
AND2_X1 _15613_ ( .A1(_05671_ ), .A2(_05670_ ), .ZN(_07576_ ) );
AND2_X1 _15614_ ( .A1(_05672_ ), .A2(_05673_ ), .ZN(_07577_ ) );
AOI21_X1 _15615_ ( .A(_05778_ ), .B1(_07576_ ), .B2(_07577_ ), .ZN(_07578_ ) );
OAI21_X1 _15616_ ( .A(_06288_ ), .B1(_07578_ ), .B2(_05668_ ), .ZN(_07579_ ) );
AND3_X1 _15617_ ( .A1(_05035_ ), .A2(_04235_ ), .A3(_04281_ ), .ZN(_07580_ ) );
OAI21_X1 _15618_ ( .A(_04190_ ), .B1(_07580_ ), .B2(_05039_ ), .ZN(_07581_ ) );
NAND2_X1 _15619_ ( .A1(_04188_ ), .A2(_02565_ ), .ZN(_07582_ ) );
NAND2_X1 _15620_ ( .A1(_07581_ ), .A2(_07582_ ), .ZN(_07583_ ) );
AOI21_X1 _15621_ ( .A(_06576_ ), .B1(_07583_ ), .B2(_04213_ ), .ZN(_07584_ ) );
OAI21_X1 _15622_ ( .A(_07584_ ), .B1(_04213_ ), .B2(_07583_ ), .ZN(_07585_ ) );
AOI22_X1 _15623_ ( .A1(_05679_ ), .A2(_06560_ ), .B1(\ID_EX_imm [7] ), .B2(_06564_ ), .ZN(_07586_ ) );
AOI21_X1 _15624_ ( .A(_07197_ ), .B1(_07585_ ), .B2(_07586_ ), .ZN(_07587_ ) );
OR2_X1 _15625_ ( .A1(_07587_ ), .A2(_05609_ ), .ZN(_07588_ ) );
AND3_X1 _15626_ ( .A1(_06763_ ), .A2(_06766_ ), .A3(_06867_ ), .ZN(_07589_ ) );
AND2_X1 _15627_ ( .A1(_07233_ ), .A2(_06814_ ), .ZN(_07590_ ) );
AND3_X1 _15628_ ( .A1(_07447_ ), .A2(_06682_ ), .A3(_07448_ ), .ZN(_07591_ ) );
NAND4_X1 _15629_ ( .A1(_06785_ ), .A2(_06801_ ), .A3(_06819_ ), .A4(_06820_ ), .ZN(_07592_ ) );
NAND3_X1 _15630_ ( .A1(_06815_ ), .A2(_06799_ ), .A3(_06795_ ), .ZN(_07593_ ) );
AND2_X1 _15631_ ( .A1(_07592_ ), .A2(_07593_ ), .ZN(_07594_ ) );
INV_X1 _15632_ ( .A(_07594_ ), .ZN(_07595_ ) );
AOI211_X1 _15633_ ( .A(_07135_ ), .B(_07591_ ), .C1(_07595_ ), .C2(_07014_ ), .ZN(_07596_ ) );
OR3_X1 _15634_ ( .A1(_07590_ ), .A2(_07596_ ), .A3(_06877_ ), .ZN(_07597_ ) );
OR3_X1 _15635_ ( .A1(_07225_ ), .A2(_06813_ ), .A3(_07226_ ), .ZN(_07598_ ) );
OAI21_X1 _15636_ ( .A(_07598_ ), .B1(_07063_ ), .B2(_07235_ ), .ZN(_07599_ ) );
NAND2_X1 _15637_ ( .A1(_07599_ ), .A2(_06877_ ), .ZN(_07600_ ) );
NAND2_X1 _15638_ ( .A1(_07597_ ), .A2(_07600_ ), .ZN(_07601_ ) );
OAI21_X1 _15639_ ( .A(_06716_ ), .B1(_07589_ ), .B2(_07601_ ), .ZN(_07602_ ) );
NAND2_X1 _15640_ ( .A1(_07601_ ), .A2(_06711_ ), .ZN(_07603_ ) );
OR3_X1 _15641_ ( .A1(_07242_ ), .A2(_07229_ ), .A3(_07457_ ), .ZN(_07604_ ) );
NAND3_X1 _15642_ ( .A1(_07602_ ), .A2(_07603_ ), .A3(_07604_ ), .ZN(_07605_ ) );
XNOR2_X1 _15643_ ( .A(_04894_ ), .B(_02565_ ), .ZN(_07606_ ) );
AND3_X1 _15644_ ( .A1(_06624_ ), .A2(_06625_ ), .A3(_06627_ ), .ZN(_07607_ ) );
OAI21_X1 _15645_ ( .A(_07606_ ), .B1(_07607_ ), .B2(_06636_ ), .ZN(_07608_ ) );
NAND2_X1 _15646_ ( .A1(_07608_ ), .A2(_04895_ ), .ZN(_07609_ ) );
OAI21_X1 _15647_ ( .A(_06589_ ), .B1(_07609_ ), .B2(_04891_ ), .ZN(_07610_ ) );
AOI21_X1 _15648_ ( .A(_07610_ ), .B1(_04891_ ), .B2(_07609_ ), .ZN(_07611_ ) );
NAND2_X1 _15649_ ( .A1(_04891_ ), .A2(_07042_ ), .ZN(_07612_ ) );
NAND2_X1 _15650_ ( .A1(_06630_ ), .A2(_07092_ ), .ZN(_07613_ ) );
OR2_X1 _15651_ ( .A1(_06631_ ), .A2(_06713_ ), .ZN(_07614_ ) );
NAND3_X1 _15652_ ( .A1(_07612_ ), .A2(_07613_ ), .A3(_07614_ ), .ZN(_07615_ ) );
OR3_X1 _15653_ ( .A1(_07605_ ), .A2(_07611_ ), .A3(_07615_ ), .ZN(_07616_ ) );
AOI21_X1 _15654_ ( .A(_07588_ ), .B1(_07616_ ), .B2(_07506_ ), .ZN(_07617_ ) );
OAI21_X1 _15655_ ( .A(_06855_ ), .B1(_05677_ ), .B2(_07542_ ), .ZN(_07618_ ) );
OAI21_X1 _15656_ ( .A(_07579_ ), .B1(_07617_ ), .B2(_07618_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_24_D ) );
AND2_X1 _15657_ ( .A1(_05692_ ), .A2(_03876_ ), .ZN(_07619_ ) );
OR2_X1 _15658_ ( .A1(_06747_ ), .A2(_06759_ ), .ZN(_07620_ ) );
INV_X1 _15659_ ( .A(_07445_ ), .ZN(_07621_ ) );
NOR4_X1 _15660_ ( .A1(_07620_ ), .A2(_06771_ ), .A3(_07621_ ), .A4(_07265_ ), .ZN(_07622_ ) );
MUX2_X1 _15661_ ( .A(_07278_ ), .B(_07270_ ), .S(_06702_ ), .Z(_07623_ ) );
NAND2_X1 _15662_ ( .A1(_07623_ ), .A2(_06877_ ), .ZN(_07624_ ) );
AND3_X1 _15663_ ( .A1(_07486_ ), .A2(_06682_ ), .A3(_07487_ ), .ZN(_07625_ ) );
OAI21_X1 _15664_ ( .A(_06951_ ), .B1(_06938_ ), .B2(_06935_ ), .ZN(_07626_ ) );
OAI211_X1 _15665_ ( .A(_07004_ ), .B(_07005_ ), .C1(_06924_ ), .C2(_06934_ ), .ZN(_07627_ ) );
AOI21_X1 _15666_ ( .A(_06693_ ), .B1(_07626_ ), .B2(_07627_ ), .ZN(_07628_ ) );
OAI21_X1 _15667_ ( .A(_06703_ ), .B1(_07625_ ), .B2(_07628_ ), .ZN(_07629_ ) );
OAI211_X1 _15668_ ( .A(_07629_ ), .B(_06838_ ), .C1(_06704_ ), .C2(_07275_ ), .ZN(_07630_ ) );
NAND2_X1 _15669_ ( .A1(_07624_ ), .A2(_07630_ ), .ZN(_07631_ ) );
OAI21_X1 _15670_ ( .A(_06716_ ), .B1(_07622_ ), .B2(_07631_ ), .ZN(_07632_ ) );
NAND2_X1 _15671_ ( .A1(_07631_ ), .A2(_06710_ ), .ZN(_07633_ ) );
AND2_X1 _15672_ ( .A1(_07290_ ), .A2(_07291_ ), .ZN(_07634_ ) );
OR3_X1 _15673_ ( .A1(_07634_ ), .A2(_06901_ ), .A3(_07457_ ), .ZN(_07635_ ) );
NAND3_X1 _15674_ ( .A1(_07632_ ), .A2(_07633_ ), .A3(_07635_ ), .ZN(_07636_ ) );
NAND3_X1 _15675_ ( .A1(_04895_ ), .A2(_04896_ ), .A3(_07041_ ), .ZN(_07637_ ) );
OR3_X1 _15676_ ( .A1(_04894_ ), .A2(_04189_ ), .A3(_04766_ ), .ZN(_07638_ ) );
NAND2_X1 _15677_ ( .A1(_04896_ ), .A2(_04770_ ), .ZN(_07639_ ) );
NAND3_X1 _15678_ ( .A1(_07637_ ), .A2(_07638_ ), .A3(_07639_ ), .ZN(_07640_ ) );
OR2_X1 _15679_ ( .A1(_07636_ ), .A2(_07640_ ), .ZN(_07641_ ) );
OR3_X1 _15680_ ( .A1(_07607_ ), .A2(_07606_ ), .A3(_06636_ ), .ZN(_07642_ ) );
AND3_X1 _15681_ ( .A1(_07642_ ), .A2(_07221_ ), .A3(_07608_ ), .ZN(_07643_ ) );
OAI21_X1 _15682_ ( .A(_06852_ ), .B1(_07641_ ), .B2(_07643_ ), .ZN(_07644_ ) );
OR3_X1 _15683_ ( .A1(_07580_ ), .A2(_04190_ ), .A3(_05039_ ), .ZN(_07645_ ) );
NAND3_X1 _15684_ ( .A1(_07645_ ), .A2(_06858_ ), .A3(_07581_ ), .ZN(_07646_ ) );
AOI22_X1 _15685_ ( .A1(_05690_ ), .A2(_06560_ ), .B1(\ID_EX_imm [6] ), .B2(_06564_ ), .ZN(_07647_ ) );
AOI21_X1 _15686_ ( .A(_06583_ ), .B1(_07646_ ), .B2(_07647_ ), .ZN(_07648_ ) );
NOR2_X1 _15687_ ( .A1(_07648_ ), .A2(_03876_ ), .ZN(_07649_ ) );
AOI21_X1 _15688_ ( .A(_07619_ ), .B1(_07644_ ), .B2(_07649_ ), .ZN(_07650_ ) );
MUX2_X1 _15689_ ( .A(_05705_ ), .B(_07650_ ), .S(_06221_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_25_D ) );
NAND3_X1 _15690_ ( .A1(_05723_ ), .A2(_05725_ ), .A3(_06434_ ), .ZN(_07651_ ) );
NAND3_X1 _15691_ ( .A1(_06562_ ), .A2(\ID_EX_imm [5] ), .A3(_06559_ ), .ZN(_07652_ ) );
OAI21_X1 _15692_ ( .A(_07652_ ), .B1(_05714_ ), .B2(_06561_ ), .ZN(_07653_ ) );
AND2_X1 _15693_ ( .A1(_04280_ ), .A2(_02611_ ), .ZN(_07654_ ) );
AOI21_X1 _15694_ ( .A(_07654_ ), .B1(_05035_ ), .B2(_04281_ ), .ZN(_07655_ ) );
XNOR2_X1 _15695_ ( .A(_07655_ ), .B(_04235_ ), .ZN(_07656_ ) );
AOI21_X1 _15696_ ( .A(_07653_ ), .B1(_07656_ ), .B2(_06974_ ), .ZN(_07657_ ) );
OAI21_X1 _15697_ ( .A(_05928_ ), .B1(_07657_ ), .B2(_06584_ ), .ZN(_07658_ ) );
NOR4_X1 _15698_ ( .A1(_06873_ ), .A2(_06872_ ), .A3(_06770_ ), .A4(_06771_ ), .ZN(_07659_ ) );
NAND2_X1 _15699_ ( .A1(_06705_ ), .A2(_07032_ ), .ZN(_07660_ ) );
NAND3_X1 _15700_ ( .A1(_07312_ ), .A2(_07315_ ), .A3(_06901_ ), .ZN(_07661_ ) );
NAND3_X1 _15701_ ( .A1(_07520_ ), .A2(_07008_ ), .A3(_07521_ ), .ZN(_07662_ ) );
NOR2_X1 _15702_ ( .A1(_07002_ ), .A2(_06827_ ), .ZN(_07663_ ) );
NAND2_X1 _15703_ ( .A1(_07663_ ), .A2(_07017_ ), .ZN(_07664_ ) );
NAND4_X1 _15704_ ( .A1(_06799_ ), .A2(_06795_ ), .A3(_07004_ ), .A4(_07005_ ), .ZN(_07665_ ) );
AND2_X1 _15705_ ( .A1(_07664_ ), .A2(_07665_ ), .ZN(_07666_ ) );
OAI211_X1 _15706_ ( .A(_07025_ ), .B(_07662_ ), .C1(_07666_ ), .C2(_07008_ ), .ZN(_07667_ ) );
NAND3_X1 _15707_ ( .A1(_07661_ ), .A2(_07000_ ), .A3(_07667_ ), .ZN(_07668_ ) );
NAND2_X1 _15708_ ( .A1(_07660_ ), .A2(_07668_ ), .ZN(_07669_ ) );
OAI21_X1 _15709_ ( .A(_06865_ ), .B1(_07659_ ), .B2(_07669_ ), .ZN(_07670_ ) );
NAND2_X1 _15710_ ( .A1(_06624_ ), .A2(_06625_ ), .ZN(_07671_ ) );
NOR2_X1 _15711_ ( .A1(_07671_ ), .A2(_04908_ ), .ZN(_07672_ ) );
NOR2_X1 _15712_ ( .A1(_07672_ ), .A2(_06634_ ), .ZN(_07673_ ) );
AOI21_X1 _15713_ ( .A(_06905_ ), .B1(_07673_ ), .B2(_04903_ ), .ZN(_07674_ ) );
OAI21_X1 _15714_ ( .A(_07674_ ), .B1(_04903_ ), .B2(_07673_ ), .ZN(_07675_ ) );
NAND2_X1 _15715_ ( .A1(_07669_ ), .A2(_06711_ ), .ZN(_07676_ ) );
OAI21_X1 _15716_ ( .A(_06959_ ), .B1(_04900_ ), .B2(_02589_ ), .ZN(_07677_ ) );
NOR3_X1 _15717_ ( .A1(_06837_ ), .A2(_07228_ ), .A3(_07457_ ), .ZN(_07678_ ) );
AOI221_X4 _15718_ ( .A(_07678_ ), .B1(_06633_ ), .B2(_06586_ ), .C1(_04902_ ), .C2(_07041_ ), .ZN(_07679_ ) );
AND3_X1 _15719_ ( .A1(_07676_ ), .A2(_07677_ ), .A3(_07679_ ), .ZN(_07680_ ) );
NAND3_X1 _15720_ ( .A1(_07670_ ), .A2(_07675_ ), .A3(_07680_ ), .ZN(_07681_ ) );
AOI21_X1 _15721_ ( .A(_07658_ ), .B1(_07681_ ), .B2(_07506_ ), .ZN(_07682_ ) );
OAI21_X1 _15722_ ( .A(_06855_ ), .B1(_05710_ ), .B2(_07542_ ), .ZN(_07683_ ) );
OAI21_X1 _15723_ ( .A(_07651_ ), .B1(_07682_ ), .B2(_07683_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_26_D ) );
AND2_X1 _15724_ ( .A1(_05742_ ), .A2(_03876_ ), .ZN(_07684_ ) );
NAND4_X1 _15725_ ( .A1(_07097_ ), .A2(_06867_ ), .A3(_06869_ ), .A4(_07445_ ), .ZN(_07685_ ) );
AND3_X1 _15726_ ( .A1(_07551_ ), .A2(_06693_ ), .A3(_07552_ ), .ZN(_07686_ ) );
NOR2_X1 _15727_ ( .A1(_06937_ ), .A2(_06944_ ), .ZN(_07687_ ) );
AND2_X1 _15728_ ( .A1(_07687_ ), .A2(_06951_ ), .ZN(_07688_ ) );
NOR3_X1 _15729_ ( .A1(_07011_ ), .A2(_06938_ ), .A3(_06935_ ), .ZN(_07689_ ) );
NOR2_X1 _15730_ ( .A1(_07688_ ), .A2(_07689_ ), .ZN(_07690_ ) );
INV_X1 _15731_ ( .A(_07690_ ), .ZN(_07691_ ) );
AOI211_X1 _15732_ ( .A(_06814_ ), .B(_07686_ ), .C1(_07691_ ), .C2(_07014_ ), .ZN(_07692_ ) );
AOI211_X1 _15733_ ( .A(_06877_ ), .B(_07692_ ), .C1(_07229_ ), .C2(_07349_ ), .ZN(_07693_ ) );
AOI21_X1 _15734_ ( .A(_07174_ ), .B1(_06894_ ), .B2(_06902_ ), .ZN(_07694_ ) );
NOR2_X1 _15735_ ( .A1(_07693_ ), .A2(_07694_ ), .ZN(_07695_ ) );
AOI21_X1 _15736_ ( .A(_06718_ ), .B1(_07685_ ), .B2(_07695_ ), .ZN(_07696_ ) );
OAI21_X1 _15737_ ( .A(_06711_ ), .B1(_07693_ ), .B2(_07694_ ), .ZN(_07697_ ) );
AOI211_X1 _15738_ ( .A(_06876_ ), .B(_06813_ ), .C1(_06950_ ), .C2(_06953_ ), .ZN(_07698_ ) );
AND2_X1 _15739_ ( .A1(_07698_ ), .A2(_05099_ ), .ZN(_07699_ ) );
AOI221_X4 _15740_ ( .A(_07699_ ), .B1(_06634_ ), .B2(_06586_ ), .C1(_04907_ ), .C2(_07041_ ), .ZN(_07700_ ) );
AOI21_X1 _15741_ ( .A(_06590_ ), .B1(_07671_ ), .B2(_04908_ ), .ZN(_07701_ ) );
OAI21_X1 _15742_ ( .A(_07701_ ), .B1(_04908_ ), .B2(_07671_ ), .ZN(_07702_ ) );
OAI21_X1 _15743_ ( .A(_06959_ ), .B1(_07032_ ), .B2(_02611_ ), .ZN(_07703_ ) );
NAND4_X1 _15744_ ( .A1(_07697_ ), .A2(_07700_ ), .A3(_07702_ ), .A4(_07703_ ), .ZN(_07704_ ) );
OAI21_X1 _15745_ ( .A(_06852_ ), .B1(_07696_ ), .B2(_07704_ ), .ZN(_07705_ ) );
AOI21_X1 _15746_ ( .A(_06575_ ), .B1(_05035_ ), .B2(_04281_ ), .ZN(_07706_ ) );
OAI21_X1 _15747_ ( .A(_07706_ ), .B1(_04281_ ), .B2(_05035_ ), .ZN(_07707_ ) );
AOI22_X1 _15748_ ( .A1(_05745_ ), .A2(_06560_ ), .B1(\ID_EX_imm [4] ), .B2(_06564_ ), .ZN(_07708_ ) );
AOI21_X1 _15749_ ( .A(_06583_ ), .B1(_07707_ ), .B2(_07708_ ), .ZN(_07709_ ) );
NOR2_X1 _15750_ ( .A1(_07709_ ), .A2(_03876_ ), .ZN(_07710_ ) );
AOI21_X1 _15751_ ( .A(_07684_ ), .B1(_07705_ ), .B2(_07710_ ), .ZN(_07711_ ) );
MUX2_X1 _15752_ ( .A(_05741_ ), .B(_07711_ ), .S(_06221_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_27_D ) );
NAND2_X1 _15753_ ( .A1(_05762_ ), .A2(_06223_ ), .ZN(_07712_ ) );
AOI21_X1 _15754_ ( .A(_04329_ ), .B1(_05031_ ), .B2(_05032_ ), .ZN(_07713_ ) );
AOI211_X1 _15755_ ( .A(_04330_ ), .B(_04304_ ), .C1(_05030_ ), .C2(_04306_ ), .ZN(_07714_ ) );
OAI21_X1 _15756_ ( .A(_06858_ ), .B1(_07713_ ), .B2(_07714_ ), .ZN(_07715_ ) );
AOI22_X1 _15757_ ( .A1(_05752_ ), .A2(_06560_ ), .B1(\ID_EX_imm [3] ), .B2(_06564_ ), .ZN(_07716_ ) );
AOI21_X1 _15758_ ( .A(_07197_ ), .B1(_07715_ ), .B2(_07716_ ), .ZN(_07717_ ) );
OR2_X1 _15759_ ( .A1(_07717_ ), .A2(_05609_ ), .ZN(_07718_ ) );
AND2_X1 _15760_ ( .A1(_07589_ ), .A2(_06996_ ), .ZN(_07719_ ) );
OAI21_X1 _15761_ ( .A(_07228_ ), .B1(_07449_ ), .B2(_07450_ ), .ZN(_07720_ ) );
NOR2_X1 _15762_ ( .A1(_06828_ ), .A2(_06831_ ), .ZN(_07721_ ) );
MUX2_X1 _15763_ ( .A(_07663_ ), .B(_07721_ ), .S(_07011_ ), .Z(_07722_ ) );
MUX2_X1 _15764_ ( .A(_07722_ ), .B(_07595_ ), .S(_06677_ ), .Z(_07723_ ) );
OAI211_X1 _15765_ ( .A(_07174_ ), .B(_07720_ ), .C1(_07723_ ), .C2(_06901_ ), .ZN(_07724_ ) );
NAND2_X1 _15766_ ( .A1(_06994_ ), .A2(_06877_ ), .ZN(_07725_ ) );
NAND2_X1 _15767_ ( .A1(_07724_ ), .A2(_07725_ ), .ZN(_07726_ ) );
OAI21_X1 _15768_ ( .A(_06865_ ), .B1(_07719_ ), .B2(_07726_ ), .ZN(_07727_ ) );
NOR2_X1 _15769_ ( .A1(_06622_ ), .A2(_06623_ ), .ZN(_07728_ ) );
OAI21_X1 _15770_ ( .A(_04877_ ), .B1(_07728_ ), .B2(_06617_ ), .ZN(_07729_ ) );
OAI221_X1 _15771_ ( .A(_06618_ ), .B1(_04884_ ), .B2(_04885_ ), .C1(_06622_ ), .C2(_06623_ ), .ZN(_07730_ ) );
NAND3_X1 _15772_ ( .A1(_07729_ ), .A2(_07730_ ), .A3(_07221_ ), .ZN(_07731_ ) );
NAND2_X1 _15773_ ( .A1(_04877_ ), .A2(_07041_ ), .ZN(_07732_ ) );
OAI221_X1 _15774_ ( .A(_07732_ ), .B1(_06616_ ), .B2(_04766_ ), .C1(_07031_ ), .C2(_07457_ ), .ZN(_07733_ ) );
AOI221_X4 _15775_ ( .A(_07733_ ), .B1(_06625_ ), .B2(_04770_ ), .C1(_07726_ ), .C2(_06711_ ), .ZN(_07734_ ) );
NAND3_X1 _15776_ ( .A1(_07727_ ), .A2(_07731_ ), .A3(_07734_ ), .ZN(_07735_ ) );
AOI21_X1 _15777_ ( .A(_07718_ ), .B1(_07735_ ), .B2(_07506_ ), .ZN(_07736_ ) );
OAI21_X1 _15778_ ( .A(_06855_ ), .B1(_05325_ ), .B2(_05750_ ), .ZN(_07737_ ) );
OAI21_X1 _15779_ ( .A(_07712_ ), .B1(_07736_ ), .B2(_07737_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_28_D ) );
NOR2_X1 _15780_ ( .A1(_05774_ ), .A2(_05775_ ), .ZN(_07738_ ) );
AOI21_X1 _15781_ ( .A(_05778_ ), .B1(_07738_ ), .B2(_06448_ ), .ZN(_07739_ ) );
OAI21_X1 _15782_ ( .A(_06556_ ), .B1(_07739_ ), .B2(_05770_ ), .ZN(_07740_ ) );
AOI21_X1 _15783_ ( .A(_06576_ ), .B1(_05030_ ), .B2(_04306_ ), .ZN(_07741_ ) );
OAI21_X1 _15784_ ( .A(_07741_ ), .B1(_04306_ ), .B2(_05030_ ), .ZN(_07742_ ) );
AOI22_X1 _15785_ ( .A1(_05767_ ), .A2(_06560_ ), .B1(\ID_EX_imm [2] ), .B2(_06564_ ), .ZN(_07743_ ) );
AOI21_X1 _15786_ ( .A(_06583_ ), .B1(_07742_ ), .B2(_07743_ ), .ZN(_07744_ ) );
OR2_X1 _15787_ ( .A1(_07744_ ), .A2(_05609_ ), .ZN(_07745_ ) );
NAND4_X1 _15788_ ( .A1(_06977_ ), .A2(_07099_ ), .A3(_06867_ ), .A4(_06996_ ), .ZN(_07746_ ) );
NAND2_X1 _15789_ ( .A1(_07064_ ), .A2(_07032_ ), .ZN(_07747_ ) );
AND3_X1 _15790_ ( .A1(_07626_ ), .A2(_06677_ ), .A3(_07627_ ), .ZN(_07748_ ) );
NOR2_X1 _15791_ ( .A1(_06945_ ), .A2(_06947_ ), .ZN(_07749_ ) );
MUX2_X1 _15792_ ( .A(_07687_ ), .B(_07749_ ), .S(_07017_ ), .Z(_07750_ ) );
AOI211_X1 _15793_ ( .A(_07228_ ), .B(_07748_ ), .C1(_06868_ ), .C2(_07750_ ), .ZN(_07751_ ) );
NOR2_X1 _15794_ ( .A1(_07490_ ), .A2(_07025_ ), .ZN(_07752_ ) );
OAI21_X1 _15795_ ( .A(_07000_ ), .B1(_07751_ ), .B2(_07752_ ), .ZN(_07753_ ) );
NAND2_X1 _15796_ ( .A1(_07747_ ), .A2(_07753_ ), .ZN(_07754_ ) );
AOI21_X1 _15797_ ( .A(_06718_ ), .B1(_07746_ ), .B2(_07754_ ), .ZN(_07755_ ) );
AND3_X1 _15798_ ( .A1(_07747_ ), .A2(_06711_ ), .A3(_07753_ ), .ZN(_07756_ ) );
AND4_X1 _15799_ ( .A1(_06708_ ), .A2(_07071_ ), .A3(_07001_ ), .A4(_05099_ ), .ZN(_07757_ ) );
NOR3_X1 _15800_ ( .A1(_07755_ ), .A2(_07756_ ), .A3(_07757_ ), .ZN(_07758_ ) );
AOI21_X1 _15801_ ( .A(_06905_ ), .B1(_06622_ ), .B2(_06623_ ), .ZN(_07759_ ) );
OAI21_X1 _15802_ ( .A(_07759_ ), .B1(_06623_ ), .B2(_06622_ ), .ZN(_07760_ ) );
AOI21_X1 _15803_ ( .A(_04771_ ), .B1(_06868_ ), .B2(_02493_ ), .ZN(_07761_ ) );
AOI221_X4 _15804_ ( .A(_07761_ ), .B1(_06617_ ), .B2(_07092_ ), .C1(_04881_ ), .C2(_07042_ ), .ZN(_07762_ ) );
NAND3_X1 _15805_ ( .A1(_07758_ ), .A2(_07760_ ), .A3(_07762_ ), .ZN(_07763_ ) );
AOI21_X1 _15806_ ( .A(_07745_ ), .B1(_07763_ ), .B2(_07506_ ), .ZN(_07764_ ) );
BUF_X4 _15807_ ( .A(_06317_ ), .Z(_07765_ ) );
OAI21_X1 _15808_ ( .A(_07765_ ), .B1(_05325_ ), .B2(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07766_ ) );
OAI21_X1 _15809_ ( .A(_07740_ ), .B1(_07764_ ), .B2(_07766_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_29_D ) );
OR3_X1 _15810_ ( .A1(_05342_ ), .A2(_05343_ ), .A3(_06317_ ), .ZN(_07767_ ) );
NOR2_X1 _15811_ ( .A1(_07420_ ), .A2(_04780_ ), .ZN(_07768_ ) );
XNOR2_X1 _15812_ ( .A(_04783_ ), .B(_02940_ ), .ZN(_07769_ ) );
OR3_X1 _15813_ ( .A1(_07768_ ), .A2(_07769_ ), .A3(_07424_ ), .ZN(_07770_ ) );
OAI21_X1 _15814_ ( .A(_07769_ ), .B1(_07768_ ), .B2(_07424_ ), .ZN(_07771_ ) );
NAND3_X1 _15815_ ( .A1(_07770_ ), .A2(_07221_ ), .A3(_07771_ ), .ZN(_07772_ ) );
OAI21_X1 _15816_ ( .A(_07228_ ), .B1(_06812_ ), .B2(_06824_ ), .ZN(_07773_ ) );
NAND4_X1 _15817_ ( .A1(_06680_ ), .A2(_06688_ ), .A3(_07004_ ), .A4(_07005_ ), .ZN(_07774_ ) );
NAND3_X1 _15818_ ( .A1(_07017_ ), .A2(_06684_ ), .A3(_06667_ ), .ZN(_07775_ ) );
NAND3_X1 _15819_ ( .A1(_07774_ ), .A2(_07775_ ), .A3(_07014_ ), .ZN(_07776_ ) );
NOR2_X1 _15820_ ( .A1(_06695_ ), .A2(_06698_ ), .ZN(_07777_ ) );
NOR2_X1 _15821_ ( .A1(_06697_ ), .A2(_06989_ ), .ZN(_07778_ ) );
MUX2_X1 _15822_ ( .A(_07777_ ), .B(_07778_ ), .S(_06815_ ), .Z(_07779_ ) );
OAI211_X1 _15823_ ( .A(_07063_ ), .B(_07776_ ), .C1(_07779_ ), .C2(_06868_ ), .ZN(_07780_ ) );
NAND3_X1 _15824_ ( .A1(_07773_ ), .A2(_06707_ ), .A3(_07780_ ), .ZN(_07781_ ) );
AND2_X1 _15825_ ( .A1(_07781_ ), .A2(_05099_ ), .ZN(_07782_ ) );
OAI21_X1 _15826_ ( .A(_07782_ ), .B1(_06708_ ), .B2(_07325_ ), .ZN(_07783_ ) );
OAI211_X1 _15827_ ( .A(_06760_ ), .B(_06762_ ), .C1(_06766_ ), .C2(_07310_ ), .ZN(_07784_ ) );
NOR3_X1 _15828_ ( .A1(_06674_ ), .A2(_07228_ ), .A3(_07008_ ), .ZN(_07785_ ) );
NAND2_X1 _15829_ ( .A1(_07785_ ), .A2(_07174_ ), .ZN(_07786_ ) );
AOI21_X1 _15830_ ( .A(_06717_ ), .B1(_07784_ ), .B2(_07786_ ), .ZN(_07787_ ) );
AND3_X1 _15831_ ( .A1(_07785_ ), .A2(_07174_ ), .A3(_06710_ ), .ZN(_07788_ ) );
NOR2_X1 _15832_ ( .A1(_07787_ ), .A2(_07788_ ), .ZN(_07789_ ) );
NAND3_X1 _15833_ ( .A1(_04783_ ), .A2(_02934_ ), .A3(_07092_ ), .ZN(_07790_ ) );
AOI22_X1 _15834_ ( .A1(_07769_ ), .A2(_07042_ ), .B1(_07423_ ), .B2(_06959_ ), .ZN(_07791_ ) );
AND4_X1 _15835_ ( .A1(_07783_ ), .A2(_07789_ ), .A3(_07790_ ), .A4(_07791_ ), .ZN(_07792_ ) );
AOI21_X1 _15836_ ( .A(_06851_ ), .B1(_07772_ ), .B2(_07792_ ), .ZN(_07793_ ) );
NOR2_X1 _15837_ ( .A1(_05322_ ), .A2(_06861_ ), .ZN(_07794_ ) );
AOI21_X1 _15838_ ( .A(_07794_ ), .B1(\ID_EX_imm [29] ), .B2(_07206_ ), .ZN(_07795_ ) );
NOR2_X1 _15839_ ( .A1(_07371_ ), .A2(_07372_ ), .ZN(_07796_ ) );
OR3_X1 _15840_ ( .A1(_07796_ ), .A2(_05062_ ), .A3(_04588_ ), .ZN(_07797_ ) );
OAI21_X1 _15841_ ( .A(_04588_ ), .B1(_07796_ ), .B2(_05062_ ), .ZN(_07798_ ) );
NAND3_X1 _15842_ ( .A1(_07797_ ), .A2(_06974_ ), .A3(_07798_ ), .ZN(_07799_ ) );
AOI21_X1 _15843_ ( .A(_06584_ ), .B1(_07795_ ), .B2(_07799_ ), .ZN(_07800_ ) );
NOR3_X1 _15844_ ( .A1(_07793_ ), .A2(_05610_ ), .A3(_07800_ ), .ZN(_07801_ ) );
OAI21_X1 _15845_ ( .A(_07765_ ), .B1(_05316_ ), .B2(_07542_ ), .ZN(_07802_ ) );
OAI21_X1 _15846_ ( .A(_07767_ ), .B1(_07801_ ), .B2(_07802_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_2_D ) );
AND2_X1 _15847_ ( .A1(_05787_ ), .A2(_05786_ ), .ZN(_07803_ ) );
AND2_X1 _15848_ ( .A1(_05788_ ), .A2(_05789_ ), .ZN(_07804_ ) );
AOI21_X1 _15849_ ( .A(_05778_ ), .B1(_07803_ ), .B2(_07804_ ), .ZN(_07805_ ) );
OAI21_X1 _15850_ ( .A(_06556_ ), .B1(_07805_ ), .B2(_05784_ ), .ZN(_07806_ ) );
OAI21_X1 _15851_ ( .A(_06858_ ), .B1(_05028_ ), .B2(_05029_ ), .ZN(_07807_ ) );
AOI21_X1 _15852_ ( .A(_07807_ ), .B1(_05029_ ), .B2(_05028_ ), .ZN(_07808_ ) );
OAI22_X1 _15853_ ( .A1(_05793_ ), .A2(_06861_ ), .B1(_02465_ ), .B2(_06566_ ), .ZN(_07809_ ) );
OAI21_X1 _15854_ ( .A(_06582_ ), .B1(_07808_ ), .B2(_07809_ ), .ZN(_07810_ ) );
NAND2_X1 _15855_ ( .A1(_07810_ ), .A2(_05347_ ), .ZN(_07811_ ) );
NAND2_X1 _15856_ ( .A1(_07097_ ), .A2(_06996_ ), .ZN(_07812_ ) );
NOR4_X1 _15857_ ( .A1(_07812_ ), .A2(_07516_ ), .A3(_06771_ ), .A4(_07621_ ), .ZN(_07813_ ) );
NAND2_X1 _15858_ ( .A1(_07127_ ), .A2(_07032_ ), .ZN(_07814_ ) );
OAI21_X1 _15859_ ( .A(_07017_ ), .B1(_06834_ ), .B2(_06830_ ), .ZN(_07815_ ) );
OAI211_X1 _15860_ ( .A(_07815_ ), .B(_07014_ ), .C1(_07017_ ), .C2(_07721_ ), .ZN(_07816_ ) );
OAI211_X1 _15861_ ( .A(_07025_ ), .B(_07816_ ), .C1(_07666_ ), .C2(_06868_ ), .ZN(_07817_ ) );
OAI211_X1 _15862_ ( .A(_07817_ ), .B(_07174_ ), .C1(_07001_ ), .C2(_07524_ ), .ZN(_07818_ ) );
NAND2_X1 _15863_ ( .A1(_07814_ ), .A2(_07818_ ), .ZN(_07819_ ) );
OAI21_X1 _15864_ ( .A(_06865_ ), .B1(_07813_ ), .B2(_07819_ ), .ZN(_07820_ ) );
OAI21_X1 _15865_ ( .A(_07221_ ), .B1(_04866_ ), .B2(_06619_ ), .ZN(_07821_ ) );
OR2_X1 _15866_ ( .A1(_07821_ ), .A2(_06621_ ), .ZN(_07822_ ) );
NAND2_X1 _15867_ ( .A1(_07819_ ), .A2(_06711_ ), .ZN(_07823_ ) );
NAND3_X1 _15868_ ( .A1(_07143_ ), .A2(_07001_ ), .A3(_07248_ ), .ZN(_07824_ ) );
OR2_X1 _15869_ ( .A1(_04865_ ), .A2(_06713_ ), .ZN(_07825_ ) );
AOI22_X1 _15870_ ( .A1(_04866_ ), .A2(_07042_ ), .B1(_04864_ ), .B2(_07092_ ), .ZN(_07826_ ) );
AND4_X1 _15871_ ( .A1(_07823_ ), .A2(_07824_ ), .A3(_07825_ ), .A4(_07826_ ), .ZN(_07827_ ) );
NAND3_X1 _15872_ ( .A1(_07820_ ), .A2(_07822_ ), .A3(_07827_ ), .ZN(_07828_ ) );
AOI21_X1 _15873_ ( .A(_07811_ ), .B1(_07828_ ), .B2(_07506_ ), .ZN(_07829_ ) );
OAI21_X1 _15874_ ( .A(_07765_ ), .B1(_05325_ ), .B2(\ID_EX_pc [1] ), .ZN(_07830_ ) );
OAI21_X1 _15875_ ( .A(_07806_ ), .B1(_07829_ ), .B2(_07830_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_30_D ) );
AND3_X1 _15876_ ( .A1(_05824_ ), .A2(_05825_ ), .A3(_05823_ ), .ZN(_07831_ ) );
AOI21_X1 _15877_ ( .A(_05778_ ), .B1(_07831_ ), .B2(_05822_ ), .ZN(_07832_ ) );
AND3_X1 _15878_ ( .A1(_05840_ ), .A2(_05841_ ), .A3(\EX_LS_result_csreg_mem [0] ), .ZN(_07833_ ) );
OAI21_X1 _15879_ ( .A(_06556_ ), .B1(_07832_ ), .B2(_07833_ ), .ZN(_07834_ ) );
AND3_X1 _15880_ ( .A1(_04764_ ), .A2(_06848_ ), .A3(_04787_ ), .ZN(_07835_ ) );
AND4_X1 _15881_ ( .A1(\ID_EX_typ [4] ), .A2(_03913_ ), .A3(\ID_EX_typ [3] ), .A4(_04769_ ), .ZN(_07836_ ) );
OAI21_X1 _15882_ ( .A(_05102_ ), .B1(_07835_ ), .B2(_07836_ ), .ZN(_07837_ ) );
AOI22_X1 _15883_ ( .A1(_04354_ ), .A2(_06974_ ), .B1(\ID_EX_imm [0] ), .B2(_07206_ ), .ZN(_07838_ ) );
NAND2_X1 _15884_ ( .A1(_07837_ ), .A2(_07838_ ), .ZN(_07839_ ) );
AND3_X1 _15885_ ( .A1(_05831_ ), .A2(_06559_ ), .A3(_06558_ ), .ZN(_07840_ ) );
OAI21_X1 _15886_ ( .A(_06582_ ), .B1(_07839_ ), .B2(_07840_ ), .ZN(_07841_ ) );
INV_X1 _15887_ ( .A(_05017_ ), .ZN(_07842_ ) );
NAND3_X1 _15888_ ( .A1(_04767_ ), .A2(_03877_ ), .A3(\ID_EX_typ [2] ), .ZN(_07843_ ) );
AOI221_X4 _15889_ ( .A(_07843_ ), .B1(_02990_ ), .B2(_05006_ ), .C1(_05021_ ), .C2(_05014_ ), .ZN(_07844_ ) );
NAND3_X1 _15890_ ( .A1(_05015_ ), .A2(_07842_ ), .A3(_07844_ ), .ZN(_07845_ ) );
NAND4_X1 _15891_ ( .A1(_07097_ ), .A2(_04900_ ), .A3(_06865_ ), .A4(_06761_ ), .ZN(_07846_ ) );
OAI21_X1 _15892_ ( .A(_06589_ ), .B1(_06952_ ), .B2(_04870_ ), .ZN(_07847_ ) );
NOR2_X1 _15893_ ( .A1(_07749_ ), .A2(_06951_ ), .ZN(_07848_ ) );
MUX2_X1 _15894_ ( .A(_04236_ ), .B(_06479_ ), .S(_06768_ ), .Z(_07849_ ) );
AOI211_X1 _15895_ ( .A(_06682_ ), .B(_07848_ ), .C1(_07017_ ), .C2(_07849_ ), .ZN(_07850_ ) );
AOI211_X1 _15896_ ( .A(_06814_ ), .B(_07850_ ), .C1(_07008_ ), .C2(_07691_ ), .ZN(_07851_ ) );
NOR3_X1 _15897_ ( .A1(_07553_ ), .A2(_07554_ ), .A3(_06704_ ), .ZN(_07852_ ) );
OAI21_X1 _15898_ ( .A(_06707_ ), .B1(_07851_ ), .B2(_07852_ ), .ZN(_07853_ ) );
OAI211_X1 _15899_ ( .A(_07853_ ), .B(_07237_ ), .C1(_07000_ ), .C2(_07173_ ), .ZN(_07854_ ) );
OAI21_X1 _15900_ ( .A(_04770_ ), .B1(_06664_ ), .B2(_04331_ ), .ZN(_07855_ ) );
NAND3_X1 _15901_ ( .A1(_07186_ ), .A2(_07063_ ), .A3(_07248_ ), .ZN(_07856_ ) );
OAI21_X1 _15902_ ( .A(_05025_ ), .B1(_06952_ ), .B2(_04870_ ), .ZN(_07857_ ) );
NAND3_X1 _15903_ ( .A1(_06664_ ), .A2(_04331_ ), .A3(_06586_ ), .ZN(_07858_ ) );
AND3_X1 _15904_ ( .A1(_07856_ ), .A2(_07857_ ), .A3(_07858_ ), .ZN(_07859_ ) );
AND4_X1 _15905_ ( .A1(_07847_ ), .A2(_07854_ ), .A3(_07855_ ), .A4(_07859_ ), .ZN(_07860_ ) );
NAND3_X1 _15906_ ( .A1(_07845_ ), .A2(_07846_ ), .A3(_07860_ ), .ZN(_07861_ ) );
AOI21_X1 _15907_ ( .A(_03892_ ), .B1(_07861_ ), .B2(_06852_ ), .ZN(_07862_ ) );
AND2_X1 _15908_ ( .A1(_07841_ ), .A2(_07862_ ), .ZN(_07863_ ) );
OAI21_X1 _15909_ ( .A(_07765_ ), .B1(_05325_ ), .B2(\ID_EX_pc [0] ), .ZN(_07864_ ) );
OAI21_X1 _15910_ ( .A(_07834_ ), .B1(_07863_ ), .B2(_07864_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_31_D ) );
NOR2_X1 _15911_ ( .A1(_05600_ ), .A2(_05598_ ), .ZN(_07865_ ) );
NAND4_X1 _15912_ ( .A1(_07865_ ), .A2(_05293_ ), .A3(_05719_ ), .A4(_05597_ ), .ZN(_07866_ ) );
INV_X1 _15913_ ( .A(\EX_LS_result_csreg_mem [28] ), .ZN(_07867_ ) );
NAND3_X1 _15914_ ( .A1(_05840_ ), .A2(_05841_ ), .A3(_07867_ ), .ZN(_07868_ ) );
NAND3_X1 _15915_ ( .A1(_07866_ ), .A2(_07868_ ), .A3(_06434_ ), .ZN(_07869_ ) );
AND2_X1 _15916_ ( .A1(_05593_ ), .A2(_07205_ ), .ZN(_07870_ ) );
OAI21_X1 _15917_ ( .A(_06858_ ), .B1(_07371_ ), .B2(_07372_ ), .ZN(_07871_ ) );
AOI21_X1 _15918_ ( .A(_07871_ ), .B1(_07372_ ), .B2(_07371_ ), .ZN(_07872_ ) );
AND3_X1 _15919_ ( .A1(_06562_ ), .A2(\ID_EX_imm [28] ), .A3(_06559_ ), .ZN(_07873_ ) );
NOR3_X1 _15920_ ( .A1(_07870_ ), .A2(_07872_ ), .A3(_07873_ ), .ZN(_07874_ ) );
OAI21_X1 _15921_ ( .A(_05928_ ), .B1(_07874_ ), .B2(_06584_ ), .ZN(_07875_ ) );
NOR3_X1 _15922_ ( .A1(_07417_ ), .A2(_04779_ ), .A3(_07419_ ), .ZN(_07876_ ) );
OR3_X1 _15923_ ( .A1(_07768_ ), .A2(_06905_ ), .A3(_07876_ ), .ZN(_07877_ ) );
NAND2_X1 _15924_ ( .A1(_04779_ ), .A2(_07042_ ), .ZN(_07878_ ) );
OAI21_X1 _15925_ ( .A(_06959_ ), .B1(_04777_ ), .B2(_02167_ ), .ZN(_07879_ ) );
NAND3_X1 _15926_ ( .A1(_04777_ ), .A2(_02167_ ), .A3(_07092_ ), .ZN(_07880_ ) );
AND3_X1 _15927_ ( .A1(_07878_ ), .A2(_07879_ ), .A3(_07880_ ), .ZN(_07881_ ) );
OAI21_X1 _15928_ ( .A(_06901_ ), .B1(_06916_ ), .B2(_06922_ ), .ZN(_07882_ ) );
OAI21_X1 _15929_ ( .A(_07011_ ), .B1(_06878_ ), .B2(_06890_ ), .ZN(_07883_ ) );
OAI211_X1 _15930_ ( .A(_07004_ ), .B(_07005_ ), .C1(_06886_ ), .C2(_06891_ ), .ZN(_07884_ ) );
AND2_X1 _15931_ ( .A1(_07883_ ), .A2(_07884_ ), .ZN(_07885_ ) );
NOR2_X1 _15932_ ( .A1(_06881_ ), .A2(_06879_ ), .ZN(_07886_ ) );
MUX2_X1 _15933_ ( .A(_07886_ ), .B(_07389_ ), .S(_07017_ ), .Z(_07887_ ) );
MUX2_X1 _15934_ ( .A(_07885_ ), .B(_07887_ ), .S(_06868_ ), .Z(_07888_ ) );
OAI211_X1 _15935_ ( .A(_07000_ ), .B(_07882_ ), .C1(_07888_ ), .C2(_07229_ ), .ZN(_07889_ ) );
OAI21_X1 _15936_ ( .A(_07032_ ), .B1(_07358_ ), .B2(_07359_ ), .ZN(_07890_ ) );
AOI21_X1 _15937_ ( .A(_06776_ ), .B1(_07889_ ), .B2(_07890_ ), .ZN(_07891_ ) );
AND3_X1 _15938_ ( .A1(_07351_ ), .A2(_06708_ ), .A3(_06710_ ), .ZN(_07892_ ) );
NAND2_X1 _15939_ ( .A1(_07351_ ), .A2(_06708_ ), .ZN(_07893_ ) );
NAND3_X1 _15940_ ( .A1(_07097_ ), .A2(_06765_ ), .A3(_07342_ ), .ZN(_07894_ ) );
OAI211_X1 _15941_ ( .A(_07893_ ), .B(_07894_ ), .C1(_06873_ ), .C2(_06872_ ), .ZN(_07895_ ) );
AOI211_X1 _15942_ ( .A(_07891_ ), .B(_07892_ ), .C1(_07895_ ), .C2(_06865_ ), .ZN(_07896_ ) );
NAND3_X1 _15943_ ( .A1(_07877_ ), .A2(_07881_ ), .A3(_07896_ ), .ZN(_07897_ ) );
AOI21_X1 _15944_ ( .A(_07875_ ), .B1(_07897_ ), .B2(_07506_ ), .ZN(_07898_ ) );
OAI21_X1 _15945_ ( .A(_07765_ ), .B1(_05590_ ), .B2(_07542_ ), .ZN(_07899_ ) );
OAI21_X1 _15946_ ( .A(_07869_ ), .B1(_07898_ ), .B2(_07899_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_3_D ) );
NAND3_X1 _15947_ ( .A1(_05814_ ), .A2(_05816_ ), .A3(_06434_ ), .ZN(_07900_ ) );
OAI22_X1 _15948_ ( .A1(_05806_ ), .A2(_06561_ ), .B1(_02200_ ), .B2(_06565_ ), .ZN(_07901_ ) );
OAI21_X1 _15949_ ( .A(_04760_ ), .B1(_07369_ ), .B2(_05096_ ), .ZN(_07902_ ) );
NAND3_X1 _15950_ ( .A1(_07902_ ), .A2(_04758_ ), .A3(_05069_ ), .ZN(_07903_ ) );
AOI21_X1 _15951_ ( .A(_05072_ ), .B1(_07903_ ), .B2(_04685_ ), .ZN(_07904_ ) );
XNOR2_X1 _15952_ ( .A(_04706_ ), .B(_04708_ ), .ZN(_07905_ ) );
OR2_X1 _15953_ ( .A1(_07904_ ), .A2(_07905_ ), .ZN(_07906_ ) );
AOI21_X1 _15954_ ( .A(_06576_ ), .B1(_07904_ ), .B2(_07905_ ), .ZN(_07907_ ) );
AOI21_X1 _15955_ ( .A(_07901_ ), .B1(_07906_ ), .B2(_07907_ ), .ZN(_07908_ ) );
OAI21_X1 _15956_ ( .A(_05928_ ), .B1(_07908_ ), .B2(_06584_ ), .ZN(_07909_ ) );
AOI21_X1 _15957_ ( .A(_04795_ ), .B1(_07414_ ), .B2(_07416_ ), .ZN(_07910_ ) );
OR3_X1 _15958_ ( .A1(_07910_ ), .A2(_04801_ ), .A3(_04792_ ), .ZN(_07911_ ) );
OAI21_X1 _15959_ ( .A(_04801_ ), .B1(_07910_ ), .B2(_04792_ ), .ZN(_07912_ ) );
AND3_X1 _15960_ ( .A1(_07911_ ), .A2(_07221_ ), .A3(_07912_ ), .ZN(_07913_ ) );
AOI22_X1 _15961_ ( .A1(_06763_ ), .A2(_06766_ ), .B1(_07000_ ), .B2(_07453_ ), .ZN(_07914_ ) );
OAI211_X1 _15962_ ( .A(_07097_ ), .B(_06765_ ), .C1(_06867_ ), .C2(_06996_ ), .ZN(_07915_ ) );
AOI21_X1 _15963_ ( .A(_06718_ ), .B1(_07914_ ), .B2(_07915_ ), .ZN(_07916_ ) );
NAND3_X1 _15964_ ( .A1(_07778_ ), .A2(_06819_ ), .A3(_06820_ ), .ZN(_07917_ ) );
NAND3_X1 _15965_ ( .A1(_06815_ ), .A2(_06680_ ), .A3(_06688_ ), .ZN(_07918_ ) );
NAND2_X1 _15966_ ( .A1(_07917_ ), .A2(_07918_ ), .ZN(_07919_ ) );
OAI21_X1 _15967_ ( .A(_06797_ ), .B1(_06698_ ), .B2(_06695_ ), .ZN(_07920_ ) );
OAI211_X1 _15968_ ( .A(_06689_ ), .B(_06690_ ), .C1(_06816_ ), .C2(_06694_ ), .ZN(_07921_ ) );
AND2_X1 _15969_ ( .A1(_07920_ ), .A2(_07921_ ), .ZN(_07922_ ) );
MUX2_X1 _15970_ ( .A(_07919_ ), .B(_07922_ ), .S(_06682_ ), .Z(_07923_ ) );
OR2_X1 _15971_ ( .A1(_07923_ ), .A2(_06839_ ), .ZN(_07924_ ) );
NAND3_X1 _15972_ ( .A1(_07021_ ), .A2(_07024_ ), .A3(_07228_ ), .ZN(_07925_ ) );
NAND3_X1 _15973_ ( .A1(_07924_ ), .A2(_07248_ ), .A3(_07925_ ), .ZN(_07926_ ) );
AOI22_X1 _15974_ ( .A1(_04801_ ), .A2(_05025_ ), .B1(_04799_ ), .B2(_06586_ ), .ZN(_07927_ ) );
OAI211_X1 _15975_ ( .A(_07926_ ), .B(_07927_ ), .C1(_04800_ ), .C2(_06713_ ), .ZN(_07928_ ) );
NOR2_X1 _15976_ ( .A1(_06943_ ), .A2(_06776_ ), .ZN(_07929_ ) );
INV_X1 _15977_ ( .A(_07929_ ), .ZN(_07930_ ) );
AOI21_X1 _15978_ ( .A(_07930_ ), .B1(_07458_ ), .B2(_07459_ ), .ZN(_07931_ ) );
AND3_X1 _15979_ ( .A1(_07453_ ), .A2(_06707_ ), .A3(_06709_ ), .ZN(_07932_ ) );
OR3_X1 _15980_ ( .A1(_07928_ ), .A2(_07931_ ), .A3(_07932_ ), .ZN(_07933_ ) );
OR3_X1 _15981_ ( .A1(_07913_ ), .A2(_07916_ ), .A3(_07933_ ), .ZN(_07934_ ) );
AOI21_X1 _15982_ ( .A(_07909_ ), .B1(_07934_ ), .B2(_07506_ ), .ZN(_07935_ ) );
NAND2_X1 _15983_ ( .A1(_05801_ ), .A2(_03892_ ), .ZN(_07936_ ) );
NAND2_X1 _15984_ ( .A1(_07936_ ), .A2(_06422_ ), .ZN(_07937_ ) );
OAI21_X1 _15985_ ( .A(_07900_ ), .B1(_07935_ ), .B2(_07937_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_4_D ) );
AND2_X1 _15986_ ( .A1(_05844_ ), .A2(_05843_ ), .ZN(_07938_ ) );
AND2_X1 _15987_ ( .A1(_05845_ ), .A2(_05846_ ), .ZN(_07939_ ) );
AOI21_X1 _15988_ ( .A(_05778_ ), .B1(_07938_ ), .B2(_07939_ ), .ZN(_07940_ ) );
AND3_X1 _15989_ ( .A1(_05840_ ), .A2(_05841_ ), .A3(\EX_LS_result_csreg_mem [26] ), .ZN(_07941_ ) );
OAI21_X1 _15990_ ( .A(_06556_ ), .B1(_07940_ ), .B2(_07941_ ), .ZN(_07942_ ) );
OAI22_X1 _15991_ ( .A1(_05838_ ), .A2(_06561_ ), .B1(_02197_ ), .B2(_06565_ ), .ZN(_07943_ ) );
OR2_X1 _15992_ ( .A1(_07903_ ), .A2(_04685_ ), .ZN(_07944_ ) );
AOI21_X1 _15993_ ( .A(_06576_ ), .B1(_07903_ ), .B2(_04685_ ), .ZN(_07945_ ) );
AOI21_X1 _15994_ ( .A(_07943_ ), .B1(_07944_ ), .B2(_07945_ ), .ZN(_07946_ ) );
OAI21_X1 _15995_ ( .A(_05928_ ), .B1(_07946_ ), .B2(_06584_ ), .ZN(_07947_ ) );
AND3_X1 _15996_ ( .A1(_07414_ ), .A2(_04795_ ), .A3(_07416_ ), .ZN(_07948_ ) );
OR3_X1 _15997_ ( .A1(_07948_ ), .A2(_07910_ ), .A3(_06905_ ), .ZN(_07949_ ) );
AND3_X1 _15998_ ( .A1(_07500_ ), .A2(_07501_ ), .A3(_07929_ ), .ZN(_07950_ ) );
AND2_X1 _15999_ ( .A1(_07492_ ), .A2(_06838_ ), .ZN(_07951_ ) );
OR2_X1 _16000_ ( .A1(_06977_ ), .A2(_07951_ ), .ZN(_07952_ ) );
INV_X1 _16001_ ( .A(_07481_ ), .ZN(_07953_ ) );
INV_X1 _16002_ ( .A(_07483_ ), .ZN(_07954_ ) );
AOI21_X1 _16003_ ( .A(_06874_ ), .B1(_07953_ ), .B2(_07954_ ), .ZN(_07955_ ) );
OAI21_X1 _16004_ ( .A(_06716_ ), .B1(_07952_ ), .B2(_07955_ ), .ZN(_07956_ ) );
NAND3_X1 _16005_ ( .A1(_07492_ ), .A2(_06708_ ), .A3(_06710_ ), .ZN(_07957_ ) );
NAND2_X1 _16006_ ( .A1(_07956_ ), .A2(_07957_ ), .ZN(_07958_ ) );
NAND2_X1 _16007_ ( .A1(_07088_ ), .A2(_07229_ ), .ZN(_07959_ ) );
NOR2_X1 _16008_ ( .A1(_07393_ ), .A2(_07394_ ), .ZN(_07960_ ) );
MUX2_X1 _16009_ ( .A(_07387_ ), .B(_07960_ ), .S(_07008_ ), .Z(_07961_ ) );
AOI21_X1 _16010_ ( .A(_07457_ ), .B1(_07961_ ), .B2(_07001_ ), .ZN(_07962_ ) );
AOI211_X1 _16011_ ( .A(_07950_ ), .B(_07958_ ), .C1(_07959_ ), .C2(_07962_ ), .ZN(_07963_ ) );
NOR3_X1 _16012_ ( .A1(_04792_ ), .A2(_04793_ ), .A3(_05026_ ), .ZN(_07964_ ) );
NOR3_X1 _16013_ ( .A1(_04790_ ), .A2(_04791_ ), .A3(_06843_ ), .ZN(_07965_ ) );
AOI21_X1 _16014_ ( .A(_06713_ ), .B1(_04790_ ), .B2(_04791_ ), .ZN(_07966_ ) );
NOR3_X1 _16015_ ( .A1(_07964_ ), .A2(_07965_ ), .A3(_07966_ ), .ZN(_07967_ ) );
NAND3_X1 _16016_ ( .A1(_07949_ ), .A2(_07963_ ), .A3(_07967_ ), .ZN(_07968_ ) );
AOI21_X1 _16017_ ( .A(_07947_ ), .B1(_07968_ ), .B2(_07506_ ), .ZN(_07969_ ) );
OAI21_X1 _16018_ ( .A(_07765_ ), .B1(_05835_ ), .B2(_07542_ ), .ZN(_07970_ ) );
OAI21_X1 _16019_ ( .A(_07942_ ), .B1(_07969_ ), .B2(_07970_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_5_D ) );
OR2_X1 _16020_ ( .A1(_06507_ ), .A2(_06213_ ), .ZN(_07971_ ) );
NOR2_X1 _16021_ ( .A1(_07369_ ), .A2(_05096_ ), .ZN(_07972_ ) );
INV_X1 _16022_ ( .A(_04734_ ), .ZN(_00304_ ) );
NOR2_X1 _16023_ ( .A1(_07972_ ), .A2(_00304_ ), .ZN(_00305_ ) );
OR3_X1 _16024_ ( .A1(_00305_ ), .A2(_04759_ ), .A3(_05068_ ), .ZN(_00306_ ) );
OAI21_X1 _16025_ ( .A(_04759_ ), .B1(_00305_ ), .B2(_05068_ ), .ZN(_00307_ ) );
AND3_X1 _16026_ ( .A1(_00306_ ), .A2(_06858_ ), .A3(_00307_ ), .ZN(_00308_ ) );
OAI22_X1 _16027_ ( .A1(_05864_ ), .A2(_06861_ ), .B1(_02900_ ), .B2(_06566_ ), .ZN(_00309_ ) );
OAI21_X1 _16028_ ( .A(_06582_ ), .B1(_00308_ ), .B2(_00309_ ), .ZN(_00310_ ) );
NAND2_X1 _16029_ ( .A1(_00310_ ), .A2(_05347_ ), .ZN(_00311_ ) );
NAND2_X1 _16030_ ( .A1(_07413_ ), .A2(_04810_ ), .ZN(_00312_ ) );
INV_X1 _16031_ ( .A(_04808_ ), .ZN(_00313_ ) );
INV_X1 _16032_ ( .A(_04816_ ), .ZN(_00314_ ) );
AND3_X1 _16033_ ( .A1(_00312_ ), .A2(_00313_ ), .A3(_00314_ ), .ZN(_00315_ ) );
AOI21_X1 _16034_ ( .A(_00314_ ), .B1(_00312_ ), .B2(_00313_ ), .ZN(_00316_ ) );
NOR3_X1 _16035_ ( .A1(_00315_ ), .A2(_00316_ ), .A3(_06905_ ), .ZN(_00317_ ) );
AOI22_X1 _16036_ ( .A1(_07415_ ), .A2(_06959_ ), .B1(_04814_ ), .B2(_07092_ ), .ZN(_00318_ ) );
OAI21_X1 _16037_ ( .A(_00318_ ), .B1(_00314_ ), .B2(_05026_ ), .ZN(_00319_ ) );
OAI21_X1 _16038_ ( .A(_06765_ ), .B1(_07481_ ), .B2(_07517_ ), .ZN(_00320_ ) );
AND3_X1 _16039_ ( .A1(_07119_ ), .A2(_06702_ ), .A3(_07120_ ), .ZN(_00321_ ) );
AND2_X1 _16040_ ( .A1(_00321_ ), .A2(_06943_ ), .ZN(_00322_ ) );
AOI21_X1 _16041_ ( .A(_00322_ ), .B1(_06763_ ), .B2(_06764_ ), .ZN(_00323_ ) );
AOI21_X1 _16042_ ( .A(_06717_ ), .B1(_00320_ ), .B2(_00323_ ), .ZN(_00324_ ) );
AOI21_X1 _16043_ ( .A(_07930_ ), .B1(_07530_ ), .B2(_07531_ ), .ZN(_00325_ ) );
AND3_X1 _16044_ ( .A1(_00321_ ), .A2(_06838_ ), .A3(_06709_ ), .ZN(_00326_ ) );
OR2_X1 _16045_ ( .A1(_07141_ ), .A2(_06703_ ), .ZN(_00327_ ) );
NOR2_X1 _16046_ ( .A1(_07779_ ), .A2(_06677_ ), .ZN(_00328_ ) );
AOI21_X1 _16047_ ( .A(_06805_ ), .B1(_06817_ ), .B2(_06823_ ), .ZN(_00329_ ) );
OAI21_X1 _16048_ ( .A(_06704_ ), .B1(_00328_ ), .B2(_00329_ ), .ZN(_00330_ ) );
AND3_X1 _16049_ ( .A1(_00327_ ), .A2(_07247_ ), .A3(_00330_ ), .ZN(_00331_ ) );
OR4_X1 _16050_ ( .A1(_00324_ ), .A2(_00325_ ), .A3(_00326_ ), .A4(_00331_ ), .ZN(_00332_ ) );
OR3_X1 _16051_ ( .A1(_00317_ ), .A2(_00319_ ), .A3(_00332_ ), .ZN(_00333_ ) );
AOI21_X1 _16052_ ( .A(_00311_ ), .B1(_00333_ ), .B2(_06852_ ), .ZN(_00334_ ) );
OAI21_X1 _16053_ ( .A(_07765_ ), .B1(_05859_ ), .B2(_07542_ ), .ZN(_00335_ ) );
OAI21_X1 _16054_ ( .A(_07971_ ), .B1(_00334_ ), .B2(_00335_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_6_D ) );
OAI211_X1 _16055_ ( .A(_06515_ ), .B(_06333_ ), .C1(_06516_ ), .C2(_06517_ ), .ZN(_00336_ ) );
OAI21_X1 _16056_ ( .A(_06858_ ), .B1(_07972_ ), .B2(_00304_ ), .ZN(_00337_ ) );
AOI21_X1 _16057_ ( .A(_00337_ ), .B1(_00304_ ), .B2(_07972_ ), .ZN(_00338_ ) );
OAI22_X1 _16058_ ( .A1(_05880_ ), .A2(_06861_ ), .B1(_02877_ ), .B2(_06566_ ), .ZN(_00339_ ) );
OAI21_X1 _16059_ ( .A(_06582_ ), .B1(_00338_ ), .B2(_00339_ ), .ZN(_00340_ ) );
NAND2_X1 _16060_ ( .A1(_00340_ ), .A2(_05928_ ), .ZN(_00341_ ) );
OAI21_X1 _16061_ ( .A(_06589_ ), .B1(_07413_ ), .B2(_04810_ ), .ZN(_00342_ ) );
AOI21_X1 _16062_ ( .A(_00342_ ), .B1(_04810_ ), .B2(_07413_ ), .ZN(_00343_ ) );
NOR3_X1 _16063_ ( .A1(_04808_ ), .A2(_04809_ ), .A3(_05026_ ), .ZN(_00344_ ) );
NOR3_X1 _16064_ ( .A1(_04806_ ), .A2(_04807_ ), .A3(_06843_ ), .ZN(_00345_ ) );
AOI21_X1 _16065_ ( .A(_04771_ ), .B1(_04806_ ), .B2(_04807_ ), .ZN(_00346_ ) );
OR3_X1 _16066_ ( .A1(_00344_ ), .A2(_00345_ ), .A3(_00346_ ), .ZN(_00347_ ) );
OAI211_X1 _16067_ ( .A(_06760_ ), .B(_06765_ ), .C1(_06901_ ), .C2(_06721_ ), .ZN(_00348_ ) );
NOR2_X1 _16068_ ( .A1(_07172_ ), .A2(_07228_ ), .ZN(_00349_ ) );
INV_X1 _16069_ ( .A(_00349_ ), .ZN(_00350_ ) );
OAI21_X1 _16070_ ( .A(_00348_ ), .B1(_07032_ ), .B2(_00350_ ), .ZN(_00351_ ) );
OAI21_X1 _16071_ ( .A(_06716_ ), .B1(_06977_ ), .B2(_00351_ ), .ZN(_00352_ ) );
NAND3_X1 _16072_ ( .A1(_07561_ ), .A2(_07562_ ), .A3(_07929_ ), .ZN(_00353_ ) );
NAND2_X1 _16073_ ( .A1(_07179_ ), .A2(_07180_ ), .ZN(_00354_ ) );
NAND2_X1 _16074_ ( .A1(_00354_ ), .A2(_07229_ ), .ZN(_00355_ ) );
AOI21_X1 _16075_ ( .A(_06868_ ), .B1(_06918_ ), .B2(_06921_ ), .ZN(_00356_ ) );
AOI21_X1 _16076_ ( .A(_07008_ ), .B1(_07883_ ), .B2(_07884_ ), .ZN(_00357_ ) );
OAI21_X1 _16077_ ( .A(_07001_ ), .B1(_00356_ ), .B2(_00357_ ), .ZN(_00358_ ) );
NAND3_X1 _16078_ ( .A1(_00355_ ), .A2(_07248_ ), .A3(_00358_ ), .ZN(_00359_ ) );
NAND3_X1 _16079_ ( .A1(_00349_ ), .A2(_07000_ ), .A3(_06710_ ), .ZN(_00360_ ) );
NAND4_X1 _16080_ ( .A1(_00352_ ), .A2(_00353_ ), .A3(_00359_ ), .A4(_00360_ ), .ZN(_00361_ ) );
OR3_X1 _16081_ ( .A1(_00343_ ), .A2(_00347_ ), .A3(_00361_ ), .ZN(_00362_ ) );
AOI21_X1 _16082_ ( .A(_00341_ ), .B1(_00362_ ), .B2(_06852_ ), .ZN(_00363_ ) );
OAI21_X1 _16083_ ( .A(_07765_ ), .B1(_05877_ ), .B2(_07542_ ), .ZN(_00364_ ) );
OAI21_X1 _16084_ ( .A(_00336_ ), .B1(_00363_ ), .B2(_00364_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_7_D ) );
AND2_X1 _16085_ ( .A1(_05904_ ), .A2(_05903_ ), .ZN(_00365_ ) );
AND2_X1 _16086_ ( .A1(_05905_ ), .A2(_05906_ ), .ZN(_00366_ ) );
AOI21_X1 _16087_ ( .A(_05778_ ), .B1(_00365_ ), .B2(_00366_ ), .ZN(_00367_ ) );
AND3_X1 _16088_ ( .A1(_05840_ ), .A2(_05841_ ), .A3(\EX_LS_result_csreg_mem [23] ), .ZN(_00368_ ) );
OAI21_X1 _16089_ ( .A(_06556_ ), .B1(_00367_ ), .B2(_00368_ ), .ZN(_00369_ ) );
NOR4_X1 _16090_ ( .A1(_06569_ ), .A2(_04488_ ), .A3(_04512_ ), .A4(_04513_ ), .ZN(_00370_ ) );
OR2_X1 _16091_ ( .A1(_00370_ ), .A2(_05089_ ), .ZN(_00371_ ) );
AND2_X1 _16092_ ( .A1(_00371_ ), .A2(_04562_ ), .ZN(_00372_ ) );
OR3_X1 _16093_ ( .A1(_00372_ ), .A2(_04537_ ), .A3(_05093_ ), .ZN(_00373_ ) );
OAI21_X1 _16094_ ( .A(_04537_ ), .B1(_00372_ ), .B2(_05093_ ), .ZN(_00374_ ) );
NAND3_X1 _16095_ ( .A1(_00373_ ), .A2(_06974_ ), .A3(_00374_ ), .ZN(_00375_ ) );
NOR2_X1 _16096_ ( .A1(_05900_ ), .A2(_06861_ ), .ZN(_00376_ ) );
AOI21_X1 _16097_ ( .A(_00376_ ), .B1(\ID_EX_imm [23] ), .B2(_07206_ ), .ZN(_00377_ ) );
AOI21_X1 _16098_ ( .A(_06584_ ), .B1(_00375_ ), .B2(_00377_ ), .ZN(_00378_ ) );
NAND2_X1 _16099_ ( .A1(_06656_ ), .A2(_07404_ ), .ZN(_00379_ ) );
AOI21_X1 _16100_ ( .A(_07406_ ), .B1(_00379_ ), .B2(_07407_ ), .ZN(_00380_ ) );
NOR2_X1 _16101_ ( .A1(_04938_ ), .A2(_04538_ ), .ZN(_00381_ ) );
OR3_X1 _16102_ ( .A1(_00380_ ), .A2(_04946_ ), .A3(_00381_ ), .ZN(_00382_ ) );
OAI21_X1 _16103_ ( .A(_04946_ ), .B1(_00380_ ), .B2(_00381_ ), .ZN(_00383_ ) );
NAND3_X1 _16104_ ( .A1(_00382_ ), .A2(_07221_ ), .A3(_00383_ ), .ZN(_00384_ ) );
OAI211_X1 _16105_ ( .A(_06760_ ), .B(_06762_ ), .C1(_06766_ ), .C2(_06867_ ), .ZN(_00385_ ) );
NAND2_X1 _16106_ ( .A1(_07599_ ), .A2(_07174_ ), .ZN(_00386_ ) );
AOI21_X1 _16107_ ( .A(_06717_ ), .B1(_00385_ ), .B2(_00386_ ), .ZN(_00387_ ) );
AND3_X1 _16108_ ( .A1(_07599_ ), .A2(_06707_ ), .A3(_06710_ ), .ZN(_00388_ ) );
OR2_X1 _16109_ ( .A1(_00387_ ), .A2(_00388_ ), .ZN(_00389_ ) );
NOR3_X1 _16110_ ( .A1(_04942_ ), .A2(_04943_ ), .A3(_06843_ ), .ZN(_00390_ ) );
OAI22_X1 _16111_ ( .A1(_07408_ ), .A2(_05026_ ), .B1(_04945_ ), .B2(_06713_ ), .ZN(_00391_ ) );
OR3_X1 _16112_ ( .A1(_07242_ ), .A2(_06707_ ), .A3(_07228_ ), .ZN(_00392_ ) );
OAI21_X1 _16113_ ( .A(_06901_ ), .B1(_07244_ ), .B2(_07245_ ), .ZN(_00393_ ) );
AOI21_X1 _16114_ ( .A(_07008_ ), .B1(_07920_ ), .B2(_07921_ ), .ZN(_00394_ ) );
AOI21_X1 _16115_ ( .A(_07014_ ), .B1(_07022_ ), .B2(_07023_ ), .ZN(_00395_ ) );
NOR2_X1 _16116_ ( .A1(_00394_ ), .A2(_00395_ ), .ZN(_00396_ ) );
OAI211_X1 _16117_ ( .A(_00393_ ), .B(_07174_ ), .C1(_07229_ ), .C2(_00396_ ), .ZN(_00397_ ) );
AOI21_X1 _16118_ ( .A(_06776_ ), .B1(_00392_ ), .B2(_00397_ ), .ZN(_00398_ ) );
NOR4_X1 _16119_ ( .A1(_00389_ ), .A2(_00390_ ), .A3(_00391_ ), .A4(_00398_ ), .ZN(_00399_ ) );
AOI21_X1 _16120_ ( .A(_06851_ ), .B1(_00384_ ), .B2(_00399_ ), .ZN(_00400_ ) );
NOR3_X1 _16121_ ( .A1(_00378_ ), .A2(_05610_ ), .A3(_00400_ ), .ZN(_00401_ ) );
OAI21_X1 _16122_ ( .A(_07765_ ), .B1(_05894_ ), .B2(_07542_ ), .ZN(_00402_ ) );
OAI21_X1 _16123_ ( .A(_00369_ ), .B1(_00401_ ), .B2(_00402_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_8_D ) );
OR2_X1 _16124_ ( .A1(_06537_ ), .A2(_06213_ ), .ZN(_00403_ ) );
NOR3_X1 _16125_ ( .A1(_00370_ ), .A2(_04562_ ), .A3(_05089_ ), .ZN(_00404_ ) );
NOR3_X1 _16126_ ( .A1(_00372_ ), .A2(_00404_ ), .A3(_06576_ ), .ZN(_00405_ ) );
OAI22_X1 _16127_ ( .A1(_05917_ ), .A2(_06861_ ), .B1(_02271_ ), .B2(_06566_ ), .ZN(_00406_ ) );
OAI21_X1 _16128_ ( .A(_06582_ ), .B1(_00405_ ), .B2(_00406_ ), .ZN(_00407_ ) );
NAND2_X1 _16129_ ( .A1(_00407_ ), .A2(_05928_ ), .ZN(_00408_ ) );
AND2_X1 _16130_ ( .A1(_07623_ ), .A2(_06838_ ), .ZN(_00409_ ) );
NOR4_X1 _16131_ ( .A1(_07620_ ), .A2(_06771_ ), .A3(_06874_ ), .A4(_07265_ ), .ZN(_00410_ ) );
OR3_X1 _16132_ ( .A1(_06977_ ), .A2(_00409_ ), .A3(_00410_ ), .ZN(_00411_ ) );
NAND2_X1 _16133_ ( .A1(_00411_ ), .A2(_06716_ ), .ZN(_00412_ ) );
AOI21_X1 _16134_ ( .A(_07063_ ), .B1(_07287_ ), .B2(_07288_ ), .ZN(_00413_ ) );
AOI211_X1 _16135_ ( .A(_06877_ ), .B(_00413_ ), .C1(_07001_ ), .C2(_07396_ ), .ZN(_00414_ ) );
AOI211_X1 _16136_ ( .A(_07174_ ), .B(_06901_ ), .C1(_07290_ ), .C2(_07291_ ), .ZN(_00415_ ) );
OAI21_X1 _16137_ ( .A(_05099_ ), .B1(_00414_ ), .B2(_00415_ ), .ZN(_00416_ ) );
NAND3_X1 _16138_ ( .A1(_07623_ ), .A2(_06708_ ), .A3(_06711_ ), .ZN(_00417_ ) );
NAND3_X1 _16139_ ( .A1(_00412_ ), .A2(_00416_ ), .A3(_00417_ ), .ZN(_00418_ ) );
AND3_X1 _16140_ ( .A1(_00379_ ), .A2(_07406_ ), .A3(_07407_ ), .ZN(_00419_ ) );
NOR3_X1 _16141_ ( .A1(_00419_ ), .A2(_00380_ ), .A3(_06590_ ), .ZN(_00420_ ) );
NAND3_X1 _16142_ ( .A1(_04936_ ), .A2(_04538_ ), .A3(_04937_ ), .ZN(_00421_ ) );
AOI22_X1 _16143_ ( .A1(_00381_ ), .A2(_07092_ ), .B1(_00421_ ), .B2(_04770_ ), .ZN(_00422_ ) );
OAI21_X1 _16144_ ( .A(_00422_ ), .B1(_07406_ ), .B2(_05026_ ), .ZN(_00423_ ) );
OR3_X1 _16145_ ( .A1(_00418_ ), .A2(_00420_ ), .A3(_00423_ ), .ZN(_00424_ ) );
AOI21_X1 _16146_ ( .A(_00408_ ), .B1(_00424_ ), .B2(_06852_ ), .ZN(_00425_ ) );
OAI21_X1 _16147_ ( .A(_07765_ ), .B1(_05913_ ), .B2(_07542_ ), .ZN(_00426_ ) );
OAI21_X1 _16148_ ( .A(_00403_ ), .B1(_00425_ ), .B2(_00426_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_9_D ) );
AND2_X1 _16149_ ( .A1(_05965_ ), .A2(_05967_ ), .ZN(_00427_ ) );
AND2_X1 _16150_ ( .A1(_05966_ ), .A2(_05968_ ), .ZN(_00428_ ) );
AOI21_X1 _16151_ ( .A(_05778_ ), .B1(_00427_ ), .B2(_00428_ ), .ZN(_00429_ ) );
AND3_X1 _16152_ ( .A1(_05840_ ), .A2(_05841_ ), .A3(\EX_LS_result_csreg_mem [31] ), .ZN(_00430_ ) );
OAI21_X1 _16153_ ( .A(_06556_ ), .B1(_00429_ ), .B2(_00430_ ), .ZN(_00431_ ) );
INV_X1 _16154_ ( .A(_05013_ ), .ZN(_00432_ ) );
AOI21_X1 _16155_ ( .A(_00432_ ), .B1(_07422_ ), .B2(_07425_ ), .ZN(_00433_ ) );
INV_X1 _16156_ ( .A(_05012_ ), .ZN(_00434_ ) );
NOR2_X1 _16157_ ( .A1(_00434_ ), .A2(_02963_ ), .ZN(_00435_ ) );
OR3_X1 _16158_ ( .A1(_00433_ ), .A2(_05009_ ), .A3(_00435_ ), .ZN(_00436_ ) );
OAI21_X1 _16159_ ( .A(_05009_ ), .B1(_00433_ ), .B2(_00435_ ), .ZN(_00437_ ) );
NAND3_X1 _16160_ ( .A1(_00436_ ), .A2(_07221_ ), .A3(_00437_ ), .ZN(_00438_ ) );
AND2_X1 _16161_ ( .A1(_06761_ ), .A2(_02990_ ), .ZN(_00439_ ) );
OAI21_X1 _16162_ ( .A(_06716_ ), .B1(_06763_ ), .B2(_00439_ ), .ZN(_00440_ ) );
NAND3_X1 _16163_ ( .A1(_07243_ ), .A2(_07246_ ), .A3(_07929_ ), .ZN(_00441_ ) );
AOI221_X4 _16164_ ( .A(_06673_ ), .B1(_06888_ ), .B2(_06889_ ), .C1(_06341_ ), .C2(_06664_ ), .ZN(_00442_ ) );
AOI21_X1 _16165_ ( .A(_07011_ ), .B1(_06684_ ), .B2(_06667_ ), .ZN(_00443_ ) );
NOR2_X1 _16166_ ( .A1(_00442_ ), .A2(_00443_ ), .ZN(_00444_ ) );
MUX2_X1 _16167_ ( .A(_07919_ ), .B(_00444_ ), .S(_07014_ ), .Z(_00445_ ) );
MUX2_X1 _16168_ ( .A(_00396_ ), .B(_00445_ ), .S(_07025_ ), .Z(_00446_ ) );
NAND2_X1 _16169_ ( .A1(_00446_ ), .A2(_07248_ ), .ZN(_00447_ ) );
NAND3_X1 _16170_ ( .A1(_06761_ ), .A2(_02990_ ), .A3(_06710_ ), .ZN(_00448_ ) );
OAI21_X1 _16171_ ( .A(_04770_ ), .B1(_05018_ ), .B2(_02990_ ), .ZN(_00449_ ) );
NOR3_X1 _16172_ ( .A1(_05006_ ), .A2(_05007_ ), .A3(_04766_ ), .ZN(_00450_ ) );
AOI21_X1 _16173_ ( .A(_00450_ ), .B1(_05009_ ), .B2(_07041_ ), .ZN(_00451_ ) );
AND3_X1 _16174_ ( .A1(_00448_ ), .A2(_00449_ ), .A3(_00451_ ), .ZN(_00452_ ) );
AND4_X1 _16175_ ( .A1(_00440_ ), .A2(_00441_ ), .A3(_00447_ ), .A4(_00452_ ), .ZN(_00453_ ) );
AOI21_X1 _16176_ ( .A(_06851_ ), .B1(_00438_ ), .B2(_00453_ ), .ZN(_00454_ ) );
OR2_X1 _16177_ ( .A1(_05964_ ), .A2(_06861_ ), .ZN(_00455_ ) );
AOI21_X1 _16178_ ( .A(_05066_ ), .B1(_07374_ ), .B2(_04658_ ), .ZN(_00456_ ) );
XNOR2_X1 _16179_ ( .A(_00456_ ), .B(_04634_ ), .ZN(_00457_ ) );
AOI22_X1 _16180_ ( .A1(_00457_ ), .A2(_06974_ ), .B1(\ID_EX_imm [31] ), .B2(_07206_ ), .ZN(_00458_ ) );
AOI21_X1 _16181_ ( .A(_06584_ ), .B1(_00455_ ), .B2(_00458_ ), .ZN(_00459_ ) );
NOR3_X1 _16182_ ( .A1(_00454_ ), .A2(_05610_ ), .A3(_00459_ ), .ZN(_00460_ ) );
NAND2_X1 _16183_ ( .A1(_05976_ ), .A2(_03892_ ), .ZN(_00461_ ) );
NAND2_X1 _16184_ ( .A1(_00461_ ), .A2(_06422_ ), .ZN(_00462_ ) );
OAI21_X1 _16185_ ( .A(_00431_ ), .B1(_00460_ ), .B2(_00462_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_D ) );
AND3_X1 _16186_ ( .A1(\myexu.state_$_ANDNOT__B_Y ), .A2(_03083_ ), .A3(_03890_ ), .ZN(\myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ) );
AOI21_X1 _16187_ ( .A(_02081_ ), .B1(_02057_ ), .B2(_02088_ ), .ZN(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NAND2_X1 _16188_ ( .A1(_03365_ ), .A2(IDU_valid_EXU ), .ZN(_00463_ ) );
OAI21_X1 _16189_ ( .A(_00463_ ), .B1(_03303_ ), .B2(_03224_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _16190_ ( .A1(_03300_ ), .A2(_03224_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16191_ ( .A1(_03300_ ), .A2(_03224_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _16192_ ( .A(_03221_ ), .ZN(_00464_ ) );
NOR4_X1 _16193_ ( .A1(_03300_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03067_ ), .A4(_00464_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _16194_ ( .A1(_03618_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03067_ ), .A4(_03220_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ) );
AOI21_X1 _16195_ ( .A(_03827_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _16196_ ( .A(_00463_ ), .B1(_00464_ ), .B2(_03365_ ), .ZN(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ) );
OAI22_X1 _16197_ ( .A1(_03221_ ), .A2(_03365_ ), .B1(_01986_ ), .B2(_03872_ ), .ZN(_00465_ ) );
INV_X1 _16198_ ( .A(loaduse_clear ), .ZN(_00466_ ) );
AOI221_X4 _16199_ ( .A(_00465_ ), .B1(\myidu.state [2] ), .B2(_00466_ ), .C1(_03300_ ), .C2(_03827_ ), .ZN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ) );
NAND3_X1 _16200_ ( .A1(_03127_ ), .A2(IDU_valid_EXU ), .A3(_06000_ ), .ZN(_00467_ ) );
NAND3_X1 _16201_ ( .A1(_03127_ ), .A2(\myidu.state [2] ), .A3(loaduse_clear ), .ZN(_00468_ ) );
NAND2_X1 _16202_ ( .A1(_03222_ ), .A2(_03127_ ), .ZN(_00469_ ) );
AOI21_X1 _16203_ ( .A(_03359_ ), .B1(_03338_ ), .B2(_03062_ ), .ZN(_00470_ ) );
NAND3_X1 _16204_ ( .A1(_03284_ ), .A2(_03287_ ), .A3(_03296_ ), .ZN(_00471_ ) );
AND4_X1 _16205_ ( .A1(_03236_ ), .A2(_03241_ ), .A3(_03269_ ), .A4(_03272_ ), .ZN(_00472_ ) );
NAND3_X1 _16206_ ( .A1(_03262_ ), .A2(_00472_ ), .A3(_03371_ ), .ZN(_00473_ ) );
OAI21_X1 _16207_ ( .A(_03360_ ), .B1(_00471_ ), .B2(_00473_ ), .ZN(_00474_ ) );
INV_X1 _16208_ ( .A(_00474_ ), .ZN(_00475_ ) );
OR2_X1 _16209_ ( .A1(_00470_ ), .A2(_00475_ ), .ZN(_00476_ ) );
OAI211_X1 _16210_ ( .A(_00467_ ), .B(_00468_ ), .C1(_00469_ ), .C2(_00476_ ), .ZN(\myidu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _16211_ ( .A(_03127_ ), .B(_03873_ ), .C1(_03221_ ), .C2(_03365_ ), .ZN(\myidu.state_$_DFF_P__Q_2_D ) );
OAI211_X1 _16212_ ( .A(_03222_ ), .B(_03127_ ), .C1(_00475_ ), .C2(_00470_ ), .ZN(_00477_ ) );
NAND3_X1 _16213_ ( .A1(_03127_ ), .A2(\myidu.state [2] ), .A3(_00466_ ), .ZN(_00478_ ) );
NAND2_X1 _16214_ ( .A1(_00477_ ), .A2(_00478_ ), .ZN(\myidu.state_$_DFF_P__Q_D ) );
NOR2_X1 _16215_ ( .A1(_03218_ ), .A2(IDU_ready_IFU ), .ZN(_00479_ ) );
NOR2_X1 _16216_ ( .A1(_03218_ ), .A2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_00480_ ) );
NOR2_X1 _16217_ ( .A1(\myifu.state [0] ), .A2(\myifu.state [1] ), .ZN(_00481_ ) );
NOR4_X1 _16218_ ( .A1(_00479_ ), .A2(_00480_ ), .A3(reset ), .A4(_00481_ ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E ) );
OR3_X1 _16219_ ( .A1(_01951_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06070_ ), .ZN(_00482_ ) );
OAI211_X1 _16220_ ( .A(_03810_ ), .B(_00482_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06071_ ), .ZN(_00483_ ) );
OAI21_X2 _16221_ ( .A(_00483_ ), .B1(_03811_ ), .B2(\io_master_rdata [31] ), .ZN(_00484_ ) );
NOR2_X1 _16222_ ( .A1(_00484_ ), .A2(_06037_ ), .ZN(\myifu.data_in [31] ) );
CLKBUF_X2 _16223_ ( .A(_01951_ ), .Z(_00485_ ) );
CLKBUF_X2 _16224_ ( .A(_06070_ ), .Z(_00486_ ) );
CLKBUF_X2 _16225_ ( .A(_00486_ ), .Z(_00487_ ) );
OR3_X1 _16226_ ( .A1(_00485_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00487_ ), .ZN(_00488_ ) );
OAI211_X1 _16227_ ( .A(_03812_ ), .B(_00488_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06072_ ), .ZN(_00489_ ) );
BUF_X2 _16228_ ( .A(_03811_ ), .Z(_00490_ ) );
BUF_X2 _16229_ ( .A(_00490_ ), .Z(_00491_ ) );
OAI21_X1 _16230_ ( .A(_00489_ ), .B1(_00491_ ), .B2(\io_master_rdata [30] ), .ZN(_00492_ ) );
NOR2_X1 _16231_ ( .A1(_00492_ ), .A2(_06037_ ), .ZN(\myifu.data_in [30] ) );
MUX2_X1 _16232_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06072_ ), .Z(_00493_ ) );
AND3_X1 _16233_ ( .A1(_02065_ ), .A2(_02068_ ), .A3(_00493_ ), .ZN(_00494_ ) );
AOI21_X1 _16234_ ( .A(\io_master_rdata [21] ), .B1(_02065_ ), .B2(_02068_ ), .ZN(_00495_ ) );
NOR3_X1 _16235_ ( .A1(_00494_ ), .A2(_00495_ ), .A3(_01972_ ), .ZN(\myifu.data_in [21] ) );
OR3_X1 _16236_ ( .A1(_00485_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00496_ ) );
BUF_X4 _16237_ ( .A(_06071_ ), .Z(_00497_ ) );
OAI211_X1 _16238_ ( .A(_03812_ ), .B(_00496_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00497_ ), .ZN(_00498_ ) );
OAI21_X1 _16239_ ( .A(_00498_ ), .B1(\io_master_rdata [20] ), .B2(_03812_ ), .ZN(_00499_ ) );
NOR2_X1 _16240_ ( .A1(_00499_ ), .A2(_06037_ ), .ZN(\myifu.data_in [20] ) );
OR2_X1 _16241_ ( .A1(_03811_ ), .A2(\io_master_rdata [19] ), .ZN(_00500_ ) );
OR3_X1 _16242_ ( .A1(_00485_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00501_ ) );
OAI211_X1 _16243_ ( .A(_00490_ ), .B(_00501_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00497_ ), .ZN(_00502_ ) );
AND3_X1 _16244_ ( .A1(_00500_ ), .A2(_00502_ ), .A3(_02021_ ), .ZN(\myifu.data_in [19] ) );
OR2_X1 _16245_ ( .A1(_03813_ ), .A2(\io_master_rdata [18] ), .ZN(_00503_ ) );
CLKBUF_X2 _16246_ ( .A(_00487_ ), .Z(_00504_ ) );
OR3_X1 _16247_ ( .A1(_03816_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00505_ ) );
OAI211_X1 _16248_ ( .A(_03813_ ), .B(_00505_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06072_ ), .ZN(_00506_ ) );
AND3_X1 _16249_ ( .A1(_00503_ ), .A2(_00506_ ), .A3(_02022_ ), .ZN(\myifu.data_in [18] ) );
OR2_X1 _16250_ ( .A1(_03811_ ), .A2(\io_master_rdata [17] ), .ZN(_00507_ ) );
OR3_X1 _16251_ ( .A1(_00485_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00508_ ) );
OAI211_X1 _16252_ ( .A(_03811_ ), .B(_00508_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00497_ ), .ZN(_00509_ ) );
AND3_X1 _16253_ ( .A1(_00507_ ), .A2(_00509_ ), .A3(_02021_ ), .ZN(\myifu.data_in [17] ) );
OR2_X1 _16254_ ( .A1(_03813_ ), .A2(\io_master_rdata [16] ), .ZN(_00510_ ) );
OR3_X1 _16255_ ( .A1(_02020_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00487_ ), .ZN(_00511_ ) );
OAI211_X1 _16256_ ( .A(_03813_ ), .B(_00511_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06072_ ), .ZN(_00512_ ) );
AND3_X1 _16257_ ( .A1(_00510_ ), .A2(_00512_ ), .A3(_02021_ ), .ZN(\myifu.data_in [16] ) );
OR3_X1 _16258_ ( .A1(_01951_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06070_ ), .ZN(_00513_ ) );
OAI211_X1 _16259_ ( .A(_03811_ ), .B(_00513_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06071_ ), .ZN(_00514_ ) );
OAI21_X1 _16260_ ( .A(_00514_ ), .B1(_03811_ ), .B2(\io_master_rdata [15] ), .ZN(_00515_ ) );
NOR2_X1 _16261_ ( .A1(_00515_ ), .A2(_06036_ ), .ZN(\myifu.data_in [15] ) );
OR2_X1 _16262_ ( .A1(_00491_ ), .A2(\io_master_rdata [14] ), .ZN(_00516_ ) );
OR3_X1 _16263_ ( .A1(_02020_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00487_ ), .ZN(_00517_ ) );
OAI211_X1 _16264_ ( .A(_03813_ ), .B(_00517_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06072_ ), .ZN(_00518_ ) );
AND3_X1 _16265_ ( .A1(_00516_ ), .A2(_00518_ ), .A3(_02021_ ), .ZN(\myifu.data_in [14] ) );
BUF_X2 _16266_ ( .A(_00491_ ), .Z(_00519_ ) );
OR2_X1 _16267_ ( .A1(_00519_ ), .A2(\io_master_rdata [13] ), .ZN(_00520_ ) );
OR3_X1 _16268_ ( .A1(_03816_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00521_ ) );
OAI211_X1 _16269_ ( .A(_00519_ ), .B(_00521_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00522_ ) );
AND3_X1 _16270_ ( .A1(_00520_ ), .A2(_00522_ ), .A3(_02021_ ), .ZN(\myifu.data_in [13] ) );
OR2_X1 _16271_ ( .A1(_00491_ ), .A2(\io_master_rdata [12] ), .ZN(_00523_ ) );
OR3_X1 _16272_ ( .A1(_02020_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00487_ ), .ZN(_00524_ ) );
OAI211_X1 _16273_ ( .A(_03813_ ), .B(_00524_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06072_ ), .ZN(_00525_ ) );
AND3_X1 _16274_ ( .A1(_00523_ ), .A2(_00525_ ), .A3(_02021_ ), .ZN(\myifu.data_in [12] ) );
OR2_X1 _16275_ ( .A1(_00519_ ), .A2(\io_master_rdata [29] ), .ZN(_00526_ ) );
OR3_X1 _16276_ ( .A1(_03816_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00527_ ) );
OAI211_X1 _16277_ ( .A(_00519_ ), .B(_00527_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00528_ ) );
AND3_X1 _16278_ ( .A1(_00526_ ), .A2(_00528_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [29] ) );
OR2_X1 _16279_ ( .A1(_00491_ ), .A2(\io_master_rdata [11] ), .ZN(_00529_ ) );
OR3_X1 _16280_ ( .A1(_02020_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00487_ ), .ZN(_00530_ ) );
OAI211_X1 _16281_ ( .A(_00491_ ), .B(_00530_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06072_ ), .ZN(_00531_ ) );
AND3_X1 _16282_ ( .A1(_00529_ ), .A2(_00531_ ), .A3(_02022_ ), .ZN(\myifu.data_in [11] ) );
OR2_X1 _16283_ ( .A1(_00519_ ), .A2(\io_master_rdata [10] ), .ZN(_00532_ ) );
OR3_X1 _16284_ ( .A1(_02021_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00533_ ) );
OAI211_X1 _16285_ ( .A(_03814_ ), .B(_00533_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00534_ ) );
AND3_X1 _16286_ ( .A1(_00532_ ), .A2(_00534_ ), .A3(_02022_ ), .ZN(\myifu.data_in [10] ) );
OR2_X1 _16287_ ( .A1(_00491_ ), .A2(\io_master_rdata [9] ), .ZN(_00535_ ) );
OR3_X1 _16288_ ( .A1(_02020_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00487_ ), .ZN(_00536_ ) );
OAI211_X1 _16289_ ( .A(_00491_ ), .B(_00536_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06072_ ), .ZN(_00537_ ) );
AND3_X1 _16290_ ( .A1(_00535_ ), .A2(_00537_ ), .A3(_02022_ ), .ZN(\myifu.data_in [9] ) );
OR2_X1 _16291_ ( .A1(_00519_ ), .A2(\io_master_rdata [8] ), .ZN(_00538_ ) );
OR3_X1 _16292_ ( .A1(_03816_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00539_ ) );
OAI211_X1 _16293_ ( .A(_03814_ ), .B(_00539_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00540_ ) );
AND3_X1 _16294_ ( .A1(_00538_ ), .A2(_00540_ ), .A3(_02022_ ), .ZN(\myifu.data_in [8] ) );
OR3_X1 _16295_ ( .A1(_00485_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00541_ ) );
OAI211_X1 _16296_ ( .A(_00490_ ), .B(_00541_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00497_ ), .ZN(_00542_ ) );
OAI21_X1 _16297_ ( .A(_00542_ ), .B1(_00491_ ), .B2(\io_master_rdata [7] ), .ZN(_00543_ ) );
NOR2_X1 _16298_ ( .A1(_00543_ ), .A2(_06036_ ), .ZN(\myifu.data_in [7] ) );
OR3_X1 _16299_ ( .A1(_00485_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00544_ ) );
OAI211_X1 _16300_ ( .A(_00490_ ), .B(_00544_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00497_ ), .ZN(_00545_ ) );
OAI21_X1 _16301_ ( .A(_00545_ ), .B1(_03812_ ), .B2(\io_master_rdata [6] ), .ZN(_00546_ ) );
NOR2_X1 _16302_ ( .A1(_00546_ ), .A2(_06036_ ), .ZN(\myifu.data_in [6] ) );
OR3_X1 _16303_ ( .A1(_03816_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00547_ ) );
OAI211_X1 _16304_ ( .A(_00519_ ), .B(_00547_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00548_ ) );
OAI21_X1 _16305_ ( .A(_00548_ ), .B1(_03814_ ), .B2(\io_master_rdata [5] ), .ZN(_00549_ ) );
NOR2_X1 _16306_ ( .A1(_00549_ ), .A2(_06036_ ), .ZN(\myifu.data_in [5] ) );
OR3_X1 _16307_ ( .A1(_00485_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00550_ ) );
OAI211_X1 _16308_ ( .A(_00490_ ), .B(_00550_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00497_ ), .ZN(_00551_ ) );
OAI21_X1 _16309_ ( .A(_00551_ ), .B1(_03812_ ), .B2(\io_master_rdata [4] ), .ZN(_00552_ ) );
NOR2_X1 _16310_ ( .A1(_00552_ ), .A2(_06036_ ), .ZN(\myifu.data_in [4] ) );
OR3_X1 _16311_ ( .A1(_00485_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00553_ ) );
OAI211_X1 _16312_ ( .A(_03811_ ), .B(_00553_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00497_ ), .ZN(_00554_ ) );
OAI21_X1 _16313_ ( .A(_00554_ ), .B1(_00490_ ), .B2(\io_master_rdata [3] ), .ZN(_00555_ ) );
NOR2_X1 _16314_ ( .A1(_00555_ ), .A2(_01972_ ), .ZN(\myifu.data_in [3] ) );
OR3_X1 _16315_ ( .A1(_03816_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00556_ ) );
OAI211_X1 _16316_ ( .A(_00519_ ), .B(_00556_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00557_ ) );
OAI21_X1 _16317_ ( .A(_00557_ ), .B1(_03814_ ), .B2(\io_master_rdata [2] ), .ZN(_00558_ ) );
NOR2_X1 _16318_ ( .A1(_00558_ ), .A2(_01972_ ), .ZN(\myifu.data_in [2] ) );
OR3_X1 _16319_ ( .A1(_02020_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00487_ ), .ZN(_00559_ ) );
OAI211_X1 _16320_ ( .A(_03812_ ), .B(_00559_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06072_ ), .ZN(_00560_ ) );
OAI21_X1 _16321_ ( .A(_00560_ ), .B1(_00491_ ), .B2(\io_master_rdata [28] ), .ZN(_00561_ ) );
NOR2_X1 _16322_ ( .A1(_00561_ ), .A2(_06036_ ), .ZN(\myifu.data_in [28] ) );
OR3_X1 _16323_ ( .A1(_00485_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00562_ ) );
OAI211_X1 _16324_ ( .A(_03811_ ), .B(_00562_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06071_ ), .ZN(_00563_ ) );
OAI21_X1 _16325_ ( .A(_00563_ ), .B1(_00490_ ), .B2(\io_master_rdata [1] ), .ZN(_00564_ ) );
NOR2_X1 _16326_ ( .A1(_00564_ ), .A2(_01972_ ), .ZN(\myifu.data_in [1] ) );
OR3_X1 _16327_ ( .A1(_03816_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_00504_ ), .ZN(_00565_ ) );
OAI211_X1 _16328_ ( .A(_00519_ ), .B(_00565_ ), .C1(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .C2(\io_master_araddr [2] ), .ZN(_00566_ ) );
OAI21_X1 _16329_ ( .A(_00566_ ), .B1(_03814_ ), .B2(\io_master_rdata [0] ), .ZN(_00567_ ) );
NOR2_X1 _16330_ ( .A1(_00567_ ), .A2(_01972_ ), .ZN(\myifu.data_in [0] ) );
OR2_X1 _16331_ ( .A1(_00490_ ), .A2(\io_master_rdata [27] ), .ZN(_00568_ ) );
OR3_X1 _16332_ ( .A1(_02020_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00487_ ), .ZN(_00569_ ) );
OAI211_X1 _16333_ ( .A(_03812_ ), .B(_00569_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00497_ ), .ZN(_00570_ ) );
AND3_X1 _16334_ ( .A1(_00568_ ), .A2(_00570_ ), .A3(_02021_ ), .ZN(\myifu.data_in [27] ) );
OR2_X1 _16335_ ( .A1(_03813_ ), .A2(\io_master_rdata [26] ), .ZN(_00571_ ) );
OR3_X1 _16336_ ( .A1(_03816_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00572_ ) );
OAI211_X1 _16337_ ( .A(_00519_ ), .B(_00572_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00573_ ) );
AND3_X1 _16338_ ( .A1(_00571_ ), .A2(_00573_ ), .A3(_02022_ ), .ZN(\myifu.data_in [26] ) );
OR2_X1 _16339_ ( .A1(_00490_ ), .A2(\io_master_rdata [25] ), .ZN(_00574_ ) );
OR3_X1 _16340_ ( .A1(_02020_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00487_ ), .ZN(_00575_ ) );
OAI211_X1 _16341_ ( .A(_03812_ ), .B(_00575_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00497_ ), .ZN(_00576_ ) );
AND3_X1 _16342_ ( .A1(_00574_ ), .A2(_00576_ ), .A3(_02022_ ), .ZN(\myifu.data_in [25] ) );
OR2_X1 _16343_ ( .A1(_03813_ ), .A2(\io_master_rdata [24] ), .ZN(_00577_ ) );
OR3_X1 _16344_ ( .A1(_03816_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00578_ ) );
OAI211_X1 _16345_ ( .A(_03813_ ), .B(_00578_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00579_ ) );
AND3_X1 _16346_ ( .A1(_00577_ ), .A2(_00579_ ), .A3(_02021_ ), .ZN(\myifu.data_in [24] ) );
OR3_X1 _16347_ ( .A1(_01951_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06070_ ), .ZN(_00580_ ) );
OAI211_X1 _16348_ ( .A(_03810_ ), .B(_00580_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06071_ ), .ZN(_00581_ ) );
OAI21_X1 _16349_ ( .A(_00581_ ), .B1(_03810_ ), .B2(\io_master_rdata [23] ), .ZN(_00582_ ) );
NOR2_X1 _16350_ ( .A1(_00582_ ), .A2(_06036_ ), .ZN(\myifu.data_in [23] ) );
OR3_X1 _16351_ ( .A1(_00485_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00486_ ), .ZN(_00583_ ) );
OAI211_X1 _16352_ ( .A(_00490_ ), .B(_00583_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_00497_ ), .ZN(_00584_ ) );
OAI21_X1 _16353_ ( .A(_00584_ ), .B1(\io_master_rdata [22] ), .B2(_03812_ ), .ZN(_00585_ ) );
NOR2_X1 _16354_ ( .A1(_00585_ ), .A2(_06036_ ), .ZN(\myifu.data_in [22] ) );
INV_X1 _16355_ ( .A(_00242_ ), .ZN(_00586_ ) );
NAND2_X1 _16356_ ( .A1(_00586_ ), .A2(_02059_ ), .ZN(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16357_ ( .A1(_03745_ ), .A2(fanout_net_7 ), .ZN(_00587_ ) );
INV_X1 _16358_ ( .A(\myifu.myicache.valid_data_in ), .ZN(_00588_ ) );
OAI21_X1 _16359_ ( .A(_02059_ ), .B1(_00587_ ), .B2(_00588_ ), .ZN(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16360_ ( .A1(_03753_ ), .A2(fanout_net_11 ), .ZN(_00589_ ) );
OAI21_X1 _16361_ ( .A(_02059_ ), .B1(_00589_ ), .B2(_00588_ ), .ZN(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16362_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .ZN(_00590_ ) );
OAI21_X1 _16363_ ( .A(_02059_ ), .B1(_00590_ ), .B2(_00588_ ), .ZN(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ) );
NAND2_X1 _16364_ ( .A1(_03116_ ), .A2(_03122_ ), .ZN(_00591_ ) );
NAND2_X1 _16365_ ( .A1(_03260_ ), .A2(_03122_ ), .ZN(_00592_ ) );
AND2_X1 _16366_ ( .A1(_00591_ ), .A2(_00592_ ), .ZN(_00593_ ) );
AND2_X1 _16367_ ( .A1(_00593_ ), .A2(_03120_ ), .ZN(_00594_ ) );
INV_X1 _16368_ ( .A(_00594_ ), .ZN(_00595_ ) );
OAI21_X1 _16369_ ( .A(\IF_ID_inst [8] ), .B1(_00595_ ), .B2(_03370_ ), .ZN(_00596_ ) );
AND2_X1 _16370_ ( .A1(_03262_ ), .A2(_03371_ ), .ZN(_00597_ ) );
BUF_X2 _16371_ ( .A(_00597_ ), .Z(_00598_ ) );
AND2_X1 _16372_ ( .A1(_00598_ ), .A2(_03319_ ), .ZN(_00599_ ) );
AND4_X1 _16373_ ( .A1(_03056_ ), .A2(_03053_ ), .A3(_03094_ ), .A4(_03122_ ), .ZN(_00600_ ) );
NAND3_X1 _16374_ ( .A1(_00600_ ), .A2(_03107_ ), .A3(_03100_ ), .ZN(_00601_ ) );
NOR3_X1 _16375_ ( .A1(_00601_ ), .A2(_03110_ ), .A3(_03109_ ), .ZN(_00602_ ) );
NOR2_X1 _16376_ ( .A1(_00602_ ), .A2(_03072_ ), .ZN(_00603_ ) );
AND4_X1 _16377_ ( .A1(_03339_ ), .A2(_00603_ ), .A3(_03485_ ), .A4(_03242_ ), .ZN(_00604_ ) );
NAND3_X1 _16378_ ( .A1(_00599_ ), .A2(_03297_ ), .A3(_00604_ ), .ZN(_00605_ ) );
AND2_X1 _16379_ ( .A1(_00605_ ), .A2(_03485_ ), .ZN(_00606_ ) );
OAI221_X1 _16380_ ( .A(_00596_ ), .B1(_03302_ ), .B2(_03063_ ), .C1(_00606_ ), .C2(_03070_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ) );
AND2_X1 _16381_ ( .A1(_03163_ ), .A2(\IF_ID_inst [31] ), .ZN(_00607_ ) );
INV_X1 _16382_ ( .A(_00607_ ), .ZN(_00608_ ) );
OAI221_X1 _16383_ ( .A(_00608_ ), .B1(_00599_ ), .B2(_03064_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_03338_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ) );
NOR2_X1 _16384_ ( .A1(_03337_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_00609_ ) );
AOI21_X1 _16385_ ( .A(_03064_ ), .B1(_03262_ ), .B2(_03371_ ), .ZN(_00610_ ) );
NOR2_X1 _16386_ ( .A1(_00609_ ), .A2(_00610_ ), .ZN(_00611_ ) );
BUF_X4 _16387_ ( .A(_00611_ ), .Z(_00612_ ) );
BUF_X4 _16388_ ( .A(_00608_ ), .Z(_00613_ ) );
BUF_X4 _16389_ ( .A(_03319_ ), .Z(_00614_ ) );
OAI211_X1 _16390_ ( .A(_00612_ ), .B(_00613_ ), .C1(_03069_ ), .C2(_00614_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ) );
OAI211_X1 _16391_ ( .A(_00612_ ), .B(_00613_ ), .C1(_03070_ ), .C2(_00614_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ) );
OAI211_X1 _16392_ ( .A(_00612_ ), .B(_00613_ ), .C1(_03073_ ), .C2(_00614_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ) );
OAI21_X1 _16393_ ( .A(\IF_ID_inst [31] ), .B1(_00595_ ), .B2(_03370_ ), .ZN(_00615_ ) );
BUF_X2 _16394_ ( .A(_03338_ ), .Z(_00616_ ) );
OAI221_X1 _16395_ ( .A(_00615_ ), .B1(_03158_ ), .B2(_03168_ ), .C1(_00616_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ) );
OAI221_X1 _16396_ ( .A(_00615_ ), .B1(_03171_ ), .B2(_03168_ ), .C1(_00616_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ) );
OAI221_X1 _16397_ ( .A(_00615_ ), .B1(_03172_ ), .B2(_03168_ ), .C1(_00616_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ) );
OAI221_X1 _16398_ ( .A(_00615_ ), .B1(_03302_ ), .B2(_03168_ ), .C1(_00616_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ) );
OAI221_X1 _16399_ ( .A(_00615_ ), .B1(_03093_ ), .B2(_03168_ ), .C1(_00616_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ) );
OAI221_X1 _16400_ ( .A(_00615_ ), .B1(_03233_ ), .B2(_03168_ ), .C1(_00616_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ) );
OAI221_X1 _16401_ ( .A(_00615_ ), .B1(_03117_ ), .B2(_03168_ ), .C1(_00616_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ) );
OAI221_X1 _16402_ ( .A(_00615_ ), .B1(_03057_ ), .B2(_03168_ ), .C1(_00616_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ) );
OAI211_X1 _16403_ ( .A(_00612_ ), .B(_00613_ ), .C1(_03074_ ), .C2(_00614_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ) );
AOI21_X1 _16404_ ( .A(_03064_ ), .B1(_00593_ ), .B2(_03120_ ), .ZN(_00617_ ) );
AOI21_X1 _16405_ ( .A(_00617_ ), .B1(\IF_ID_inst [7] ), .B2(_03370_ ), .ZN(_00618_ ) );
OAI211_X1 _16406_ ( .A(_03534_ ), .B(_00618_ ), .C1(_00616_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ) );
INV_X1 _16407_ ( .A(_03549_ ), .ZN(_00619_ ) );
OAI221_X1 _16408_ ( .A(_00619_ ), .B1(_00598_ ), .B2(_03069_ ), .C1(_00616_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ) );
OAI221_X1 _16409_ ( .A(_03543_ ), .B1(_00598_ ), .B2(_03074_ ), .C1(_03338_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ) );
INV_X1 _16410_ ( .A(_03500_ ), .ZN(_00620_ ) );
OAI221_X1 _16411_ ( .A(_00620_ ), .B1(_00598_ ), .B2(_03075_ ), .C1(_03338_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ) );
OAI221_X1 _16412_ ( .A(_03504_ ), .B1(_00598_ ), .B2(_03076_ ), .C1(_03338_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ) );
INV_X1 _16413_ ( .A(_03495_ ), .ZN(_00621_ ) );
OAI221_X1 _16414_ ( .A(_00621_ ), .B1(_00598_ ), .B2(_03077_ ), .C1(_03338_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ) );
INV_X1 _16415_ ( .A(_03491_ ), .ZN(_00622_ ) );
OAI221_X1 _16416_ ( .A(_00622_ ), .B1(_00598_ ), .B2(_03078_ ), .C1(_03338_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ) );
OAI211_X1 _16417_ ( .A(_00612_ ), .B(_00613_ ), .C1(_03075_ ), .C2(_00614_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ) );
OAI211_X1 _16418_ ( .A(_00612_ ), .B(_00613_ ), .C1(_03076_ ), .C2(_00614_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ) );
OAI211_X1 _16419_ ( .A(_00612_ ), .B(_00613_ ), .C1(_03077_ ), .C2(_00614_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ) );
OAI211_X1 _16420_ ( .A(_00612_ ), .B(_00613_ ), .C1(_03078_ ), .C2(_00614_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ) );
OAI211_X1 _16421_ ( .A(_00612_ ), .B(_00613_ ), .C1(_03080_ ), .C2(_00614_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ) );
OAI211_X1 _16422_ ( .A(_00612_ ), .B(_00613_ ), .C1(_03081_ ), .C2(_00614_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ) );
OAI211_X1 _16423_ ( .A(_00611_ ), .B(_00608_ ), .C1(_03082_ ), .C2(_03319_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ) );
OAI21_X1 _16424_ ( .A(\IF_ID_inst [19] ), .B1(_03059_ ), .B2(_03061_ ), .ZN(_00623_ ) );
OAI221_X1 _16425_ ( .A(_00623_ ), .B1(_03096_ ), .B2(_00598_ ), .C1(_00606_ ), .C2(_03080_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ) );
OAI21_X1 _16426_ ( .A(\IF_ID_inst [18] ), .B1(_03059_ ), .B2(_03061_ ), .ZN(_00624_ ) );
OAI221_X1 _16427_ ( .A(_00624_ ), .B1(_03097_ ), .B2(_00598_ ), .C1(_00606_ ), .C2(_03081_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ) );
OAI21_X1 _16428_ ( .A(\IF_ID_inst [17] ), .B1(_03059_ ), .B2(_03061_ ), .ZN(_00625_ ) );
OAI221_X1 _16429_ ( .A(_00625_ ), .B1(_03098_ ), .B2(_00598_ ), .C1(_00606_ ), .C2(_03082_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ) );
OAI21_X1 _16430_ ( .A(\IF_ID_inst [15] ), .B1(_03059_ ), .B2(_03061_ ), .ZN(_00626_ ) );
OAI221_X1 _16431_ ( .A(_00626_ ), .B1(_03092_ ), .B2(_03262_ ), .C1(_00605_ ), .C2(_03073_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ) );
AND3_X1 _16432_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][8] ), .ZN(_00627_ ) );
AND3_X1 _16433_ ( .A1(_03744_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][8] ), .ZN(_00628_ ) );
AOI211_X1 _16434_ ( .A(_00627_ ), .B(_00628_ ), .C1(\myifu.myicache.data[0][8] ), .C2(_05999_ ), .ZN(_00629_ ) );
NAND2_X2 _16435_ ( .A1(_00588_ ), .A2(\IF_ID_pc [2] ), .ZN(_00630_ ) );
BUF_X2 _16436_ ( .A(_00630_ ), .Z(_00631_ ) );
NAND2_X2 _16437_ ( .A1(\myifu.tmp_offset [2] ), .A2(\myifu.myicache.valid_data_in ), .ZN(_00632_ ) );
BUF_X4 _16438_ ( .A(_00632_ ), .Z(_00633_ ) );
BUF_X4 _16439_ ( .A(_00633_ ), .Z(_00634_ ) );
NAND3_X1 _16440_ ( .A1(_03753_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][8] ), .ZN(_00635_ ) );
NAND4_X1 _16441_ ( .A1(_00629_ ), .A2(_00631_ ), .A3(_00634_ ), .A4(_00635_ ), .ZN(_00636_ ) );
NOR2_X1 _16442_ ( .A1(\myifu.state [1] ), .A2(\myifu.state [2] ), .ZN(_00637_ ) );
BUF_X2 _16443_ ( .A(_00637_ ), .Z(_00638_ ) );
BUF_X4 _16444_ ( .A(_00638_ ), .Z(_00639_ ) );
CLKBUF_X2 _16445_ ( .A(_03743_ ), .Z(_00640_ ) );
BUF_X4 _16446_ ( .A(_00640_ ), .Z(_00641_ ) );
NAND3_X1 _16447_ ( .A1(_00641_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][8] ), .ZN(_00642_ ) );
NAND3_X1 _16448_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][8] ), .ZN(_00643_ ) );
AND2_X1 _16449_ ( .A1(_00642_ ), .A2(_00643_ ), .ZN(_00644_ ) );
NAND2_X1 _16450_ ( .A1(_00630_ ), .A2(_00632_ ), .ZN(_00645_ ) );
BUF_X2 _16451_ ( .A(_00645_ ), .Z(_00646_ ) );
BUF_X4 _16452_ ( .A(_03752_ ), .Z(_00647_ ) );
BUF_X4 _16453_ ( .A(_00647_ ), .Z(_00648_ ) );
NAND3_X1 _16454_ ( .A1(_00648_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][8] ), .ZN(_00649_ ) );
BUF_X4 _16455_ ( .A(_03751_ ), .Z(_00650_ ) );
BUF_X4 _16456_ ( .A(_00650_ ), .Z(_00651_ ) );
NAND3_X1 _16457_ ( .A1(_03745_ ), .A2(_00651_ ), .A3(\myifu.myicache.data[1][8] ), .ZN(_00652_ ) );
NAND4_X1 _16458_ ( .A1(_00644_ ), .A2(_00646_ ), .A3(_00649_ ), .A4(_00652_ ), .ZN(_00653_ ) );
NAND3_X1 _16459_ ( .A1(_00636_ ), .A2(_00639_ ), .A3(_00653_ ), .ZN(_00654_ ) );
OR2_X1 _16460_ ( .A1(_03808_ ), .A2(_03822_ ), .ZN(_00655_ ) );
XOR2_X1 _16461_ ( .A(\IF_ID_pc [2] ), .B(\myifu.tmp_offset [2] ), .Z(_00656_ ) );
NAND2_X1 _16462_ ( .A1(_03470_ ), .A2(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ), .ZN(_00657_ ) );
NOR2_X1 _16463_ ( .A1(_00656_ ), .A2(_00657_ ), .ZN(_00658_ ) );
INV_X2 _16464_ ( .A(_00658_ ), .ZN(_00659_ ) );
NOR2_X1 _16465_ ( .A1(_00655_ ), .A2(_00659_ ), .ZN(_00660_ ) );
BUF_X4 _16466_ ( .A(_00660_ ), .Z(_00661_ ) );
OAI21_X1 _16467_ ( .A(\myifu.state [2] ), .B1(_00661_ ), .B2(_03467_ ), .ZN(_00662_ ) );
BUF_X4 _16468_ ( .A(_00659_ ), .Z(_00663_ ) );
NOR4_X1 _16469_ ( .A1(\myifu.data_in [8] ), .A2(_03809_ ), .A3(_03823_ ), .A4(_00663_ ), .ZN(_00664_ ) );
OAI21_X1 _16470_ ( .A(_00654_ ), .B1(_00662_ ), .B2(_00664_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ) );
AND3_X1 _16471_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][31] ), .ZN(_00665_ ) );
AND3_X1 _16472_ ( .A1(_03744_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][31] ), .ZN(_00666_ ) );
AOI211_X1 _16473_ ( .A(_00665_ ), .B(_00666_ ), .C1(\myifu.myicache.data[0][31] ), .C2(_05999_ ), .ZN(_00667_ ) );
NAND3_X1 _16474_ ( .A1(_03753_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][31] ), .ZN(_00668_ ) );
NAND4_X1 _16475_ ( .A1(_00667_ ), .A2(_00631_ ), .A3(_00634_ ), .A4(_00668_ ), .ZN(_00669_ ) );
NAND3_X1 _16476_ ( .A1(_00641_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][31] ), .ZN(_00670_ ) );
NAND3_X1 _16477_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][31] ), .ZN(_00671_ ) );
AND2_X1 _16478_ ( .A1(_00670_ ), .A2(_00671_ ), .ZN(_00672_ ) );
NAND3_X1 _16479_ ( .A1(_00648_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][31] ), .ZN(_00673_ ) );
NAND3_X1 _16480_ ( .A1(_03745_ ), .A2(_00651_ ), .A3(\myifu.myicache.data[1][31] ), .ZN(_00674_ ) );
NAND4_X1 _16481_ ( .A1(_00672_ ), .A2(_00646_ ), .A3(_00673_ ), .A4(_00674_ ), .ZN(_00675_ ) );
NAND3_X1 _16482_ ( .A1(_00669_ ), .A2(_00639_ ), .A3(_00675_ ), .ZN(_00676_ ) );
OAI21_X1 _16483_ ( .A(\myifu.state [2] ), .B1(_00661_ ), .B2(_03267_ ), .ZN(_00677_ ) );
BUF_X4 _16484_ ( .A(_00655_ ), .Z(_00678_ ) );
BUF_X4 _16485_ ( .A(_00678_ ), .Z(_00679_ ) );
BUF_X4 _16486_ ( .A(_00663_ ), .Z(_00680_ ) );
NOR3_X1 _16487_ ( .A1(_00679_ ), .A2(\myifu.data_in [31] ), .A3(_00680_ ), .ZN(_00681_ ) );
OAI21_X1 _16488_ ( .A(_00676_ ), .B1(_00677_ ), .B2(_00681_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ) );
AND3_X1 _16489_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][30] ), .ZN(_00682_ ) );
AND3_X1 _16490_ ( .A1(_03744_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][30] ), .ZN(_00683_ ) );
AOI211_X1 _16491_ ( .A(_00682_ ), .B(_00683_ ), .C1(\myifu.myicache.data[0][30] ), .C2(_05999_ ), .ZN(_00684_ ) );
NAND3_X1 _16492_ ( .A1(_03753_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][30] ), .ZN(_00685_ ) );
NAND4_X1 _16493_ ( .A1(_00684_ ), .A2(_00631_ ), .A3(_00634_ ), .A4(_00685_ ), .ZN(_00686_ ) );
NAND3_X1 _16494_ ( .A1(_00641_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][30] ), .ZN(_00687_ ) );
NAND3_X1 _16495_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][30] ), .ZN(_00688_ ) );
AND2_X1 _16496_ ( .A1(_00687_ ), .A2(_00688_ ), .ZN(_00689_ ) );
NAND3_X1 _16497_ ( .A1(_00648_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][30] ), .ZN(_00690_ ) );
NAND3_X1 _16498_ ( .A1(_03745_ ), .A2(_00651_ ), .A3(\myifu.myicache.data[1][30] ), .ZN(_00691_ ) );
NAND4_X1 _16499_ ( .A1(_00689_ ), .A2(_00646_ ), .A3(_00690_ ), .A4(_00691_ ), .ZN(_00692_ ) );
NAND3_X1 _16500_ ( .A1(_00686_ ), .A2(_00639_ ), .A3(_00692_ ), .ZN(_00693_ ) );
OAI21_X1 _16501_ ( .A(\myifu.state [2] ), .B1(_00661_ ), .B2(_03550_ ), .ZN(_00694_ ) );
NOR3_X1 _16502_ ( .A1(_00679_ ), .A2(\myifu.data_in [30] ), .A3(_00680_ ), .ZN(_00695_ ) );
OAI21_X1 _16503_ ( .A(_00693_ ), .B1(_00694_ ), .B2(_00695_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ) );
INV_X1 _16504_ ( .A(\myifu.state [2] ), .ZN(_00696_ ) );
BUF_X4 _16505_ ( .A(_00696_ ), .Z(_00697_ ) );
NOR3_X1 _16506_ ( .A1(_00678_ ), .A2(\myifu.data_in [21] ), .A3(_00663_ ), .ZN(_00698_ ) );
INV_X2 _16507_ ( .A(_00660_ ), .ZN(_00699_ ) );
BUF_X4 _16508_ ( .A(_00699_ ), .Z(_00700_ ) );
AOI211_X1 _16509_ ( .A(_00697_ ), .B(_00698_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00700_ ), .ZN(_00701_ ) );
AND3_X1 _16510_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][21] ), .ZN(_00702_ ) );
BUF_X4 _16511_ ( .A(_03742_ ), .Z(_00703_ ) );
AND3_X1 _16512_ ( .A1(_00703_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][21] ), .ZN(_00704_ ) );
BUF_X4 _16513_ ( .A(_05998_ ), .Z(_00705_ ) );
AOI211_X1 _16514_ ( .A(_00702_ ), .B(_00704_ ), .C1(\myifu.myicache.data[0][21] ), .C2(_00705_ ), .ZN(_00706_ ) );
BUF_X4 _16515_ ( .A(_00630_ ), .Z(_00707_ ) );
BUF_X4 _16516_ ( .A(_03752_ ), .Z(_00708_ ) );
NAND3_X1 _16517_ ( .A1(_00708_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][21] ), .ZN(_00709_ ) );
NAND4_X1 _16518_ ( .A1(_00706_ ), .A2(_00707_ ), .A3(_00633_ ), .A4(_00709_ ), .ZN(_00710_ ) );
NAND3_X1 _16519_ ( .A1(_00640_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][21] ), .ZN(_00711_ ) );
NAND3_X1 _16520_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][21] ), .ZN(_00712_ ) );
AND2_X1 _16521_ ( .A1(_00711_ ), .A2(_00712_ ), .ZN(_00713_ ) );
BUF_X4 _16522_ ( .A(_00645_ ), .Z(_00714_ ) );
NAND3_X1 _16523_ ( .A1(_00647_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][21] ), .ZN(_00715_ ) );
BUF_X4 _16524_ ( .A(_00703_ ), .Z(_00716_ ) );
NAND3_X1 _16525_ ( .A1(_00716_ ), .A2(_00650_ ), .A3(\myifu.myicache.data[1][21] ), .ZN(_00717_ ) );
NAND4_X1 _16526_ ( .A1(_00713_ ), .A2(_00714_ ), .A3(_00715_ ), .A4(_00717_ ), .ZN(_00718_ ) );
AND3_X1 _16527_ ( .A1(_00710_ ), .A2(_00638_ ), .A3(_00718_ ), .ZN(_00719_ ) );
OR2_X1 _16528_ ( .A1(_00701_ ), .A2(_00719_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ) );
AND3_X1 _16529_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][20] ), .ZN(_00720_ ) );
AND3_X1 _16530_ ( .A1(_03744_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][20] ), .ZN(_00721_ ) );
AOI211_X1 _16531_ ( .A(_00720_ ), .B(_00721_ ), .C1(\myifu.myicache.data[0][20] ), .C2(_05999_ ), .ZN(_00722_ ) );
NAND3_X1 _16532_ ( .A1(_03753_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][20] ), .ZN(_00723_ ) );
NAND4_X1 _16533_ ( .A1(_00722_ ), .A2(_00631_ ), .A3(_00634_ ), .A4(_00723_ ), .ZN(_00724_ ) );
NAND3_X1 _16534_ ( .A1(_00641_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][20] ), .ZN(_00725_ ) );
NAND3_X1 _16535_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][20] ), .ZN(_00726_ ) );
AND2_X1 _16536_ ( .A1(_00725_ ), .A2(_00726_ ), .ZN(_00727_ ) );
BUF_X4 _16537_ ( .A(_00714_ ), .Z(_00728_ ) );
NAND3_X1 _16538_ ( .A1(_00648_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][20] ), .ZN(_00729_ ) );
NAND3_X1 _16539_ ( .A1(_03745_ ), .A2(_00651_ ), .A3(\myifu.myicache.data[1][20] ), .ZN(_00730_ ) );
NAND4_X1 _16540_ ( .A1(_00727_ ), .A2(_00728_ ), .A3(_00729_ ), .A4(_00730_ ), .ZN(_00731_ ) );
NAND3_X1 _16541_ ( .A1(_00724_ ), .A2(_00639_ ), .A3(_00731_ ), .ZN(_00732_ ) );
OAI21_X1 _16542_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_00679_ ), .B2(_00680_ ), .ZN(_00733_ ) );
NAND2_X1 _16543_ ( .A1(_00733_ ), .A2(\myifu.state [2] ), .ZN(_00734_ ) );
NOR3_X1 _16544_ ( .A1(_00679_ ), .A2(\myifu.data_in [20] ), .A3(_00680_ ), .ZN(_00735_ ) );
OAI21_X1 _16545_ ( .A(_00732_ ), .B1(_00734_ ), .B2(_00735_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ) );
BUF_X4 _16546_ ( .A(_00659_ ), .Z(_00736_ ) );
NOR3_X1 _16547_ ( .A1(_00678_ ), .A2(\myifu.data_in [19] ), .A3(_00736_ ), .ZN(_00737_ ) );
AOI211_X1 _16548_ ( .A(_00697_ ), .B(_00737_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00700_ ), .ZN(_00738_ ) );
AND3_X1 _16549_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][19] ), .ZN(_00739_ ) );
CLKBUF_X2 _16550_ ( .A(_03742_ ), .Z(_00740_ ) );
AND3_X1 _16551_ ( .A1(_00740_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][19] ), .ZN(_00741_ ) );
AOI211_X1 _16552_ ( .A(_00739_ ), .B(_00741_ ), .C1(\myifu.myicache.data[0][19] ), .C2(_00705_ ), .ZN(_00742_ ) );
BUF_X4 _16553_ ( .A(_03752_ ), .Z(_00743_ ) );
NAND3_X1 _16554_ ( .A1(_00743_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][19] ), .ZN(_00744_ ) );
NAND4_X1 _16555_ ( .A1(_00742_ ), .A2(_00707_ ), .A3(_00633_ ), .A4(_00744_ ), .ZN(_00745_ ) );
BUF_X4 _16556_ ( .A(_03743_ ), .Z(_00746_ ) );
NAND3_X1 _16557_ ( .A1(_00746_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][19] ), .ZN(_00747_ ) );
NAND3_X1 _16558_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][19] ), .ZN(_00748_ ) );
AND2_X1 _16559_ ( .A1(_00747_ ), .A2(_00748_ ), .ZN(_00749_ ) );
NAND3_X1 _16560_ ( .A1(_00647_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][19] ), .ZN(_00750_ ) );
NAND3_X1 _16561_ ( .A1(_00716_ ), .A2(_00650_ ), .A3(\myifu.myicache.data[1][19] ), .ZN(_00751_ ) );
NAND4_X1 _16562_ ( .A1(_00749_ ), .A2(_00714_ ), .A3(_00750_ ), .A4(_00751_ ), .ZN(_00752_ ) );
AND3_X1 _16563_ ( .A1(_00745_ ), .A2(_00638_ ), .A3(_00752_ ), .ZN(_00753_ ) );
OR2_X1 _16564_ ( .A1(_00738_ ), .A2(_00753_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ) );
NOR4_X1 _16565_ ( .A1(\myifu.data_in [18] ), .A2(_03809_ ), .A3(_03823_ ), .A4(_00659_ ), .ZN(_00754_ ) );
AOI211_X1 _16566_ ( .A(_00697_ ), .B(_00754_ ), .C1(_00700_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00755_ ) );
AND3_X1 _16567_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][18] ), .ZN(_00756_ ) );
AND3_X1 _16568_ ( .A1(_00740_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][18] ), .ZN(_00757_ ) );
BUF_X4 _16569_ ( .A(_05998_ ), .Z(_00758_ ) );
AOI211_X1 _16570_ ( .A(_00756_ ), .B(_00757_ ), .C1(\myifu.myicache.data[0][18] ), .C2(_00758_ ), .ZN(_00759_ ) );
NAND3_X1 _16571_ ( .A1(_00743_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][18] ), .ZN(_00760_ ) );
NAND4_X1 _16572_ ( .A1(_00759_ ), .A2(_00707_ ), .A3(_00633_ ), .A4(_00760_ ), .ZN(_00761_ ) );
NAND3_X1 _16573_ ( .A1(_00746_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][18] ), .ZN(_00762_ ) );
NAND3_X1 _16574_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][18] ), .ZN(_00763_ ) );
AND2_X1 _16575_ ( .A1(_00762_ ), .A2(_00763_ ), .ZN(_00764_ ) );
BUF_X4 _16576_ ( .A(_03752_ ), .Z(_00765_ ) );
NAND3_X1 _16577_ ( .A1(_00765_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][18] ), .ZN(_00766_ ) );
NAND3_X1 _16578_ ( .A1(_00716_ ), .A2(_00650_ ), .A3(\myifu.myicache.data[1][18] ), .ZN(_00767_ ) );
NAND4_X1 _16579_ ( .A1(_00764_ ), .A2(_00714_ ), .A3(_00766_ ), .A4(_00767_ ), .ZN(_00768_ ) );
AND3_X1 _16580_ ( .A1(_00761_ ), .A2(_00638_ ), .A3(_00768_ ), .ZN(_00769_ ) );
OR2_X1 _16581_ ( .A1(_00755_ ), .A2(_00769_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ) );
NOR3_X1 _16582_ ( .A1(_00678_ ), .A2(\myifu.data_in [17] ), .A3(_00736_ ), .ZN(_00770_ ) );
AOI211_X1 _16583_ ( .A(_00697_ ), .B(_00770_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00700_ ), .ZN(_00771_ ) );
AND3_X1 _16584_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][17] ), .ZN(_00772_ ) );
AND3_X1 _16585_ ( .A1(_00740_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][17] ), .ZN(_00773_ ) );
AOI211_X1 _16586_ ( .A(_00772_ ), .B(_00773_ ), .C1(\myifu.myicache.data[0][17] ), .C2(_00758_ ), .ZN(_00774_ ) );
NAND3_X1 _16587_ ( .A1(_00743_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][17] ), .ZN(_00775_ ) );
NAND4_X1 _16588_ ( .A1(_00774_ ), .A2(_00707_ ), .A3(_00633_ ), .A4(_00775_ ), .ZN(_00776_ ) );
NAND3_X1 _16589_ ( .A1(_00746_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][17] ), .ZN(_00777_ ) );
NAND3_X1 _16590_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][17] ), .ZN(_00778_ ) );
AND2_X1 _16591_ ( .A1(_00777_ ), .A2(_00778_ ), .ZN(_00779_ ) );
NAND3_X1 _16592_ ( .A1(_00765_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][17] ), .ZN(_00780_ ) );
BUF_X4 _16593_ ( .A(_03751_ ), .Z(_00781_ ) );
NAND3_X1 _16594_ ( .A1(_00716_ ), .A2(_00781_ ), .A3(\myifu.myicache.data[1][17] ), .ZN(_00782_ ) );
NAND4_X1 _16595_ ( .A1(_00779_ ), .A2(_00714_ ), .A3(_00780_ ), .A4(_00782_ ), .ZN(_00783_ ) );
AND3_X1 _16596_ ( .A1(_00776_ ), .A2(_00638_ ), .A3(_00783_ ), .ZN(_00784_ ) );
OR2_X1 _16597_ ( .A1(_00771_ ), .A2(_00784_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ) );
NOR3_X1 _16598_ ( .A1(_00678_ ), .A2(\myifu.data_in [16] ), .A3(_00736_ ), .ZN(_00785_ ) );
AOI211_X1 _16599_ ( .A(_00697_ ), .B(_00785_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00700_ ), .ZN(_00786_ ) );
AND3_X1 _16600_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][16] ), .ZN(_00787_ ) );
AND3_X1 _16601_ ( .A1(_00740_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][16] ), .ZN(_00788_ ) );
AOI211_X1 _16602_ ( .A(_00787_ ), .B(_00788_ ), .C1(\myifu.myicache.data[0][16] ), .C2(_00758_ ), .ZN(_00789_ ) );
BUF_X4 _16603_ ( .A(_00632_ ), .Z(_00790_ ) );
NAND3_X1 _16604_ ( .A1(_00743_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][16] ), .ZN(_00791_ ) );
NAND4_X1 _16605_ ( .A1(_00789_ ), .A2(_00707_ ), .A3(_00790_ ), .A4(_00791_ ), .ZN(_00792_ ) );
NAND3_X1 _16606_ ( .A1(_00746_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][16] ), .ZN(_00793_ ) );
NAND3_X1 _16607_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][16] ), .ZN(_00794_ ) );
AND2_X1 _16608_ ( .A1(_00793_ ), .A2(_00794_ ), .ZN(_00795_ ) );
NAND3_X1 _16609_ ( .A1(_00765_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][16] ), .ZN(_00796_ ) );
NAND3_X1 _16610_ ( .A1(_00716_ ), .A2(_00781_ ), .A3(\myifu.myicache.data[1][16] ), .ZN(_00797_ ) );
NAND4_X1 _16611_ ( .A1(_00795_ ), .A2(_00714_ ), .A3(_00796_ ), .A4(_00797_ ), .ZN(_00798_ ) );
AND3_X1 _16612_ ( .A1(_00792_ ), .A2(_00638_ ), .A3(_00798_ ), .ZN(_00799_ ) );
OR2_X1 _16613_ ( .A1(_00786_ ), .A2(_00799_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ) );
NOR3_X1 _16614_ ( .A1(_00678_ ), .A2(\myifu.data_in [15] ), .A3(_00736_ ), .ZN(_00800_ ) );
AOI211_X1 _16615_ ( .A(_00697_ ), .B(_00800_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00700_ ), .ZN(_00801_ ) );
AND3_X1 _16616_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][15] ), .ZN(_00802_ ) );
AND3_X1 _16617_ ( .A1(_00740_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][15] ), .ZN(_00803_ ) );
AOI211_X1 _16618_ ( .A(_00802_ ), .B(_00803_ ), .C1(\myifu.myicache.data[0][15] ), .C2(_00758_ ), .ZN(_00804_ ) );
BUF_X4 _16619_ ( .A(_00630_ ), .Z(_00805_ ) );
NAND3_X1 _16620_ ( .A1(_00743_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][15] ), .ZN(_00806_ ) );
NAND4_X1 _16621_ ( .A1(_00804_ ), .A2(_00805_ ), .A3(_00790_ ), .A4(_00806_ ), .ZN(_00807_ ) );
CLKBUF_X2 _16622_ ( .A(_00637_ ), .Z(_00808_ ) );
NAND3_X1 _16623_ ( .A1(_00746_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][15] ), .ZN(_00809_ ) );
NAND3_X1 _16624_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][15] ), .ZN(_00810_ ) );
AND2_X1 _16625_ ( .A1(_00809_ ), .A2(_00810_ ), .ZN(_00811_ ) );
NAND3_X1 _16626_ ( .A1(_00765_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][15] ), .ZN(_00812_ ) );
BUF_X4 _16627_ ( .A(_00703_ ), .Z(_00813_ ) );
NAND3_X1 _16628_ ( .A1(_00813_ ), .A2(_00781_ ), .A3(\myifu.myicache.data[1][15] ), .ZN(_00814_ ) );
NAND4_X1 _16629_ ( .A1(_00811_ ), .A2(_00714_ ), .A3(_00812_ ), .A4(_00814_ ), .ZN(_00815_ ) );
AND3_X1 _16630_ ( .A1(_00807_ ), .A2(_00808_ ), .A3(_00815_ ), .ZN(_00816_ ) );
OR2_X1 _16631_ ( .A1(_00801_ ), .A2(_00816_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ) );
NOR3_X1 _16632_ ( .A1(_00678_ ), .A2(\myifu.data_in [14] ), .A3(_00736_ ), .ZN(_00817_ ) );
AOI211_X1 _16633_ ( .A(_00697_ ), .B(_00817_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00700_ ), .ZN(_00818_ ) );
AND3_X1 _16634_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][14] ), .ZN(_00819_ ) );
AND3_X1 _16635_ ( .A1(_00740_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][14] ), .ZN(_00820_ ) );
AOI211_X1 _16636_ ( .A(_00819_ ), .B(_00820_ ), .C1(\myifu.myicache.data[0][14] ), .C2(_00758_ ), .ZN(_00821_ ) );
NAND3_X1 _16637_ ( .A1(_00743_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][14] ), .ZN(_00822_ ) );
NAND4_X1 _16638_ ( .A1(_00821_ ), .A2(_00805_ ), .A3(_00790_ ), .A4(_00822_ ), .ZN(_00823_ ) );
NAND3_X1 _16639_ ( .A1(_00746_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][14] ), .ZN(_00824_ ) );
NAND3_X1 _16640_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][14] ), .ZN(_00825_ ) );
AND2_X1 _16641_ ( .A1(_00824_ ), .A2(_00825_ ), .ZN(_00826_ ) );
NAND3_X1 _16642_ ( .A1(_00765_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][14] ), .ZN(_00827_ ) );
NAND3_X1 _16643_ ( .A1(_00813_ ), .A2(_00781_ ), .A3(\myifu.myicache.data[1][14] ), .ZN(_00828_ ) );
NAND4_X1 _16644_ ( .A1(_00826_ ), .A2(_00714_ ), .A3(_00827_ ), .A4(_00828_ ), .ZN(_00829_ ) );
AND3_X1 _16645_ ( .A1(_00823_ ), .A2(_00808_ ), .A3(_00829_ ), .ZN(_00830_ ) );
OR2_X1 _16646_ ( .A1(_00818_ ), .A2(_00830_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ) );
BUF_X4 _16647_ ( .A(_00655_ ), .Z(_00831_ ) );
NOR3_X1 _16648_ ( .A1(_00831_ ), .A2(\myifu.data_in [13] ), .A3(_00736_ ), .ZN(_00832_ ) );
AOI211_X1 _16649_ ( .A(_00697_ ), .B(_00832_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00700_ ), .ZN(_00833_ ) );
AND3_X1 _16650_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][13] ), .ZN(_00834_ ) );
AND3_X1 _16651_ ( .A1(_00740_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][13] ), .ZN(_00835_ ) );
AOI211_X1 _16652_ ( .A(_00834_ ), .B(_00835_ ), .C1(\myifu.myicache.data[0][13] ), .C2(_00758_ ), .ZN(_00836_ ) );
NAND3_X1 _16653_ ( .A1(_00743_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][13] ), .ZN(_00837_ ) );
NAND4_X1 _16654_ ( .A1(_00836_ ), .A2(_00805_ ), .A3(_00790_ ), .A4(_00837_ ), .ZN(_00838_ ) );
NAND3_X1 _16655_ ( .A1(_00746_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][13] ), .ZN(_00839_ ) );
NAND3_X1 _16656_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][13] ), .ZN(_00840_ ) );
AND2_X1 _16657_ ( .A1(_00839_ ), .A2(_00840_ ), .ZN(_00841_ ) );
NAND3_X1 _16658_ ( .A1(_00765_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][13] ), .ZN(_00842_ ) );
NAND3_X1 _16659_ ( .A1(_00813_ ), .A2(_00781_ ), .A3(\myifu.myicache.data[1][13] ), .ZN(_00843_ ) );
NAND4_X1 _16660_ ( .A1(_00841_ ), .A2(_00714_ ), .A3(_00842_ ), .A4(_00843_ ), .ZN(_00844_ ) );
AND3_X1 _16661_ ( .A1(_00838_ ), .A2(_00808_ ), .A3(_00844_ ), .ZN(_00845_ ) );
OR2_X1 _16662_ ( .A1(_00833_ ), .A2(_00845_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ) );
NOR4_X1 _16663_ ( .A1(\myifu.data_in [12] ), .A2(_03808_ ), .A3(_03822_ ), .A4(_00659_ ), .ZN(_00846_ ) );
AOI211_X1 _16664_ ( .A(_00697_ ), .B(_00846_ ), .C1(_00700_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00847_ ) );
AND3_X1 _16665_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][12] ), .ZN(_00848_ ) );
AND3_X1 _16666_ ( .A1(_00740_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][12] ), .ZN(_00849_ ) );
AOI211_X1 _16667_ ( .A(_00848_ ), .B(_00849_ ), .C1(\myifu.myicache.data[0][12] ), .C2(_00758_ ), .ZN(_00850_ ) );
NAND3_X1 _16668_ ( .A1(_00743_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][12] ), .ZN(_00851_ ) );
NAND4_X1 _16669_ ( .A1(_00850_ ), .A2(_00805_ ), .A3(_00790_ ), .A4(_00851_ ), .ZN(_00852_ ) );
NAND3_X1 _16670_ ( .A1(_00746_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][12] ), .ZN(_00853_ ) );
NAND3_X1 _16671_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][12] ), .ZN(_00854_ ) );
AND2_X1 _16672_ ( .A1(_00853_ ), .A2(_00854_ ), .ZN(_00855_ ) );
BUF_X4 _16673_ ( .A(_00645_ ), .Z(_00856_ ) );
NAND3_X1 _16674_ ( .A1(_00765_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][12] ), .ZN(_00857_ ) );
NAND3_X1 _16675_ ( .A1(_00813_ ), .A2(_00781_ ), .A3(\myifu.myicache.data[1][12] ), .ZN(_00858_ ) );
NAND4_X1 _16676_ ( .A1(_00855_ ), .A2(_00856_ ), .A3(_00857_ ), .A4(_00858_ ), .ZN(_00859_ ) );
AND3_X1 _16677_ ( .A1(_00852_ ), .A2(_00808_ ), .A3(_00859_ ), .ZN(_00860_ ) );
OR2_X1 _16678_ ( .A1(_00847_ ), .A2(_00860_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ) );
AND3_X1 _16679_ ( .A1(fanout_net_13 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][29] ), .ZN(_00861_ ) );
AND3_X1 _16680_ ( .A1(_03744_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][29] ), .ZN(_00862_ ) );
AOI211_X1 _16681_ ( .A(_00861_ ), .B(_00862_ ), .C1(\myifu.myicache.data[0][29] ), .C2(_05999_ ), .ZN(_00863_ ) );
BUF_X4 _16682_ ( .A(_00708_ ), .Z(_00864_ ) );
NAND3_X1 _16683_ ( .A1(_00864_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][29] ), .ZN(_00865_ ) );
NAND4_X1 _16684_ ( .A1(_00863_ ), .A2(_00631_ ), .A3(_00634_ ), .A4(_00865_ ), .ZN(_00866_ ) );
NAND3_X1 _16685_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][29] ), .ZN(_00867_ ) );
NAND3_X1 _16686_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][29] ), .ZN(_00868_ ) );
AND2_X1 _16687_ ( .A1(_00867_ ), .A2(_00868_ ), .ZN(_00869_ ) );
NAND3_X1 _16688_ ( .A1(_00648_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][29] ), .ZN(_00870_ ) );
BUF_X4 _16689_ ( .A(_00716_ ), .Z(_00871_ ) );
NAND3_X1 _16690_ ( .A1(_00871_ ), .A2(_00651_ ), .A3(\myifu.myicache.data[1][29] ), .ZN(_00872_ ) );
NAND4_X1 _16691_ ( .A1(_00869_ ), .A2(_00728_ ), .A3(_00870_ ), .A4(_00872_ ), .ZN(_00873_ ) );
NAND3_X1 _16692_ ( .A1(_00866_ ), .A2(_00639_ ), .A3(_00873_ ), .ZN(_00874_ ) );
OAI21_X1 _16693_ ( .A(\myifu.state [2] ), .B1(_00661_ ), .B2(_03544_ ), .ZN(_00875_ ) );
NOR4_X1 _16694_ ( .A1(\myifu.data_in [29] ), .A2(_03809_ ), .A3(_03823_ ), .A4(_00663_ ), .ZN(_00876_ ) );
OAI21_X1 _16695_ ( .A(_00874_ ), .B1(_00875_ ), .B2(_00876_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ) );
AND3_X1 _16696_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][11] ), .ZN(_00877_ ) );
AND3_X1 _16697_ ( .A1(_03744_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][11] ), .ZN(_00878_ ) );
AOI211_X1 _16698_ ( .A(_00877_ ), .B(_00878_ ), .C1(\myifu.myicache.data[0][11] ), .C2(_05999_ ), .ZN(_00879_ ) );
NAND3_X1 _16699_ ( .A1(_00864_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][11] ), .ZN(_00880_ ) );
NAND4_X1 _16700_ ( .A1(_00879_ ), .A2(_00631_ ), .A3(_00634_ ), .A4(_00880_ ), .ZN(_00881_ ) );
NAND3_X1 _16701_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][11] ), .ZN(_00882_ ) );
NAND3_X1 _16702_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][11] ), .ZN(_00883_ ) );
AND2_X1 _16703_ ( .A1(_00882_ ), .A2(_00883_ ), .ZN(_00884_ ) );
NAND3_X1 _16704_ ( .A1(_00648_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][11] ), .ZN(_00885_ ) );
NAND3_X1 _16705_ ( .A1(_00871_ ), .A2(_00651_ ), .A3(\myifu.myicache.data[1][11] ), .ZN(_00886_ ) );
NAND4_X1 _16706_ ( .A1(_00884_ ), .A2(_00728_ ), .A3(_00885_ ), .A4(_00886_ ), .ZN(_00887_ ) );
NAND3_X1 _16707_ ( .A1(_00881_ ), .A2(_00639_ ), .A3(_00887_ ), .ZN(_00888_ ) );
OAI21_X1 _16708_ ( .A(\myifu.state [2] ), .B1(_00661_ ), .B2(_03483_ ), .ZN(_00889_ ) );
NOR4_X1 _16709_ ( .A1(\myifu.data_in [11] ), .A2(_03809_ ), .A3(_03823_ ), .A4(_00663_ ), .ZN(_00890_ ) );
OAI21_X1 _16710_ ( .A(_00888_ ), .B1(_00889_ ), .B2(_00890_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ) );
AND3_X1 _16711_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][10] ), .ZN(_00891_ ) );
AND3_X1 _16712_ ( .A1(_00640_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][10] ), .ZN(_00892_ ) );
AOI211_X1 _16713_ ( .A(_00891_ ), .B(_00892_ ), .C1(\myifu.myicache.data[0][10] ), .C2(_00705_ ), .ZN(_00893_ ) );
NAND3_X1 _16714_ ( .A1(_00864_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][10] ), .ZN(_00894_ ) );
NAND4_X1 _16715_ ( .A1(_00893_ ), .A2(_00631_ ), .A3(_00634_ ), .A4(_00894_ ), .ZN(_00895_ ) );
NAND3_X1 _16716_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][10] ), .ZN(_00896_ ) );
NAND3_X1 _16717_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][10] ), .ZN(_00897_ ) );
AND2_X1 _16718_ ( .A1(_00896_ ), .A2(_00897_ ), .ZN(_00898_ ) );
NAND3_X1 _16719_ ( .A1(_00648_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][10] ), .ZN(_00899_ ) );
NAND3_X1 _16720_ ( .A1(_00871_ ), .A2(_00708_ ), .A3(\myifu.myicache.data[1][10] ), .ZN(_00900_ ) );
NAND4_X1 _16721_ ( .A1(_00898_ ), .A2(_00728_ ), .A3(_00899_ ), .A4(_00900_ ), .ZN(_00901_ ) );
NAND3_X1 _16722_ ( .A1(_00895_ ), .A2(_00639_ ), .A3(_00901_ ), .ZN(_00902_ ) );
OAI21_X1 _16723_ ( .A(\myifu.state [2] ), .B1(_00661_ ), .B2(_03476_ ), .ZN(_00903_ ) );
NOR4_X1 _16724_ ( .A1(\myifu.data_in [10] ), .A2(_03809_ ), .A3(_03823_ ), .A4(_00663_ ), .ZN(_00904_ ) );
OAI21_X1 _16725_ ( .A(_00902_ ), .B1(_00903_ ), .B2(_00904_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ) );
AND3_X1 _16726_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][9] ), .ZN(_00905_ ) );
AND3_X1 _16727_ ( .A1(_00640_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][9] ), .ZN(_00906_ ) );
AOI211_X1 _16728_ ( .A(_00905_ ), .B(_00906_ ), .C1(\myifu.myicache.data[0][9] ), .C2(_00705_ ), .ZN(_00907_ ) );
NAND3_X1 _16729_ ( .A1(_00864_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][9] ), .ZN(_00908_ ) );
NAND4_X1 _16730_ ( .A1(_00907_ ), .A2(_00631_ ), .A3(_00634_ ), .A4(_00908_ ), .ZN(_00909_ ) );
NAND3_X1 _16731_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][9] ), .ZN(_00910_ ) );
NAND3_X1 _16732_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][9] ), .ZN(_00911_ ) );
AND2_X1 _16733_ ( .A1(_00910_ ), .A2(_00911_ ), .ZN(_00912_ ) );
NAND3_X1 _16734_ ( .A1(_00648_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][9] ), .ZN(_00913_ ) );
NAND3_X1 _16735_ ( .A1(_00871_ ), .A2(_00708_ ), .A3(\myifu.myicache.data[1][9] ), .ZN(_00914_ ) );
NAND4_X1 _16736_ ( .A1(_00912_ ), .A2(_00728_ ), .A3(_00913_ ), .A4(_00914_ ), .ZN(_00915_ ) );
NAND3_X1 _16737_ ( .A1(_00909_ ), .A2(_00639_ ), .A3(_00915_ ), .ZN(_00916_ ) );
OAI21_X1 _16738_ ( .A(\myifu.state [2] ), .B1(_00661_ ), .B2(_03463_ ), .ZN(_00917_ ) );
NOR3_X1 _16739_ ( .A1(_00679_ ), .A2(\myifu.data_in [9] ), .A3(_00680_ ), .ZN(_00918_ ) );
OAI21_X1 _16740_ ( .A(_00916_ ), .B1(_00917_ ), .B2(_00918_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ) );
BUF_X4 _16741_ ( .A(_00696_ ), .Z(_00919_ ) );
NOR3_X1 _16742_ ( .A1(_00831_ ), .A2(\myifu.data_in [7] ), .A3(_00736_ ), .ZN(_00920_ ) );
AOI211_X1 _16743_ ( .A(_00919_ ), .B(_00920_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00700_ ), .ZN(_00921_ ) );
AND3_X1 _16744_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][7] ), .ZN(_00922_ ) );
AND3_X1 _16745_ ( .A1(_00740_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][7] ), .ZN(_00923_ ) );
AOI211_X1 _16746_ ( .A(_00922_ ), .B(_00923_ ), .C1(\myifu.myicache.data[0][7] ), .C2(_00758_ ), .ZN(_00924_ ) );
NAND3_X1 _16747_ ( .A1(_00743_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][7] ), .ZN(_00925_ ) );
NAND4_X1 _16748_ ( .A1(_00924_ ), .A2(_00805_ ), .A3(_00790_ ), .A4(_00925_ ), .ZN(_00926_ ) );
NAND3_X1 _16749_ ( .A1(_00746_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][7] ), .ZN(_00927_ ) );
NAND3_X1 _16750_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][7] ), .ZN(_00928_ ) );
AND2_X1 _16751_ ( .A1(_00927_ ), .A2(_00928_ ), .ZN(_00929_ ) );
NAND3_X1 _16752_ ( .A1(_00765_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][7] ), .ZN(_00930_ ) );
NAND3_X1 _16753_ ( .A1(_00813_ ), .A2(_00781_ ), .A3(\myifu.myicache.data[1][7] ), .ZN(_00931_ ) );
NAND4_X1 _16754_ ( .A1(_00929_ ), .A2(_00856_ ), .A3(_00930_ ), .A4(_00931_ ), .ZN(_00932_ ) );
AND3_X1 _16755_ ( .A1(_00926_ ), .A2(_00808_ ), .A3(_00932_ ), .ZN(_00933_ ) );
OR2_X1 _16756_ ( .A1(_00921_ ), .A2(_00933_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ) );
AND3_X1 _16757_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][6] ), .ZN(_00934_ ) );
AND3_X1 _16758_ ( .A1(_00640_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][6] ), .ZN(_00935_ ) );
AOI211_X1 _16759_ ( .A(_00934_ ), .B(_00935_ ), .C1(\myifu.myicache.data[0][6] ), .C2(_00705_ ), .ZN(_00936_ ) );
NAND3_X1 _16760_ ( .A1(_00864_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][6] ), .ZN(_00937_ ) );
NAND4_X1 _16761_ ( .A1(_00936_ ), .A2(_00631_ ), .A3(_00634_ ), .A4(_00937_ ), .ZN(_00938_ ) );
NAND3_X1 _16762_ ( .A1(_00641_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][6] ), .ZN(_00939_ ) );
NAND3_X1 _16763_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][6] ), .ZN(_00940_ ) );
AND2_X1 _16764_ ( .A1(_00939_ ), .A2(_00940_ ), .ZN(_00941_ ) );
NAND3_X1 _16765_ ( .A1(_00648_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][6] ), .ZN(_00942_ ) );
NAND3_X1 _16766_ ( .A1(_00871_ ), .A2(_00708_ ), .A3(\myifu.myicache.data[1][6] ), .ZN(_00943_ ) );
NAND4_X1 _16767_ ( .A1(_00941_ ), .A2(_00728_ ), .A3(_00942_ ), .A4(_00943_ ), .ZN(_00944_ ) );
NAND3_X1 _16768_ ( .A1(_00938_ ), .A2(_00639_ ), .A3(_00944_ ), .ZN(_00945_ ) );
OAI21_X1 _16769_ ( .A(\myifu.state [2] ), .B1(_00661_ ), .B2(_03159_ ), .ZN(_00946_ ) );
NOR3_X1 _16770_ ( .A1(_00679_ ), .A2(\myifu.data_in [6] ), .A3(_00680_ ), .ZN(_00947_ ) );
OAI21_X1 _16771_ ( .A(_00945_ ), .B1(_00946_ ), .B2(_00947_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ) );
NOR3_X1 _16772_ ( .A1(_00831_ ), .A2(\myifu.data_in [5] ), .A3(_00736_ ), .ZN(_00948_ ) );
AOI211_X1 _16773_ ( .A(_00919_ ), .B(_00948_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00699_ ), .ZN(_00949_ ) );
AND3_X1 _16774_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][5] ), .ZN(_00950_ ) );
AND3_X1 _16775_ ( .A1(_00740_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][5] ), .ZN(_00951_ ) );
AOI211_X1 _16776_ ( .A(_00950_ ), .B(_00951_ ), .C1(\myifu.myicache.data[0][5] ), .C2(_00758_ ), .ZN(_00952_ ) );
NAND3_X1 _16777_ ( .A1(_00743_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][5] ), .ZN(_00953_ ) );
NAND4_X1 _16778_ ( .A1(_00952_ ), .A2(_00805_ ), .A3(_00790_ ), .A4(_00953_ ), .ZN(_00954_ ) );
NAND3_X1 _16779_ ( .A1(_00746_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][5] ), .ZN(_00955_ ) );
NAND3_X1 _16780_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][5] ), .ZN(_00956_ ) );
AND2_X1 _16781_ ( .A1(_00955_ ), .A2(_00956_ ), .ZN(_00957_ ) );
NAND3_X1 _16782_ ( .A1(_00765_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][5] ), .ZN(_00958_ ) );
NAND3_X1 _16783_ ( .A1(_00813_ ), .A2(_00781_ ), .A3(\myifu.myicache.data[1][5] ), .ZN(_00959_ ) );
NAND4_X1 _16784_ ( .A1(_00957_ ), .A2(_00856_ ), .A3(_00958_ ), .A4(_00959_ ), .ZN(_00960_ ) );
AND3_X1 _16785_ ( .A1(_00954_ ), .A2(_00808_ ), .A3(_00960_ ), .ZN(_00961_ ) );
OR2_X1 _16786_ ( .A1(_00949_ ), .A2(_00961_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ) );
NOR3_X1 _16787_ ( .A1(_00831_ ), .A2(\myifu.data_in [4] ), .A3(_00736_ ), .ZN(_00962_ ) );
AOI211_X1 _16788_ ( .A(_00919_ ), .B(_00962_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00699_ ), .ZN(_00963_ ) );
AND3_X1 _16789_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][4] ), .ZN(_00964_ ) );
AND3_X1 _16790_ ( .A1(_03743_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][4] ), .ZN(_00965_ ) );
AOI211_X1 _16791_ ( .A(_00964_ ), .B(_00965_ ), .C1(\myifu.myicache.data[0][4] ), .C2(_00758_ ), .ZN(_00966_ ) );
NAND3_X1 _16792_ ( .A1(_00647_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][4] ), .ZN(_00967_ ) );
NAND4_X1 _16793_ ( .A1(_00966_ ), .A2(_00805_ ), .A3(_00790_ ), .A4(_00967_ ), .ZN(_00968_ ) );
NAND3_X1 _16794_ ( .A1(_00703_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][4] ), .ZN(_00969_ ) );
NAND3_X1 _16795_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][4] ), .ZN(_00970_ ) );
AND2_X1 _16796_ ( .A1(_00969_ ), .A2(_00970_ ), .ZN(_00971_ ) );
NAND3_X1 _16797_ ( .A1(_00765_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][4] ), .ZN(_00972_ ) );
NAND3_X1 _16798_ ( .A1(_00813_ ), .A2(_00781_ ), .A3(\myifu.myicache.data[1][4] ), .ZN(_00973_ ) );
NAND4_X1 _16799_ ( .A1(_00971_ ), .A2(_00856_ ), .A3(_00972_ ), .A4(_00973_ ), .ZN(_00974_ ) );
AND3_X1 _16800_ ( .A1(_00968_ ), .A2(_00808_ ), .A3(_00974_ ), .ZN(_00975_ ) );
OR2_X1 _16801_ ( .A1(_00963_ ), .A2(_00975_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ) );
NOR3_X1 _16802_ ( .A1(_00831_ ), .A2(\myifu.data_in [3] ), .A3(_00736_ ), .ZN(_00976_ ) );
AOI211_X1 _16803_ ( .A(_00919_ ), .B(_00976_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00699_ ), .ZN(_00977_ ) );
AND3_X1 _16804_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][3] ), .ZN(_00978_ ) );
AND3_X1 _16805_ ( .A1(_03743_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][3] ), .ZN(_00979_ ) );
AOI211_X1 _16806_ ( .A(_00978_ ), .B(_00979_ ), .C1(\myifu.myicache.data[0][3] ), .C2(_05998_ ), .ZN(_00980_ ) );
NAND3_X1 _16807_ ( .A1(_00647_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][3] ), .ZN(_00981_ ) );
NAND4_X1 _16808_ ( .A1(_00980_ ), .A2(_00805_ ), .A3(_00790_ ), .A4(_00981_ ), .ZN(_00982_ ) );
NAND3_X1 _16809_ ( .A1(_00703_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][3] ), .ZN(_00983_ ) );
NAND3_X1 _16810_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][3] ), .ZN(_00984_ ) );
AND2_X1 _16811_ ( .A1(_00983_ ), .A2(_00984_ ), .ZN(_00985_ ) );
NAND3_X1 _16812_ ( .A1(_00650_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][3] ), .ZN(_00986_ ) );
NAND3_X1 _16813_ ( .A1(_00813_ ), .A2(_00781_ ), .A3(\myifu.myicache.data[1][3] ), .ZN(_00987_ ) );
NAND4_X1 _16814_ ( .A1(_00985_ ), .A2(_00856_ ), .A3(_00986_ ), .A4(_00987_ ), .ZN(_00988_ ) );
AND3_X1 _16815_ ( .A1(_00982_ ), .A2(_00808_ ), .A3(_00988_ ), .ZN(_00989_ ) );
OR2_X1 _16816_ ( .A1(_00977_ ), .A2(_00989_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ) );
NOR3_X1 _16817_ ( .A1(_00831_ ), .A2(\myifu.data_in [2] ), .A3(_00659_ ), .ZN(_00990_ ) );
AOI211_X1 _16818_ ( .A(_00919_ ), .B(_00990_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00699_ ), .ZN(_00991_ ) );
AND3_X1 _16819_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][2] ), .ZN(_00992_ ) );
AND3_X1 _16820_ ( .A1(_03743_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][2] ), .ZN(_00993_ ) );
AOI211_X1 _16821_ ( .A(_00992_ ), .B(_00993_ ), .C1(\myifu.myicache.data[0][2] ), .C2(_05998_ ), .ZN(_00994_ ) );
NAND3_X1 _16822_ ( .A1(_00647_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][2] ), .ZN(_00995_ ) );
NAND4_X1 _16823_ ( .A1(_00994_ ), .A2(_00805_ ), .A3(_00790_ ), .A4(_00995_ ), .ZN(_00996_ ) );
NAND3_X1 _16824_ ( .A1(_00703_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][2] ), .ZN(_00997_ ) );
NAND3_X1 _16825_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][2] ), .ZN(_00998_ ) );
AND2_X1 _16826_ ( .A1(_00997_ ), .A2(_00998_ ), .ZN(_00999_ ) );
NAND3_X1 _16827_ ( .A1(_00650_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][2] ), .ZN(_01000_ ) );
NAND3_X1 _16828_ ( .A1(_00813_ ), .A2(_03752_ ), .A3(\myifu.myicache.data[1][2] ), .ZN(_01001_ ) );
NAND4_X1 _16829_ ( .A1(_00999_ ), .A2(_00856_ ), .A3(_01000_ ), .A4(_01001_ ), .ZN(_01002_ ) );
AND3_X1 _16830_ ( .A1(_00996_ ), .A2(_00808_ ), .A3(_01002_ ), .ZN(_01003_ ) );
OR2_X1 _16831_ ( .A1(_00991_ ), .A2(_01003_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ) );
NOR3_X1 _16832_ ( .A1(_00831_ ), .A2(\myifu.data_in [1] ), .A3(_00659_ ), .ZN(_01004_ ) );
AOI211_X1 _16833_ ( .A(_00919_ ), .B(_01004_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00699_ ), .ZN(_01005_ ) );
AND3_X1 _16834_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][1] ), .ZN(_01006_ ) );
AND3_X1 _16835_ ( .A1(_03743_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][1] ), .ZN(_01007_ ) );
AOI211_X1 _16836_ ( .A(_01006_ ), .B(_01007_ ), .C1(\myifu.myicache.data[0][1] ), .C2(_05998_ ), .ZN(_01008_ ) );
NAND3_X1 _16837_ ( .A1(_00647_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][1] ), .ZN(_01009_ ) );
NAND4_X1 _16838_ ( .A1(_01008_ ), .A2(_00805_ ), .A3(_00632_ ), .A4(_01009_ ), .ZN(_01010_ ) );
NAND3_X1 _16839_ ( .A1(_00703_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][1] ), .ZN(_01011_ ) );
NAND3_X1 _16840_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][1] ), .ZN(_01012_ ) );
AND2_X1 _16841_ ( .A1(_01011_ ), .A2(_01012_ ), .ZN(_01013_ ) );
NAND3_X1 _16842_ ( .A1(_00650_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][1] ), .ZN(_01014_ ) );
NAND3_X1 _16843_ ( .A1(_00813_ ), .A2(_03752_ ), .A3(\myifu.myicache.data[1][1] ), .ZN(_01015_ ) );
NAND4_X1 _16844_ ( .A1(_01013_ ), .A2(_00856_ ), .A3(_01014_ ), .A4(_01015_ ), .ZN(_01016_ ) );
AND3_X1 _16845_ ( .A1(_01010_ ), .A2(_00808_ ), .A3(_01016_ ), .ZN(_01017_ ) );
OR2_X1 _16846_ ( .A1(_01005_ ), .A2(_01017_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ) );
AND3_X1 _16847_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][28] ), .ZN(_01018_ ) );
AND3_X1 _16848_ ( .A1(_00640_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][28] ), .ZN(_01019_ ) );
AOI211_X1 _16849_ ( .A(_01018_ ), .B(_01019_ ), .C1(\myifu.myicache.data[0][28] ), .C2(_00705_ ), .ZN(_01020_ ) );
NAND3_X1 _16850_ ( .A1(_00864_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][28] ), .ZN(_01021_ ) );
NAND4_X1 _16851_ ( .A1(_01020_ ), .A2(_00707_ ), .A3(_00633_ ), .A4(_01021_ ), .ZN(_01022_ ) );
NAND3_X1 _16852_ ( .A1(_00641_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][28] ), .ZN(_01023_ ) );
NAND3_X1 _16853_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][28] ), .ZN(_01024_ ) );
AND2_X1 _16854_ ( .A1(_01023_ ), .A2(_01024_ ), .ZN(_01025_ ) );
NAND3_X1 _16855_ ( .A1(_00648_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][28] ), .ZN(_01026_ ) );
NAND3_X1 _16856_ ( .A1(_00871_ ), .A2(_00708_ ), .A3(\myifu.myicache.data[1][28] ), .ZN(_01027_ ) );
NAND4_X1 _16857_ ( .A1(_01025_ ), .A2(_00728_ ), .A3(_01026_ ), .A4(_01027_ ), .ZN(_01028_ ) );
NAND3_X1 _16858_ ( .A1(_01022_ ), .A2(_00639_ ), .A3(_01028_ ), .ZN(_01029_ ) );
OAI21_X1 _16859_ ( .A(\myifu.state [2] ), .B1(_00661_ ), .B2(_03501_ ), .ZN(_01030_ ) );
NOR3_X1 _16860_ ( .A1(_00679_ ), .A2(\myifu.data_in [28] ), .A3(_00680_ ), .ZN(_01031_ ) );
OAI21_X1 _16861_ ( .A(_01029_ ), .B1(_01030_ ), .B2(_01031_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ) );
NOR3_X1 _16862_ ( .A1(_00831_ ), .A2(\myifu.data_in [0] ), .A3(_00659_ ), .ZN(_01032_ ) );
AOI211_X1 _16863_ ( .A(_00919_ ), .B(_01032_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00699_ ), .ZN(_01033_ ) );
AND3_X1 _16864_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][0] ), .ZN(_01034_ ) );
AND3_X1 _16865_ ( .A1(_03743_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][0] ), .ZN(_01035_ ) );
AOI211_X1 _16866_ ( .A(_01034_ ), .B(_01035_ ), .C1(\myifu.myicache.data[0][0] ), .C2(_05998_ ), .ZN(_01036_ ) );
NAND3_X1 _16867_ ( .A1(_00647_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][0] ), .ZN(_01037_ ) );
NAND4_X1 _16868_ ( .A1(_01036_ ), .A2(_00630_ ), .A3(_00632_ ), .A4(_01037_ ), .ZN(_01038_ ) );
NAND3_X1 _16869_ ( .A1(_00703_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][0] ), .ZN(_01039_ ) );
NAND3_X1 _16870_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][0] ), .ZN(_01040_ ) );
AND2_X1 _16871_ ( .A1(_01039_ ), .A2(_01040_ ), .ZN(_01041_ ) );
NAND3_X1 _16872_ ( .A1(_00650_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][0] ), .ZN(_01042_ ) );
NAND3_X1 _16873_ ( .A1(_03744_ ), .A2(_03752_ ), .A3(\myifu.myicache.data[1][0] ), .ZN(_01043_ ) );
NAND4_X1 _16874_ ( .A1(_01041_ ), .A2(_00856_ ), .A3(_01042_ ), .A4(_01043_ ), .ZN(_01044_ ) );
AND3_X1 _16875_ ( .A1(_01038_ ), .A2(_00637_ ), .A3(_01044_ ), .ZN(_01045_ ) );
OR2_X1 _16876_ ( .A1(_01033_ ), .A2(_01045_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ) );
NOR3_X1 _16877_ ( .A1(_00831_ ), .A2(\myifu.data_in [27] ), .A3(_00659_ ), .ZN(_01046_ ) );
AOI211_X1 _16878_ ( .A(_00919_ ), .B(_01046_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00699_ ), .ZN(_01047_ ) );
AND3_X1 _16879_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][27] ), .ZN(_01048_ ) );
AND3_X1 _16880_ ( .A1(_03743_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][27] ), .ZN(_01049_ ) );
AOI211_X1 _16881_ ( .A(_01048_ ), .B(_01049_ ), .C1(\myifu.myicache.data[0][27] ), .C2(_05998_ ), .ZN(_01050_ ) );
NAND3_X1 _16882_ ( .A1(_00647_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][27] ), .ZN(_01051_ ) );
NAND4_X1 _16883_ ( .A1(_01050_ ), .A2(_00630_ ), .A3(_00632_ ), .A4(_01051_ ), .ZN(_01052_ ) );
NAND3_X1 _16884_ ( .A1(_00703_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][27] ), .ZN(_01053_ ) );
NAND3_X1 _16885_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][27] ), .ZN(_01054_ ) );
AND2_X1 _16886_ ( .A1(_01053_ ), .A2(_01054_ ), .ZN(_01055_ ) );
NAND3_X1 _16887_ ( .A1(_00650_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][27] ), .ZN(_01056_ ) );
NAND3_X1 _16888_ ( .A1(_03744_ ), .A2(_03752_ ), .A3(\myifu.myicache.data[1][27] ), .ZN(_01057_ ) );
NAND4_X1 _16889_ ( .A1(_01055_ ), .A2(_00856_ ), .A3(_01056_ ), .A4(_01057_ ), .ZN(_01058_ ) );
AND3_X1 _16890_ ( .A1(_01052_ ), .A2(_00637_ ), .A3(_01058_ ), .ZN(_01059_ ) );
OR2_X1 _16891_ ( .A1(_01047_ ), .A2(_01059_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ) );
AND3_X1 _16892_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][26] ), .ZN(_01060_ ) );
AND3_X1 _16893_ ( .A1(_00640_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][26] ), .ZN(_01061_ ) );
AOI211_X1 _16894_ ( .A(_01060_ ), .B(_01061_ ), .C1(\myifu.myicache.data[0][26] ), .C2(_00705_ ), .ZN(_01062_ ) );
NAND3_X1 _16895_ ( .A1(_00864_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][26] ), .ZN(_01063_ ) );
NAND4_X1 _16896_ ( .A1(_01062_ ), .A2(_00707_ ), .A3(_00633_ ), .A4(_01063_ ), .ZN(_01064_ ) );
NAND3_X1 _16897_ ( .A1(_00716_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][26] ), .ZN(_01065_ ) );
NAND3_X1 _16898_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][26] ), .ZN(_01066_ ) );
AND2_X1 _16899_ ( .A1(_01065_ ), .A2(_01066_ ), .ZN(_01067_ ) );
NAND3_X1 _16900_ ( .A1(_00651_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][26] ), .ZN(_01068_ ) );
NAND3_X1 _16901_ ( .A1(_00871_ ), .A2(_00708_ ), .A3(\myifu.myicache.data[1][26] ), .ZN(_01069_ ) );
NAND4_X1 _16902_ ( .A1(_01067_ ), .A2(_00728_ ), .A3(_01068_ ), .A4(_01069_ ), .ZN(_01070_ ) );
NAND3_X1 _16903_ ( .A1(_01064_ ), .A2(_00638_ ), .A3(_01070_ ), .ZN(_01071_ ) );
OAI21_X1 _16904_ ( .A(\myifu.state [2] ), .B1(_00661_ ), .B2(_03496_ ), .ZN(_01072_ ) );
NOR3_X1 _16905_ ( .A1(_00679_ ), .A2(\myifu.data_in [26] ), .A3(_00680_ ), .ZN(_01073_ ) );
OAI21_X1 _16906_ ( .A(_01071_ ), .B1(_01072_ ), .B2(_01073_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ) );
AND3_X1 _16907_ ( .A1(\IF_ID_pc [4] ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][25] ), .ZN(_01074_ ) );
AND3_X1 _16908_ ( .A1(_00640_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][25] ), .ZN(_01075_ ) );
AOI211_X1 _16909_ ( .A(_01074_ ), .B(_01075_ ), .C1(\myifu.myicache.data[0][25] ), .C2(_00705_ ), .ZN(_01076_ ) );
NAND3_X1 _16910_ ( .A1(_00864_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][25] ), .ZN(_01077_ ) );
NAND4_X1 _16911_ ( .A1(_01076_ ), .A2(_00707_ ), .A3(_00633_ ), .A4(_01077_ ), .ZN(_01078_ ) );
NAND3_X1 _16912_ ( .A1(_00716_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][25] ), .ZN(_01079_ ) );
NAND3_X1 _16913_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][25] ), .ZN(_01080_ ) );
AND2_X1 _16914_ ( .A1(_01079_ ), .A2(_01080_ ), .ZN(_01081_ ) );
NAND3_X1 _16915_ ( .A1(_00651_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][25] ), .ZN(_01082_ ) );
NAND3_X1 _16916_ ( .A1(_00871_ ), .A2(_00708_ ), .A3(\myifu.myicache.data[1][25] ), .ZN(_01083_ ) );
NAND4_X1 _16917_ ( .A1(_01081_ ), .A2(_00728_ ), .A3(_01082_ ), .A4(_01083_ ), .ZN(_01084_ ) );
NAND3_X1 _16918_ ( .A1(_01078_ ), .A2(_00638_ ), .A3(_01084_ ), .ZN(_01085_ ) );
OAI21_X1 _16919_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .B1(_00678_ ), .B2(_00663_ ), .ZN(_01086_ ) );
NAND2_X1 _16920_ ( .A1(_01086_ ), .A2(\myifu.state [2] ), .ZN(_01087_ ) );
NOR4_X1 _16921_ ( .A1(\myifu.data_in [25] ), .A2(_03809_ ), .A3(_03823_ ), .A4(_00663_ ), .ZN(_01088_ ) );
OAI21_X1 _16922_ ( .A(_01085_ ), .B1(_01087_ ), .B2(_01088_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ) );
NOR3_X1 _16923_ ( .A1(_00831_ ), .A2(\myifu.data_in [24] ), .A3(_00659_ ), .ZN(_01089_ ) );
AOI211_X1 _16924_ ( .A(_00919_ ), .B(_01089_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00699_ ), .ZN(_01090_ ) );
AND3_X1 _16925_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][24] ), .ZN(_01091_ ) );
AND3_X1 _16926_ ( .A1(_03743_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][24] ), .ZN(_01092_ ) );
AOI211_X1 _16927_ ( .A(_01091_ ), .B(_01092_ ), .C1(\myifu.myicache.data[0][24] ), .C2(_05998_ ), .ZN(_01093_ ) );
NAND3_X1 _16928_ ( .A1(_00647_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][24] ), .ZN(_01094_ ) );
NAND4_X1 _16929_ ( .A1(_01093_ ), .A2(_00630_ ), .A3(_00632_ ), .A4(_01094_ ), .ZN(_01095_ ) );
NAND3_X1 _16930_ ( .A1(_00703_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][24] ), .ZN(_01096_ ) );
NAND3_X1 _16931_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][24] ), .ZN(_01097_ ) );
AND2_X1 _16932_ ( .A1(_01096_ ), .A2(_01097_ ), .ZN(_01098_ ) );
NAND3_X1 _16933_ ( .A1(_00650_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][24] ), .ZN(_01099_ ) );
NAND3_X1 _16934_ ( .A1(_03744_ ), .A2(_03752_ ), .A3(\myifu.myicache.data[1][24] ), .ZN(_01100_ ) );
NAND4_X1 _16935_ ( .A1(_01098_ ), .A2(_00856_ ), .A3(_01099_ ), .A4(_01100_ ), .ZN(_01101_ ) );
AND3_X1 _16936_ ( .A1(_01095_ ), .A2(_00637_ ), .A3(_01101_ ), .ZN(_01102_ ) );
OR2_X1 _16937_ ( .A1(_01090_ ), .A2(_01102_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ) );
AND3_X1 _16938_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][23] ), .ZN(_01103_ ) );
AND3_X1 _16939_ ( .A1(_00640_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][23] ), .ZN(_01104_ ) );
AOI211_X1 _16940_ ( .A(_01103_ ), .B(_01104_ ), .C1(\myifu.myicache.data[0][23] ), .C2(_00705_ ), .ZN(_01105_ ) );
NAND3_X1 _16941_ ( .A1(_00864_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][23] ), .ZN(_01106_ ) );
NAND4_X1 _16942_ ( .A1(_01105_ ), .A2(_00707_ ), .A3(_00633_ ), .A4(_01106_ ), .ZN(_01107_ ) );
NAND3_X1 _16943_ ( .A1(_00716_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][23] ), .ZN(_01108_ ) );
NAND3_X1 _16944_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][23] ), .ZN(_01109_ ) );
AND2_X1 _16945_ ( .A1(_01108_ ), .A2(_01109_ ), .ZN(_01110_ ) );
NAND3_X1 _16946_ ( .A1(_00651_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][23] ), .ZN(_01111_ ) );
NAND3_X1 _16947_ ( .A1(_00871_ ), .A2(_00708_ ), .A3(\myifu.myicache.data[1][23] ), .ZN(_01112_ ) );
NAND4_X1 _16948_ ( .A1(_01110_ ), .A2(_00728_ ), .A3(_01111_ ), .A4(_01112_ ), .ZN(_01113_ ) );
NAND3_X1 _16949_ ( .A1(_01107_ ), .A2(_00638_ ), .A3(_01113_ ), .ZN(_01114_ ) );
OAI21_X1 _16950_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B1(_00678_ ), .B2(_00663_ ), .ZN(_01115_ ) );
NAND2_X1 _16951_ ( .A1(_01115_ ), .A2(\myifu.state [2] ), .ZN(_01116_ ) );
NOR3_X1 _16952_ ( .A1(_00679_ ), .A2(\myifu.data_in [23] ), .A3(_00680_ ), .ZN(_01117_ ) );
OAI21_X1 _16953_ ( .A(_01114_ ), .B1(_01116_ ), .B2(_01117_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ) );
AND3_X1 _16954_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][22] ), .ZN(_01118_ ) );
AND3_X1 _16955_ ( .A1(_00640_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][22] ), .ZN(_01119_ ) );
AOI211_X1 _16956_ ( .A(_01118_ ), .B(_01119_ ), .C1(\myifu.myicache.data[0][22] ), .C2(_00705_ ), .ZN(_01120_ ) );
NAND3_X1 _16957_ ( .A1(_00864_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][22] ), .ZN(_01121_ ) );
NAND4_X1 _16958_ ( .A1(_01120_ ), .A2(_00707_ ), .A3(_00633_ ), .A4(_01121_ ), .ZN(_01122_ ) );
NAND3_X1 _16959_ ( .A1(_00716_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][22] ), .ZN(_01123_ ) );
NAND3_X1 _16960_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][22] ), .ZN(_01124_ ) );
AND2_X1 _16961_ ( .A1(_01123_ ), .A2(_01124_ ), .ZN(_01125_ ) );
NAND3_X1 _16962_ ( .A1(_00651_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][22] ), .ZN(_01126_ ) );
NAND3_X1 _16963_ ( .A1(_00871_ ), .A2(_00708_ ), .A3(\myifu.myicache.data[1][22] ), .ZN(_01127_ ) );
NAND4_X1 _16964_ ( .A1(_01125_ ), .A2(_00714_ ), .A3(_01126_ ), .A4(_01127_ ), .ZN(_01128_ ) );
NAND3_X1 _16965_ ( .A1(_01122_ ), .A2(_00638_ ), .A3(_01128_ ), .ZN(_01129_ ) );
OAI21_X1 _16966_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .B1(_00678_ ), .B2(_00663_ ), .ZN(_01130_ ) );
NAND2_X1 _16967_ ( .A1(_01130_ ), .A2(\myifu.state [2] ), .ZN(_01131_ ) );
NOR3_X1 _16968_ ( .A1(_00679_ ), .A2(\myifu.data_in [22] ), .A3(_00680_ ), .ZN(_01132_ ) );
OAI21_X1 _16969_ ( .A(_01129_ ), .B1(_01131_ ), .B2(_01132_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ) );
AOI211_X1 _16970_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .B(_03218_ ), .C1(_03627_ ), .C2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_E ) );
OR4_X1 _16971_ ( .A1(_01795_ ), .A2(_01827_ ), .A3(_01847_ ), .A4(_01859_ ), .ZN(_01133_ ) );
NAND2_X1 _16972_ ( .A1(_01906_ ), .A2(_01945_ ), .ZN(_01134_ ) );
INV_X1 _16973_ ( .A(\myifu.state [0] ), .ZN(_01135_ ) );
NOR4_X1 _16974_ ( .A1(_01133_ ), .A2(_01134_ ), .A3(\myidu.stall_quest_fencei ), .A4(_01135_ ), .ZN(_01136_ ) );
NOR4_X1 _16975_ ( .A1(_03809_ ), .A2(_00919_ ), .A3(_03815_ ), .A4(_03823_ ), .ZN(_01137_ ) );
AOI211_X1 _16976_ ( .A(_01136_ ), .B(_01137_ ), .C1(_03365_ ), .C2(\myifu.state [1] ), .ZN(_01138_ ) );
NOR2_X1 _16977_ ( .A1(_01138_ ), .A2(reset ), .ZN(\myifu.state_$_DFF_P__Q_1_D ) );
NOR2_X1 _16978_ ( .A1(_05989_ ), .A2(_06036_ ), .ZN(_01139_ ) );
NOR2_X1 _16979_ ( .A1(_01133_ ), .A2(_01134_ ), .ZN(_01140_ ) );
NOR4_X1 _16980_ ( .A1(_01139_ ), .A2(\myidu.stall_quest_fencei ), .A3(_01135_ ), .A4(_01140_ ), .ZN(_01141_ ) );
AND2_X1 _16981_ ( .A1(\myidu.stall_quest_fencei ), .A2(\myifu.state [0] ), .ZN(_01142_ ) );
OR4_X1 _16982_ ( .A1(reset ), .A2(_01141_ ), .A3(\myifu.pc_$_SDFFE_PP1P__Q_E ), .A4(_01142_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D ) );
NAND3_X1 _16983_ ( .A1(_03824_ ), .A2(_01618_ ), .A3(\myifu.state [2] ), .ZN(_01143_ ) );
NAND2_X1 _16984_ ( .A1(_01139_ ), .A2(_02071_ ), .ZN(_01144_ ) );
NAND2_X1 _16985_ ( .A1(_01143_ ), .A2(_01144_ ), .ZN(\myifu.state_$_DFF_P__Q_D ) );
NOR3_X1 _16986_ ( .A1(_03809_ ), .A2(_00697_ ), .A3(_03823_ ), .ZN(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ) );
INV_X1 _16987_ ( .A(\myifu.wen_$_ANDNOT__A_Y ), .ZN(_01145_ ) );
NOR3_X1 _16988_ ( .A1(_01145_ ), .A2(_00589_ ), .A3(_00646_ ), .ZN(\myifu.myicache.data[4]_$_DFFE_PP__Q_E ) );
NOR3_X1 _16989_ ( .A1(_01145_ ), .A2(_00590_ ), .A3(_00646_ ), .ZN(\myifu.myicache.data[6]_$_DFFE_PP__Q_E ) );
AND4_X1 _16990_ ( .A1(\IF_ID_pc [4] ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00646_ ), .ZN(\myifu.myicache.data[7]_$_DFFE_PP__Q_E ) );
AND4_X1 _16991_ ( .A1(\IF_ID_pc [4] ), .A2(_05997_ ), .A3(_03753_ ), .A4(_00646_ ), .ZN(\myifu.myicache.data[5]_$_DFFE_PP__Q_E ) );
NOR3_X1 _16992_ ( .A1(_01145_ ), .A2(_00587_ ), .A3(_00646_ ), .ZN(\myifu.myicache.data[2]_$_DFFE_PP__Q_E ) );
AND4_X1 _16993_ ( .A1(_03745_ ), .A2(_05997_ ), .A3(\IF_ID_pc [3] ), .A4(_00646_ ), .ZN(\myifu.myicache.data[3]_$_DFFE_PP__Q_E ) );
AND3_X1 _16994_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_05999_ ), .A3(_00646_ ), .ZN(\myifu.myicache.data[1]_$_DFFE_PP__Q_E ) );
AND4_X1 _16995_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_05999_ ), .A3(_00631_ ), .A4(_00634_ ), .ZN(\myifu.myicache.data[0]_$_DFFE_PP__Q_E ) );
AND3_X1 _16996_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_03745_ ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.myicache.tag[1]_$_DFFE_PP__Q_E ) );
AND3_X1 _16997_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(_03753_ ), .ZN(\myifu.myicache.tag[2]_$_DFFE_PP__Q_E ) );
AND3_X1 _16998_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.myicache.tag[3]_$_DFFE_PP__Q_E ) );
AND3_X1 _16999_ ( .A1(_02059_ ), .A2(_05999_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(\myifu.myicache.tag[0]_$_DFFE_PP__Q_E ) );
NOR2_X1 _17000_ ( .A1(_01139_ ), .A2(_01135_ ), .ZN(_01146_ ) );
AND2_X1 _17001_ ( .A1(_00481_ ), .A2(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01147_ ) );
NOR2_X1 _17002_ ( .A1(_01146_ ), .A2(_01147_ ), .ZN(_01148_ ) );
NOR2_X1 _17003_ ( .A1(_01946_ ), .A2(_01135_ ), .ZN(_01149_ ) );
INV_X1 _17004_ ( .A(_01149_ ), .ZN(_01150_ ) );
NOR3_X1 _17005_ ( .A1(_03809_ ), .A2(_03815_ ), .A3(_03823_ ), .ZN(_01151_ ) );
OAI211_X1 _17006_ ( .A(_01148_ ), .B(_01150_ ), .C1(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .C2(_01151_ ), .ZN(_01152_ ) );
NOR4_X1 _17007_ ( .A1(_01152_ ), .A2(_03219_ ), .A3(_00479_ ), .A4(_01142_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _17008_ ( .A1(_03618_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03220_ ), .ZN(\myidu.typ_$_SDFFE_PP0P__Q_E ) );
AND4_X1 _17009_ ( .A1(_03139_ ), .A2(_03141_ ), .A3(_03143_ ), .A4(_03144_ ), .ZN(_01153_ ) );
AND2_X1 _17010_ ( .A1(_03151_ ), .A2(_01153_ ), .ZN(_01154_ ) );
INV_X1 _17011_ ( .A(_01154_ ), .ZN(_01155_ ) );
AOI211_X1 _17012_ ( .A(_03365_ ), .B(_00464_ ), .C1(_03063_ ), .C2(_01155_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ) );
OR4_X1 _17013_ ( .A1(reset ), .A2(_01147_ ), .A3(_00479_ ), .A4(_01142_ ), .ZN(_01156_ ) );
AOI211_X1 _17014_ ( .A(_03219_ ), .B(_01156_ ), .C1(_01946_ ), .C2(\myifu.state [0] ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
INV_X2 _17015_ ( .A(\mylsu.state [3] ), .ZN(_01157_ ) );
MUX2_X1 _17016_ ( .A(_01157_ ), .B(_01986_ ), .S(\mylsu.state [0] ), .Z(_01158_ ) );
AOI21_X1 _17017_ ( .A(_01158_ ), .B1(_06092_ ), .B2(\mylsu.state [3] ), .ZN(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ) );
AOI211_X1 _17018_ ( .A(_05299_ ), .B(_01158_ ), .C1(_06092_ ), .C2(\mylsu.state [3] ), .ZN(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ) );
AND2_X1 _17019_ ( .A1(_03887_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ) );
NAND3_X1 _17020_ ( .A1(_06014_ ), .A2(_03844_ ), .A3(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .ZN(_01159_ ) );
OAI22_X1 _17021_ ( .A1(_05993_ ), .A2(_01159_ ), .B1(_06091_ ), .B2(_06021_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D ) );
AND2_X1 _17022_ ( .A1(_02045_ ), .A2(_03887_ ), .ZN(_01160_ ) );
INV_X1 _17023_ ( .A(io_master_wready ), .ZN(_01161_ ) );
NAND2_X1 _17024_ ( .A1(_01161_ ), .A2(_05986_ ), .ZN(_01162_ ) );
AND4_X1 _17025_ ( .A1(_01987_ ), .A2(_02055_ ), .A3(_01160_ ), .A4(_01162_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
NAND4_X1 _17026_ ( .A1(_03890_ ), .A2(\mylsu.state [2] ), .A3(_05985_ ), .A4(_01161_ ), .ZN(_01163_ ) );
AND2_X1 _17027_ ( .A1(io_master_wready ), .A2(io_master_awready ), .ZN(_01164_ ) );
NOR2_X1 _17028_ ( .A1(_03839_ ), .A2(_01164_ ), .ZN(_01165_ ) );
NAND4_X1 _17029_ ( .A1(_06077_ ), .A2(io_master_awready ), .A3(_03887_ ), .A4(_01165_ ), .ZN(_01166_ ) );
OAI21_X1 _17030_ ( .A(_01163_ ), .B1(_02079_ ), .B2(_01166_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D ) );
NOR2_X1 _17031_ ( .A1(_03839_ ), .A2(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_01167_ ) );
AND3_X1 _17032_ ( .A1(_01160_ ), .A2(\mylsu.state [0] ), .A3(_01167_ ), .ZN(_01168_ ) );
NAND3_X1 _17033_ ( .A1(_02055_ ), .A2(_01168_ ), .A3(_01164_ ), .ZN(_01169_ ) );
NAND3_X1 _17034_ ( .A1(_03887_ ), .A2(\mylsu.state [4] ), .A3(io_master_awready ), .ZN(_01170_ ) );
AND3_X1 _17035_ ( .A1(_03885_ ), .A2(io_master_wready ), .A3(_03065_ ), .ZN(_01171_ ) );
NAND2_X1 _17036_ ( .A1(_01171_ ), .A2(\mylsu.state [2] ), .ZN(_01172_ ) );
NAND3_X1 _17037_ ( .A1(_06087_ ), .A2(\mylsu.state [1] ), .A3(_03887_ ), .ZN(_01173_ ) );
NAND4_X1 _17038_ ( .A1(_01169_ ), .A2(_01170_ ), .A3(_01172_ ), .A4(_01173_ ), .ZN(\mylsu.state_$_DFF_P__Q_3_D ) );
NAND2_X1 _17039_ ( .A1(_06091_ ), .A2(_00283_ ), .ZN(_01174_ ) );
OAI211_X1 _17040_ ( .A(_06013_ ), .B(_02040_ ), .C1(_02023_ ), .C2(_02045_ ), .ZN(_01175_ ) );
NAND2_X1 _17041_ ( .A1(_01175_ ), .A2(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .ZN(_01176_ ) );
AND3_X1 _17042_ ( .A1(_02045_ ), .A2(\mylsu.state [0] ), .A3(_05986_ ), .ZN(_01177_ ) );
AND4_X1 _17043_ ( .A1(_01161_ ), .A2(_01177_ ), .A3(_05995_ ), .A4(_01165_ ), .ZN(_01178_ ) );
NAND2_X1 _17044_ ( .A1(_02055_ ), .A2(_01178_ ), .ZN(_01179_ ) );
OAI21_X1 _17045_ ( .A(_01168_ ), .B1(_02046_ ), .B2(_02054_ ), .ZN(_01180_ ) );
AOI221_X4 _17046_ ( .A(_05299_ ), .B1(\mylsu.state [0] ), .B2(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .C1(_06086_ ), .C2(\mylsu.state [1] ), .ZN(_01181_ ) );
AND4_X1 _17047_ ( .A1(_01176_ ), .A2(_01179_ ), .A3(_01180_ ), .A4(_01181_ ), .ZN(_01182_ ) );
OAI211_X1 _17048_ ( .A(_01174_ ), .B(_01182_ ), .C1(_05992_ ), .C2(_01159_ ), .ZN(\mylsu.state_$_DFF_P__Q_4_D ) );
NAND3_X1 _17049_ ( .A1(_03887_ ), .A2(\mylsu.state [4] ), .A3(_05986_ ), .ZN(_01183_ ) );
NAND3_X1 _17050_ ( .A1(_01177_ ), .A2(_01167_ ), .A3(_01171_ ), .ZN(_01184_ ) );
OAI21_X1 _17051_ ( .A(_01183_ ), .B1(_02079_ ), .B2(_01184_ ), .ZN(\mylsu.state_$_DFF_P__Q_D ) );
MUX2_X1 _17052_ ( .A(\LS_WB_wdata_csreg [21] ), .B(\EX_LS_result_csreg_mem [21] ), .S(_03834_ ), .Z(_01185_ ) );
NAND2_X2 _17053_ ( .A1(_03831_ ), .A2(_03840_ ), .ZN(_01186_ ) );
BUF_X4 _17054_ ( .A(_01186_ ), .Z(_01187_ ) );
MUX2_X1 _17055_ ( .A(_01185_ ), .B(\EX_LS_pc [21] ), .S(_01187_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ) );
AOI21_X1 _17056_ ( .A(\EX_LS_pc [20] ), .B1(_03832_ ), .B2(_03843_ ), .ZN(_01188_ ) );
BUF_X4 _17057_ ( .A(_05285_ ), .Z(_01189_ ) );
OAI21_X1 _17058_ ( .A(_03841_ ), .B1(_01189_ ), .B2(_06114_ ), .ZN(_01190_ ) );
BUF_X4 _17059_ ( .A(_05285_ ), .Z(_01191_ ) );
BUF_X4 _17060_ ( .A(_02045_ ), .Z(_01192_ ) );
AOI221_X4 _17061_ ( .A(_01190_ ), .B1(\LS_WB_wdata_csreg [20] ), .B2(_01191_ ), .C1(_02079_ ), .C2(_01192_ ), .ZN(_01193_ ) );
NOR2_X1 _17062_ ( .A1(_01188_ ), .A2(_01193_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _17063_ ( .A(\LS_WB_wdata_csreg [19] ), .B(\EX_LS_result_csreg_mem [19] ), .S(_03834_ ), .Z(_01194_ ) );
MUX2_X1 _17064_ ( .A(_01194_ ), .B(\EX_LS_pc [19] ), .S(_01187_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ) );
AOI21_X1 _17065_ ( .A(\EX_LS_pc [18] ), .B1(_03832_ ), .B2(_03843_ ), .ZN(_01195_ ) );
OAI21_X1 _17066_ ( .A(_03841_ ), .B1(_01189_ ), .B2(_06119_ ), .ZN(_01196_ ) );
AOI221_X4 _17067_ ( .A(_01196_ ), .B1(\LS_WB_wdata_csreg [18] ), .B2(_01191_ ), .C1(_02079_ ), .C2(_01192_ ), .ZN(_01197_ ) );
NOR2_X1 _17068_ ( .A1(_01195_ ), .A2(_01197_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _17069_ ( .A(\LS_WB_wdata_csreg [17] ), .B(\EX_LS_result_csreg_mem [17] ), .S(_03834_ ), .Z(_01198_ ) );
MUX2_X1 _17070_ ( .A(_01198_ ), .B(\EX_LS_pc [17] ), .S(_01187_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _17071_ ( .A(\LS_WB_wdata_csreg [16] ), .B(\EX_LS_result_csreg_mem [16] ), .S(_03834_ ), .Z(_01199_ ) );
MUX2_X1 _17072_ ( .A(_01199_ ), .B(\EX_LS_pc [16] ), .S(_01187_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ) );
AOI221_X4 _17073_ ( .A(_01186_ ), .B1(\LS_WB_wdata_csreg [15] ), .B2(_01191_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [15] ), .ZN(_01200_ ) );
BUF_X4 _17074_ ( .A(_03831_ ), .Z(_01201_ ) );
AOI21_X1 _17075_ ( .A(\EX_LS_pc [15] ), .B1(_01201_ ), .B2(_03842_ ), .ZN(_01202_ ) );
NOR2_X1 _17076_ ( .A1(_01200_ ), .A2(_01202_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ) );
AOI21_X1 _17077_ ( .A(\EX_LS_pc [14] ), .B1(_03832_ ), .B2(_03843_ ), .ZN(_01203_ ) );
OAI21_X1 _17078_ ( .A(_03841_ ), .B1(_01189_ ), .B2(_06134_ ), .ZN(_01204_ ) );
AOI221_X4 _17079_ ( .A(_01204_ ), .B1(\LS_WB_wdata_csreg [14] ), .B2(_01191_ ), .C1(_02079_ ), .C2(_01192_ ), .ZN(_01205_ ) );
NOR2_X1 _17080_ ( .A1(_01203_ ), .A2(_01205_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ) );
AOI21_X1 _17081_ ( .A(\EX_LS_pc [13] ), .B1(_03832_ ), .B2(_03843_ ), .ZN(_01206_ ) );
OAI21_X1 _17082_ ( .A(_03841_ ), .B1(_01189_ ), .B2(_06110_ ), .ZN(_01207_ ) );
AOI221_X4 _17083_ ( .A(_01207_ ), .B1(\LS_WB_wdata_csreg [13] ), .B2(_01191_ ), .C1(_02079_ ), .C2(_01192_ ), .ZN(_01208_ ) );
NOR2_X1 _17084_ ( .A1(_01206_ ), .A2(_01208_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _17085_ ( .A(\LS_WB_wdata_csreg [12] ), .B(\EX_LS_result_csreg_mem [12] ), .S(_03834_ ), .Z(_01209_ ) );
MUX2_X1 _17086_ ( .A(_01209_ ), .B(\EX_LS_pc [12] ), .S(_01187_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ) );
MUX2_X1 _17087_ ( .A(\LS_WB_wdata_csreg [30] ), .B(\EX_LS_result_csreg_mem [30] ), .S(_03833_ ), .Z(_01210_ ) );
MUX2_X1 _17088_ ( .A(_01210_ ), .B(\EX_LS_pc [30] ), .S(_01187_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ) );
OAI22_X1 _17089_ ( .A1(_03834_ ), .A2(_02077_ ), .B1(_02049_ ), .B2(_05580_ ), .ZN(_01211_ ) );
MUX2_X1 _17090_ ( .A(_01211_ ), .B(\EX_LS_pc [11] ), .S(_01187_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ) );
AOI21_X1 _17091_ ( .A(\EX_LS_pc [10] ), .B1(_03832_ ), .B2(_03843_ ), .ZN(_01212_ ) );
OAI21_X1 _17092_ ( .A(_03841_ ), .B1(_01189_ ), .B2(_06120_ ), .ZN(_01213_ ) );
AOI221_X4 _17093_ ( .A(_01213_ ), .B1(\LS_WB_wdata_csreg [10] ), .B2(_01191_ ), .C1(_02079_ ), .C2(_01192_ ), .ZN(_01214_ ) );
NOR2_X1 _17094_ ( .A1(_01212_ ), .A2(_01214_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _17095_ ( .A(\LS_WB_wdata_csreg [9] ), .B(\EX_LS_result_csreg_mem [9] ), .S(_03833_ ), .Z(_01215_ ) );
MUX2_X1 _17096_ ( .A(_01215_ ), .B(\EX_LS_pc [9] ), .S(_01187_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _17097_ ( .A(\LS_WB_wdata_csreg [8] ), .B(\EX_LS_result_csreg_mem [8] ), .S(_03833_ ), .Z(_01216_ ) );
MUX2_X1 _17098_ ( .A(_01216_ ), .B(\EX_LS_pc [8] ), .S(_01187_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ) );
AOI21_X1 _17099_ ( .A(\EX_LS_pc [7] ), .B1(_03832_ ), .B2(_03843_ ), .ZN(_01217_ ) );
OAI21_X1 _17100_ ( .A(_03841_ ), .B1(_05285_ ), .B2(_06106_ ), .ZN(_01218_ ) );
AOI221_X4 _17101_ ( .A(_01218_ ), .B1(\LS_WB_wdata_csreg [7] ), .B2(_01191_ ), .C1(_02079_ ), .C2(_01192_ ), .ZN(_01219_ ) );
NOR2_X1 _17102_ ( .A1(_01217_ ), .A2(_01219_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _17103_ ( .A(\LS_WB_wdata_csreg [6] ), .B(\EX_LS_result_csreg_mem [6] ), .S(_03833_ ), .Z(_01220_ ) );
MUX2_X1 _17104_ ( .A(_01220_ ), .B(\EX_LS_pc [6] ), .S(_01187_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ) );
AOI21_X1 _17105_ ( .A(\EX_LS_pc [5] ), .B1(_03832_ ), .B2(_03843_ ), .ZN(_01221_ ) );
OAI21_X1 _17106_ ( .A(_03841_ ), .B1(_05285_ ), .B2(_05724_ ), .ZN(_01222_ ) );
AOI221_X4 _17107_ ( .A(_01222_ ), .B1(\LS_WB_wdata_csreg [5] ), .B2(_01191_ ), .C1(_02079_ ), .C2(_01192_ ), .ZN(_01223_ ) );
NOR2_X1 _17108_ ( .A1(_01221_ ), .A2(_01223_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _17109_ ( .A(\LS_WB_wdata_csreg [4] ), .B(\EX_LS_result_csreg_mem [4] ), .S(_03833_ ), .Z(_01224_ ) );
MUX2_X1 _17110_ ( .A(_01224_ ), .B(\EX_LS_pc [4] ), .S(_01186_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _17111_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\EX_LS_result_csreg_mem [3] ), .S(_03833_ ), .Z(_01225_ ) );
MUX2_X1 _17112_ ( .A(_01225_ ), .B(\EX_LS_pc [3] ), .S(_01186_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ) );
AOI21_X1 _17113_ ( .A(\EX_LS_pc [2] ), .B1(_03832_ ), .B2(_03843_ ), .ZN(_01226_ ) );
OAI21_X1 _17114_ ( .A(_03841_ ), .B1(_05285_ ), .B2(_06097_ ), .ZN(_01227_ ) );
AOI221_X4 _17115_ ( .A(_01227_ ), .B1(\LS_WB_wdata_csreg [2] ), .B2(_01189_ ), .C1(_02056_ ), .C2(_01192_ ), .ZN(_01228_ ) );
NOR2_X1 _17116_ ( .A1(_01226_ ), .A2(_01228_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ) );
AOI221_X4 _17117_ ( .A(_01186_ ), .B1(\LS_WB_wdata_csreg [29] ), .B2(_01191_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [29] ), .ZN(_01229_ ) );
AOI21_X1 _17118_ ( .A(\EX_LS_pc [29] ), .B1(_01201_ ), .B2(_03842_ ), .ZN(_01230_ ) );
NOR2_X1 _17119_ ( .A1(_01229_ ), .A2(_01230_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ) );
AOI21_X1 _17120_ ( .A(\EX_LS_pc [1] ), .B1(_01201_ ), .B2(_03843_ ), .ZN(_01231_ ) );
OAI21_X1 _17121_ ( .A(_03841_ ), .B1(_05285_ ), .B2(_06098_ ), .ZN(_01232_ ) );
AOI221_X4 _17122_ ( .A(_01232_ ), .B1(\LS_WB_wdata_csreg [1] ), .B2(_01189_ ), .C1(_02056_ ), .C2(_01192_ ), .ZN(_01233_ ) );
NOR2_X1 _17123_ ( .A1(_01231_ ), .A2(_01233_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ) );
AOI221_X4 _17124_ ( .A(_01186_ ), .B1(_02049_ ), .B2(\LS_WB_wdata_csreg [0] ), .C1(\EX_LS_result_csreg_mem [0] ), .C2(_03834_ ), .ZN(_01234_ ) );
AOI21_X1 _17125_ ( .A(\EX_LS_pc [0] ), .B1(_01201_ ), .B2(_03842_ ), .ZN(_01235_ ) );
NOR2_X1 _17126_ ( .A1(_01234_ ), .A2(_01235_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ) );
AOI21_X1 _17127_ ( .A(\EX_LS_pc [28] ), .B1(_01201_ ), .B2(_03842_ ), .ZN(_01236_ ) );
OAI21_X1 _17128_ ( .A(_03840_ ), .B1(_05285_ ), .B2(_07867_ ), .ZN(_01237_ ) );
AOI221_X4 _17129_ ( .A(_01237_ ), .B1(\LS_WB_wdata_csreg [28] ), .B2(_01189_ ), .C1(_02056_ ), .C2(_01192_ ), .ZN(_01238_ ) );
NOR2_X1 _17130_ ( .A1(_01236_ ), .A2(_01238_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ) );
AOI21_X1 _17131_ ( .A(\EX_LS_pc [27] ), .B1(_01201_ ), .B2(_03842_ ), .ZN(_01239_ ) );
OAI21_X1 _17132_ ( .A(_03840_ ), .B1(_05285_ ), .B2(_05815_ ), .ZN(_01240_ ) );
AOI221_X4 _17133_ ( .A(_01240_ ), .B1(\LS_WB_wdata_csreg [27] ), .B2(_01189_ ), .C1(_02056_ ), .C2(_02045_ ), .ZN(_01241_ ) );
NOR2_X1 _17134_ ( .A1(_01239_ ), .A2(_01241_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ) );
AOI21_X1 _17135_ ( .A(\EX_LS_pc [26] ), .B1(_01201_ ), .B2(_03842_ ), .ZN(_01242_ ) );
MUX2_X1 _17136_ ( .A(\LS_WB_wdata_csreg [26] ), .B(\EX_LS_result_csreg_mem [26] ), .S(_03833_ ), .Z(_01243_ ) );
NOR4_X1 _17137_ ( .A1(_03830_ ), .A2(_03839_ ), .A3(_03837_ ), .A4(_01243_ ), .ZN(_01244_ ) );
NOR2_X1 _17138_ ( .A1(_01242_ ), .A2(_01244_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ) );
AOI221_X4 _17139_ ( .A(_01186_ ), .B1(\LS_WB_wdata_csreg [25] ), .B2(_01191_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [25] ), .ZN(_01245_ ) );
AOI21_X1 _17140_ ( .A(\EX_LS_pc [25] ), .B1(_01201_ ), .B2(_03842_ ), .ZN(_01246_ ) );
NOR2_X1 _17141_ ( .A1(_01245_ ), .A2(_01246_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ) );
AOI21_X1 _17142_ ( .A(\EX_LS_pc [24] ), .B1(_01201_ ), .B2(_03842_ ), .ZN(_01247_ ) );
OAI21_X1 _17143_ ( .A(_03840_ ), .B1(_05285_ ), .B2(_05888_ ), .ZN(_01248_ ) );
AOI221_X4 _17144_ ( .A(_01248_ ), .B1(\LS_WB_wdata_csreg [24] ), .B2(_01189_ ), .C1(_02056_ ), .C2(_02045_ ), .ZN(_01249_ ) );
NOR2_X1 _17145_ ( .A1(_01247_ ), .A2(_01249_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _17146_ ( .A(\LS_WB_wdata_csreg [23] ), .B(\EX_LS_result_csreg_mem [23] ), .S(_03833_ ), .Z(_01250_ ) );
MUX2_X1 _17147_ ( .A(_01250_ ), .B(\EX_LS_pc [23] ), .S(_01186_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ) );
OAI22_X1 _17148_ ( .A1(_03834_ ), .A2(_02078_ ), .B1(_02049_ ), .B2(_05919_ ), .ZN(_01251_ ) );
MUX2_X1 _17149_ ( .A(_01251_ ), .B(\EX_LS_pc [22] ), .S(_01186_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ) );
AOI21_X1 _17150_ ( .A(\EX_LS_pc [31] ), .B1(_01201_ ), .B2(_03842_ ), .ZN(_01252_ ) );
MUX2_X1 _17151_ ( .A(\LS_WB_wdata_csreg [31] ), .B(\EX_LS_result_csreg_mem [31] ), .S(_03833_ ), .Z(_01253_ ) );
NOR4_X1 _17152_ ( .A1(_03830_ ), .A2(_03839_ ), .A3(_03837_ ), .A4(_01253_ ), .ZN(_01254_ ) );
NOR2_X1 _17153_ ( .A1(_01252_ ), .A2(_01254_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ) );
BUF_X2 _17154_ ( .A(_05990_ ), .Z(_01255_ ) );
NOR2_X1 _17155_ ( .A1(_00543_ ), .A2(_01255_ ), .ZN(_01256_ ) );
NOR2_X1 _17156_ ( .A1(_00515_ ), .A2(_05990_ ), .ZN(_01257_ ) );
NOR2_X1 _17157_ ( .A1(_00484_ ), .A2(_05990_ ), .ZN(_01258_ ) );
NOR2_X1 _17158_ ( .A1(_00582_ ), .A2(_05990_ ), .ZN(_01259_ ) );
NOR2_X1 _17159_ ( .A1(_06029_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01260_ ) );
MUX2_X2 _17160_ ( .A(_01258_ ), .B(_01259_ ), .S(_01260_ ), .Z(_01261_ ) );
NOR2_X1 _17161_ ( .A1(_06032_ ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01262_ ) );
INV_X1 _17162_ ( .A(_01262_ ), .ZN(_01263_ ) );
MUX2_X2 _17163_ ( .A(_01257_ ), .B(_01261_ ), .S(_01263_ ), .Z(_01264_ ) );
NOR2_X2 _17164_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01265_ ) );
INV_X1 _17165_ ( .A(_01265_ ), .ZN(_01266_ ) );
MUX2_X2 _17166_ ( .A(_01256_ ), .B(_01264_ ), .S(_01266_ ), .Z(_01267_ ) );
NOR2_X1 _17167_ ( .A1(\mylsu.typ_tmp [0] ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01268_ ) );
AND2_X1 _17168_ ( .A1(_01268_ ), .A2(\mylsu.typ_tmp_$_NOT__A_Y ), .ZN(_01269_ ) );
BUF_X4 _17169_ ( .A(_01269_ ), .Z(_01270_ ) );
AND2_X4 _17170_ ( .A1(_01267_ ), .A2(_01270_ ), .ZN(_01271_ ) );
MUX2_X1 _17171_ ( .A(_01258_ ), .B(_01257_ ), .S(_01265_ ), .Z(_01272_ ) );
AND2_X1 _17172_ ( .A1(\mylsu.typ_tmp_$_NOT__A_Y ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01273_ ) );
INV_X1 _17173_ ( .A(\mylsu.typ_tmp [0] ), .ZN(_01274_ ) );
AND2_X2 _17174_ ( .A1(_01273_ ), .A2(_01274_ ), .ZN(_01275_ ) );
INV_X1 _17175_ ( .A(_01275_ ), .ZN(_01276_ ) );
OR2_X4 _17176_ ( .A1(_01272_ ), .A2(_01276_ ), .ZN(_01277_ ) );
BUF_X2 _17177_ ( .A(_01273_ ), .Z(_01278_ ) );
AND2_X1 _17178_ ( .A1(_01278_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01279_ ) );
BUF_X4 _17179_ ( .A(_01279_ ), .Z(_01280_ ) );
NOR4_X1 _17180_ ( .A1(_00494_ ), .A2(_00495_ ), .A3(_05991_ ), .A4(_01280_ ), .ZN(_01281_ ) );
OR2_X1 _17181_ ( .A1(_01281_ ), .A2(_01275_ ), .ZN(_01282_ ) );
OR2_X1 _17182_ ( .A1(_01274_ ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01283_ ) );
NOR2_X1 _17183_ ( .A1(_01283_ ), .A2(\mylsu.typ_tmp [2] ), .ZN(_01284_ ) );
NOR2_X1 _17184_ ( .A1(_01284_ ), .A2(_01269_ ), .ZN(_01285_ ) );
AND3_X1 _17185_ ( .A1(_01277_ ), .A2(_01282_ ), .A3(_01285_ ), .ZN(_01286_ ) );
OAI21_X1 _17186_ ( .A(\mylsu.state [3] ), .B1(_01271_ ), .B2(_01286_ ), .ZN(_01287_ ) );
OAI21_X1 _17187_ ( .A(_01287_ ), .B1(\mylsu.state [3] ), .B2(_04508_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ) );
OR2_X1 _17188_ ( .A1(_00499_ ), .A2(_05991_ ), .ZN(_01288_ ) );
OAI21_X1 _17189_ ( .A(_01276_ ), .B1(_01288_ ), .B2(_01280_ ), .ZN(_01289_ ) );
AND3_X1 _17190_ ( .A1(_01277_ ), .A2(_01285_ ), .A3(_01289_ ), .ZN(_01290_ ) );
OR2_X4 _17191_ ( .A1(_01271_ ), .A2(_01290_ ), .ZN(_01291_ ) );
MUX2_X2 _17192_ ( .A(\EX_LS_result_reg [20] ), .B(_01291_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ) );
NAND3_X1 _17193_ ( .A1(_00500_ ), .A2(_00502_ ), .A3(\io_master_arid [1] ), .ZN(_01292_ ) );
OAI21_X1 _17194_ ( .A(_01276_ ), .B1(_01292_ ), .B2(_01280_ ), .ZN(_01293_ ) );
AND3_X1 _17195_ ( .A1(_01277_ ), .A2(_01285_ ), .A3(_01293_ ), .ZN(_01294_ ) );
OAI21_X1 _17196_ ( .A(\mylsu.state [3] ), .B1(_01271_ ), .B2(_01294_ ), .ZN(_01295_ ) );
OAI21_X1 _17197_ ( .A(_01295_ ), .B1(\mylsu.state [3] ), .B2(_04384_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ) );
NAND3_X1 _17198_ ( .A1(_00503_ ), .A2(_00506_ ), .A3(_06073_ ), .ZN(_01296_ ) );
OAI21_X1 _17199_ ( .A(_01276_ ), .B1(_01296_ ), .B2(_01280_ ), .ZN(_01297_ ) );
AND3_X1 _17200_ ( .A1(_01277_ ), .A2(_01285_ ), .A3(_01297_ ), .ZN(_01298_ ) );
OR2_X4 _17201_ ( .A1(_01271_ ), .A2(_01298_ ), .ZN(_01299_ ) );
MUX2_X2 _17202_ ( .A(\EX_LS_result_reg [18] ), .B(_01299_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ) );
NAND3_X1 _17203_ ( .A1(_00507_ ), .A2(_00509_ ), .A3(\io_master_arid [1] ), .ZN(_01300_ ) );
OAI21_X1 _17204_ ( .A(_01276_ ), .B1(_01300_ ), .B2(_01280_ ), .ZN(_01301_ ) );
AND3_X1 _17205_ ( .A1(_01277_ ), .A2(_01285_ ), .A3(_01301_ ), .ZN(_01302_ ) );
OAI21_X1 _17206_ ( .A(\mylsu.state [3] ), .B1(_01271_ ), .B2(_01302_ ), .ZN(_01303_ ) );
OAI21_X1 _17207_ ( .A(_01303_ ), .B1(\mylsu.state [3] ), .B2(_04427_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ) );
NAND3_X1 _17208_ ( .A1(_00510_ ), .A2(_00512_ ), .A3(_06073_ ), .ZN(_01304_ ) );
OAI21_X1 _17209_ ( .A(_01276_ ), .B1(_01304_ ), .B2(_01280_ ), .ZN(_01305_ ) );
AND3_X1 _17210_ ( .A1(_01277_ ), .A2(_01285_ ), .A3(_01305_ ), .ZN(_01306_ ) );
OR2_X4 _17211_ ( .A1(_01271_ ), .A2(_01306_ ), .ZN(_01307_ ) );
MUX2_X2 _17212_ ( .A(\EX_LS_result_reg [16] ), .B(_01307_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ) );
NOR2_X2 _17213_ ( .A1(_01271_ ), .A2(_01157_ ), .ZN(_01308_ ) );
AND2_X1 _17214_ ( .A1(_01272_ ), .A2(_01278_ ), .ZN(_01309_ ) );
NOR3_X1 _17215_ ( .A1(_01284_ ), .A2(_01270_ ), .A3(_01278_ ), .ZN(_01310_ ) );
AOI21_X1 _17216_ ( .A(_01309_ ), .B1(_01257_ ), .B2(_01310_ ), .ZN(_01311_ ) );
BUF_X4 _17217_ ( .A(_01157_ ), .Z(_01312_ ) );
AOI22_X1 _17218_ ( .A1(_01308_ ), .A2(_01311_ ), .B1(_01312_ ), .B2(_04110_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ) );
INV_X4 _17219_ ( .A(_01271_ ), .ZN(_01313_ ) );
NAND2_X1 _17220_ ( .A1(_01266_ ), .A2(_01278_ ), .ZN(_01314_ ) );
OR3_X1 _17221_ ( .A1(_00492_ ), .A2(_06027_ ), .A3(_01314_ ), .ZN(_01315_ ) );
NAND2_X1 _17222_ ( .A1(_01285_ ), .A2(_01314_ ), .ZN(_01316_ ) );
NOR2_X1 _17223_ ( .A1(_05991_ ), .A2(_01316_ ), .ZN(_01317_ ) );
NAND3_X1 _17224_ ( .A1(_00516_ ), .A2(_00518_ ), .A3(_01317_ ), .ZN(_01318_ ) );
NAND3_X1 _17225_ ( .A1(_01313_ ), .A2(_01315_ ), .A3(_01318_ ), .ZN(_01319_ ) );
MUX2_X1 _17226_ ( .A(\EX_LS_result_reg [14] ), .B(_01319_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ) );
INV_X1 _17227_ ( .A(_01278_ ), .ZN(_01320_ ) );
NOR2_X1 _17228_ ( .A1(_01320_ ), .A2(_01265_ ), .ZN(_01321_ ) );
AND4_X1 _17229_ ( .A1(\io_master_arid [1] ), .A2(_00526_ ), .A3(_00528_ ), .A4(_01321_ ), .ZN(_01322_ ) );
AND3_X1 _17230_ ( .A1(_00520_ ), .A2(_00522_ ), .A3(_01317_ ), .ZN(_01323_ ) );
NOR2_X1 _17231_ ( .A1(_01322_ ), .A2(_01323_ ), .ZN(_01324_ ) );
AOI22_X1 _17232_ ( .A1(_01308_ ), .A2(_01324_ ), .B1(_01312_ ), .B2(_04051_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ) );
AND3_X1 _17233_ ( .A1(_00523_ ), .A2(_00525_ ), .A3(_01317_ ), .ZN(_01325_ ) );
NOR2_X1 _17234_ ( .A1(_00561_ ), .A2(_06028_ ), .ZN(_01326_ ) );
AOI21_X1 _17235_ ( .A(_01325_ ), .B1(_01326_ ), .B2(_01321_ ), .ZN(_01327_ ) );
AOI22_X1 _17236_ ( .A1(_01308_ ), .A2(_01327_ ), .B1(_01312_ ), .B2(_04080_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ) );
AND2_X1 _17237_ ( .A1(_01277_ ), .A2(_01285_ ), .ZN(_01328_ ) );
BUF_X4 _17238_ ( .A(_01328_ ), .Z(_01329_ ) );
BUF_X4 _17239_ ( .A(_01275_ ), .Z(_01330_ ) );
NOR3_X1 _17240_ ( .A1(_00492_ ), .A2(_06027_ ), .A3(_01278_ ), .ZN(_01331_ ) );
OAI21_X1 _17241_ ( .A(_01329_ ), .B1(_01330_ ), .B2(_01331_ ), .ZN(_01332_ ) );
NAND2_X1 _17242_ ( .A1(_01313_ ), .A2(_01332_ ), .ZN(_01333_ ) );
MUX2_X1 _17243_ ( .A(\EX_LS_result_reg [30] ), .B(_01333_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ) );
NAND4_X1 _17244_ ( .A1(_00568_ ), .A2(_00570_ ), .A3(\io_master_arid [1] ), .A4(_01321_ ), .ZN(_01334_ ) );
NAND3_X1 _17245_ ( .A1(_00529_ ), .A2(_00531_ ), .A3(_01317_ ), .ZN(_01335_ ) );
AND2_X1 _17246_ ( .A1(_01334_ ), .A2(_01335_ ), .ZN(_01336_ ) );
AOI22_X1 _17247_ ( .A1(_01308_ ), .A2(_01336_ ), .B1(_01312_ ), .B2(_03926_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ) );
AND3_X1 _17248_ ( .A1(_00532_ ), .A2(_00534_ ), .A3(_01317_ ), .ZN(_01337_ ) );
AND4_X1 _17249_ ( .A1(_06073_ ), .A2(_00571_ ), .A3(_00573_ ), .A4(_01321_ ), .ZN(_01338_ ) );
OR3_X4 _17250_ ( .A1(_01271_ ), .A2(_01337_ ), .A3(_01338_ ), .ZN(_01339_ ) );
MUX2_X2 _17251_ ( .A(\EX_LS_result_reg [10] ), .B(_01339_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ) );
NAND4_X1 _17252_ ( .A1(_00574_ ), .A2(_00576_ ), .A3(\io_master_arid [1] ), .A4(_01321_ ), .ZN(_01340_ ) );
NAND3_X1 _17253_ ( .A1(_00535_ ), .A2(_00537_ ), .A3(_01317_ ), .ZN(_01341_ ) );
AND2_X1 _17254_ ( .A1(_01340_ ), .A2(_01341_ ), .ZN(_01342_ ) );
AOI22_X1 _17255_ ( .A1(_01308_ ), .A2(_01342_ ), .B1(_01312_ ), .B2(_04025_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ) );
AND3_X1 _17256_ ( .A1(_00538_ ), .A2(_00540_ ), .A3(_01317_ ), .ZN(_01343_ ) );
AND4_X1 _17257_ ( .A1(_06073_ ), .A2(_00577_ ), .A3(_00579_ ), .A4(_01321_ ), .ZN(_01344_ ) );
OR3_X4 _17258_ ( .A1(_01271_ ), .A2(_01343_ ), .A3(_01344_ ), .ZN(_01345_ ) );
MUX2_X2 _17259_ ( .A(\EX_LS_result_reg [8] ), .B(_01345_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ) );
NAND2_X1 _17260_ ( .A1(_01157_ ), .A2(\EX_LS_result_reg [7] ), .ZN(_01346_ ) );
NOR2_X1 _17261_ ( .A1(_01267_ ), .A2(_01285_ ), .ZN(_01347_ ) );
OAI221_X1 _17262_ ( .A(\mylsu.state [3] ), .B1(_01259_ ), .B2(_01314_ ), .C1(_01256_ ), .C2(_01316_ ), .ZN(_01348_ ) );
OAI21_X1 _17263_ ( .A(_01346_ ), .B1(_01347_ ), .B2(_01348_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ) );
INV_X1 _17264_ ( .A(_01260_ ), .ZN(_01349_ ) );
NOR3_X1 _17265_ ( .A1(_00585_ ), .A2(_05991_ ), .A3(_01349_ ), .ZN(_01350_ ) );
NOR3_X1 _17266_ ( .A1(_00492_ ), .A2(_01255_ ), .A3(_01260_ ), .ZN(_01351_ ) );
OAI21_X1 _17267_ ( .A(_01263_ ), .B1(_01350_ ), .B2(_01351_ ), .ZN(_01352_ ) );
NAND4_X1 _17268_ ( .A1(_00516_ ), .A2(_00518_ ), .A3(_06073_ ), .A4(_01262_ ), .ZN(_01353_ ) );
AOI21_X1 _17269_ ( .A(_01265_ ), .B1(_01352_ ), .B2(_01353_ ), .ZN(_01354_ ) );
NOR3_X1 _17270_ ( .A1(_00546_ ), .A2(_01255_ ), .A3(_01266_ ), .ZN(_01355_ ) );
OAI21_X1 _17271_ ( .A(_01270_ ), .B1(_01354_ ), .B2(_01355_ ), .ZN(_01356_ ) );
NOR3_X1 _17272_ ( .A1(_00585_ ), .A2(_01255_ ), .A3(_01265_ ), .ZN(_01357_ ) );
OAI21_X1 _17273_ ( .A(_01280_ ), .B1(_01357_ ), .B2(_01355_ ), .ZN(_01358_ ) );
OR3_X1 _17274_ ( .A1(_00546_ ), .A2(_05991_ ), .A3(_01279_ ), .ZN(_01359_ ) );
AOI21_X1 _17275_ ( .A(_01275_ ), .B1(_01358_ ), .B2(_01359_ ), .ZN(_01360_ ) );
INV_X1 _17276_ ( .A(_01357_ ), .ZN(_01361_ ) );
INV_X1 _17277_ ( .A(_01355_ ), .ZN(_01362_ ) );
AOI21_X1 _17278_ ( .A(_01276_ ), .B1(_01361_ ), .B2(_01362_ ), .ZN(_01363_ ) );
OAI22_X1 _17279_ ( .A1(_01360_ ), .A2(_01363_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01283_ ), .ZN(_01364_ ) );
OAI21_X1 _17280_ ( .A(_01284_ ), .B1(_01354_ ), .B2(_01355_ ), .ZN(_01365_ ) );
AND2_X1 _17281_ ( .A1(_01364_ ), .A2(_01365_ ), .ZN(_01366_ ) );
OAI21_X1 _17282_ ( .A(_01356_ ), .B1(_01366_ ), .B2(_01270_ ), .ZN(_01367_ ) );
MUX2_X1 _17283_ ( .A(\EX_LS_result_reg [6] ), .B(_01367_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ) );
NAND2_X1 _17284_ ( .A1(_01157_ ), .A2(\EX_LS_result_reg [5] ), .ZN(_01368_ ) );
NOR2_X1 _17285_ ( .A1(_01310_ ), .A2(_01265_ ), .ZN(_01369_ ) );
INV_X1 _17286_ ( .A(_01369_ ), .ZN(_01370_ ) );
AOI211_X1 _17287_ ( .A(_01157_ ), .B(_06027_ ), .C1(_00549_ ), .C2(_01370_ ), .ZN(_01371_ ) );
NOR2_X1 _17288_ ( .A1(_01285_ ), .A2(_06032_ ), .ZN(_01372_ ) );
INV_X1 _17289_ ( .A(_01372_ ), .ZN(_01373_ ) );
AND2_X1 _17290_ ( .A1(_01373_ ), .A2(_01369_ ), .ZN(_01374_ ) );
OAI21_X1 _17291_ ( .A(_01374_ ), .B1(_00494_ ), .B2(_00495_ ), .ZN(_01375_ ) );
NAND2_X1 _17292_ ( .A1(_01371_ ), .A2(_01375_ ), .ZN(_01376_ ) );
OAI211_X1 _17293_ ( .A(_00522_ ), .B(_06029_ ), .C1(\io_master_rdata [13] ), .C2(_03814_ ), .ZN(_01377_ ) );
NAND3_X1 _17294_ ( .A1(_00526_ ), .A2(_00528_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01378_ ) );
AND3_X1 _17295_ ( .A1(_01377_ ), .A2(_01372_ ), .A3(_01378_ ), .ZN(_01379_ ) );
OAI21_X1 _17296_ ( .A(_01368_ ), .B1(_01376_ ), .B2(_01379_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ) );
NOR3_X1 _17297_ ( .A1(_00561_ ), .A2(_05991_ ), .A3(_01260_ ), .ZN(_01380_ ) );
NOR3_X1 _17298_ ( .A1(_00499_ ), .A2(_01255_ ), .A3(_01349_ ), .ZN(_01381_ ) );
OAI21_X1 _17299_ ( .A(_01263_ ), .B1(_01380_ ), .B2(_01381_ ), .ZN(_01382_ ) );
NAND4_X1 _17300_ ( .A1(_00523_ ), .A2(_00525_ ), .A3(_06073_ ), .A4(_01262_ ), .ZN(_01383_ ) );
AOI21_X1 _17301_ ( .A(_01265_ ), .B1(_01382_ ), .B2(_01383_ ), .ZN(_01384_ ) );
NOR3_X1 _17302_ ( .A1(_00552_ ), .A2(_01255_ ), .A3(_01266_ ), .ZN(_01385_ ) );
OAI21_X1 _17303_ ( .A(_01270_ ), .B1(_01384_ ), .B2(_01385_ ), .ZN(_01386_ ) );
NOR3_X1 _17304_ ( .A1(_00499_ ), .A2(_01255_ ), .A3(_01265_ ), .ZN(_01387_ ) );
OAI21_X1 _17305_ ( .A(_01280_ ), .B1(_01387_ ), .B2(_01385_ ), .ZN(_01388_ ) );
OR3_X1 _17306_ ( .A1(_00552_ ), .A2(_05991_ ), .A3(_01279_ ), .ZN(_01389_ ) );
AOI21_X1 _17307_ ( .A(_01275_ ), .B1(_01388_ ), .B2(_01389_ ), .ZN(_01390_ ) );
INV_X1 _17308_ ( .A(_01387_ ), .ZN(_01391_ ) );
INV_X1 _17309_ ( .A(_01385_ ), .ZN(_01392_ ) );
AOI21_X1 _17310_ ( .A(_01276_ ), .B1(_01391_ ), .B2(_01392_ ), .ZN(_01393_ ) );
OAI22_X1 _17311_ ( .A1(_01390_ ), .A2(_01393_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01283_ ), .ZN(_01394_ ) );
OAI21_X1 _17312_ ( .A(_01284_ ), .B1(_01384_ ), .B2(_01385_ ), .ZN(_01395_ ) );
AND2_X1 _17313_ ( .A1(_01394_ ), .A2(_01395_ ), .ZN(_01396_ ) );
OAI21_X1 _17314_ ( .A(_01386_ ), .B1(_01396_ ), .B2(_01270_ ), .ZN(_01397_ ) );
MUX2_X1 _17315_ ( .A(\EX_LS_result_reg [4] ), .B(_01397_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ) );
AND4_X1 _17316_ ( .A1(_01966_ ), .A2(_00568_ ), .A3(_00570_ ), .A4(_01349_ ), .ZN(_01398_ ) );
AND4_X1 _17317_ ( .A1(_01966_ ), .A2(_00500_ ), .A3(_00502_ ), .A4(_01260_ ), .ZN(_01399_ ) );
OAI21_X1 _17318_ ( .A(_01263_ ), .B1(_01398_ ), .B2(_01399_ ), .ZN(_01400_ ) );
NAND4_X1 _17319_ ( .A1(_00529_ ), .A2(_00531_ ), .A3(_06073_ ), .A4(_01262_ ), .ZN(_01401_ ) );
AOI21_X1 _17320_ ( .A(_01265_ ), .B1(_01400_ ), .B2(_01401_ ), .ZN(_01402_ ) );
NOR3_X1 _17321_ ( .A1(_00555_ ), .A2(_01255_ ), .A3(_01266_ ), .ZN(_01403_ ) );
OAI21_X1 _17322_ ( .A(_01270_ ), .B1(_01402_ ), .B2(_01403_ ), .ZN(_01404_ ) );
AND4_X1 _17323_ ( .A1(_01966_ ), .A2(_00500_ ), .A3(_00502_ ), .A4(_01266_ ), .ZN(_01405_ ) );
OR2_X1 _17324_ ( .A1(_01403_ ), .A2(_01405_ ), .ZN(_01406_ ) );
AND2_X1 _17325_ ( .A1(_01406_ ), .A2(_01275_ ), .ZN(_01407_ ) );
OAI21_X1 _17326_ ( .A(_01280_ ), .B1(_01403_ ), .B2(_01405_ ), .ZN(_01408_ ) );
OR3_X1 _17327_ ( .A1(_00555_ ), .A2(_05991_ ), .A3(_01279_ ), .ZN(_01409_ ) );
AOI21_X1 _17328_ ( .A(_01275_ ), .B1(_01408_ ), .B2(_01409_ ), .ZN(_01410_ ) );
OAI22_X1 _17329_ ( .A1(_01407_ ), .A2(_01410_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01283_ ), .ZN(_01411_ ) );
OAI21_X1 _17330_ ( .A(_01284_ ), .B1(_01402_ ), .B2(_01403_ ), .ZN(_01412_ ) );
AND2_X1 _17331_ ( .A1(_01411_ ), .A2(_01412_ ), .ZN(_01413_ ) );
OAI21_X1 _17332_ ( .A(_01404_ ), .B1(_01413_ ), .B2(_01270_ ), .ZN(_01414_ ) );
MUX2_X1 _17333_ ( .A(\EX_LS_result_reg [3] ), .B(_01414_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ) );
AND2_X1 _17334_ ( .A1(_00558_ ), .A2(_01370_ ), .ZN(_01415_ ) );
INV_X1 _17335_ ( .A(_01374_ ), .ZN(_01416_ ) );
AOI21_X1 _17336_ ( .A(_01416_ ), .B1(_00503_ ), .B2(_00506_ ), .ZN(_01417_ ) );
OR4_X1 _17337_ ( .A1(_01157_ ), .A2(_01415_ ), .A3(_06027_ ), .A4(_01417_ ), .ZN(_01418_ ) );
OAI211_X1 _17338_ ( .A(_00534_ ), .B(_06029_ ), .C1(\io_master_rdata [10] ), .C2(_03814_ ), .ZN(_01419_ ) );
NAND3_X1 _17339_ ( .A1(_00571_ ), .A2(_00573_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01420_ ) );
AND3_X1 _17340_ ( .A1(_01419_ ), .A2(_01372_ ), .A3(_01420_ ), .ZN(_01421_ ) );
OAI22_X1 _17341_ ( .A1(_01418_ ), .A2(_01421_ ), .B1(\mylsu.state [3] ), .B2(_04302_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ) );
AND4_X1 _17342_ ( .A1(_06073_ ), .A2(_00526_ ), .A3(_00528_ ), .A4(_01320_ ), .ZN(_01422_ ) );
OAI21_X1 _17343_ ( .A(_01329_ ), .B1(_01330_ ), .B2(_01422_ ), .ZN(_01423_ ) );
NAND2_X1 _17344_ ( .A1(_01313_ ), .A2(_01423_ ), .ZN(_01424_ ) );
MUX2_X1 _17345_ ( .A(\EX_LS_result_reg [29] ), .B(_01424_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ) );
AND4_X1 _17346_ ( .A1(_01966_ ), .A2(_00574_ ), .A3(_00576_ ), .A4(_01349_ ), .ZN(_01425_ ) );
AND4_X1 _17347_ ( .A1(_01966_ ), .A2(_00507_ ), .A3(_00509_ ), .A4(_01260_ ), .ZN(_01426_ ) );
OAI21_X1 _17348_ ( .A(_01263_ ), .B1(_01425_ ), .B2(_01426_ ), .ZN(_01427_ ) );
NAND4_X1 _17349_ ( .A1(_00535_ ), .A2(_00537_ ), .A3(_01966_ ), .A4(_01262_ ), .ZN(_01428_ ) );
AOI21_X1 _17350_ ( .A(_01265_ ), .B1(_01427_ ), .B2(_01428_ ), .ZN(_01429_ ) );
NOR3_X1 _17351_ ( .A1(_00564_ ), .A2(_01255_ ), .A3(_01266_ ), .ZN(_01430_ ) );
OAI21_X1 _17352_ ( .A(_01270_ ), .B1(_01429_ ), .B2(_01430_ ), .ZN(_01431_ ) );
AND4_X1 _17353_ ( .A1(_01966_ ), .A2(_00507_ ), .A3(_00509_ ), .A4(_01266_ ), .ZN(_01432_ ) );
OR2_X1 _17354_ ( .A1(_01430_ ), .A2(_01432_ ), .ZN(_01433_ ) );
AND2_X1 _17355_ ( .A1(_01433_ ), .A2(_01275_ ), .ZN(_01434_ ) );
OAI21_X1 _17356_ ( .A(_01280_ ), .B1(_01430_ ), .B2(_01432_ ), .ZN(_01435_ ) );
OR3_X1 _17357_ ( .A1(_00564_ ), .A2(_01255_ ), .A3(_01279_ ), .ZN(_01436_ ) );
AOI21_X1 _17358_ ( .A(_01275_ ), .B1(_01435_ ), .B2(_01436_ ), .ZN(_01437_ ) );
OAI22_X1 _17359_ ( .A1(_01434_ ), .A2(_01437_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01283_ ), .ZN(_01438_ ) );
OAI21_X1 _17360_ ( .A(_01284_ ), .B1(_01429_ ), .B2(_01430_ ), .ZN(_01439_ ) );
AND2_X1 _17361_ ( .A1(_01438_ ), .A2(_01439_ ), .ZN(_01440_ ) );
OAI21_X1 _17362_ ( .A(_01431_ ), .B1(_01440_ ), .B2(_01270_ ), .ZN(_01441_ ) );
MUX2_X1 _17363_ ( .A(\EX_LS_result_reg [1] ), .B(_01441_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ) );
NAND2_X1 _17364_ ( .A1(_01157_ ), .A2(\EX_LS_result_reg [0] ), .ZN(_01442_ ) );
AND2_X1 _17365_ ( .A1(_00567_ ), .A2(_01370_ ), .ZN(_01443_ ) );
AOI21_X1 _17366_ ( .A(_01416_ ), .B1(_00510_ ), .B2(_00512_ ), .ZN(_01444_ ) );
OR4_X1 _17367_ ( .A1(_01157_ ), .A2(_01443_ ), .A3(_06027_ ), .A4(_01444_ ), .ZN(_01445_ ) );
OAI211_X1 _17368_ ( .A(_00540_ ), .B(_06029_ ), .C1(\io_master_rdata [8] ), .C2(_03814_ ), .ZN(_01446_ ) );
NAND3_X1 _17369_ ( .A1(_00577_ ), .A2(_00579_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01447_ ) );
AND3_X1 _17370_ ( .A1(_01446_ ), .A2(_01372_ ), .A3(_01447_ ), .ZN(_01448_ ) );
OAI21_X1 _17371_ ( .A(_01442_ ), .B1(_01445_ ), .B2(_01448_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ) );
NOR3_X1 _17372_ ( .A1(_00561_ ), .A2(_06027_ ), .A3(_01278_ ), .ZN(_01449_ ) );
OAI21_X1 _17373_ ( .A(_01329_ ), .B1(_01330_ ), .B2(_01449_ ), .ZN(_01450_ ) );
NAND2_X1 _17374_ ( .A1(_01313_ ), .A2(_01450_ ), .ZN(_01451_ ) );
MUX2_X1 _17375_ ( .A(\EX_LS_result_reg [28] ), .B(_01451_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ) );
AND4_X1 _17376_ ( .A1(\io_master_arid [1] ), .A2(_00568_ ), .A3(_00570_ ), .A4(_01320_ ), .ZN(_01452_ ) );
OAI21_X1 _17377_ ( .A(_01329_ ), .B1(_01330_ ), .B2(_01452_ ), .ZN(_01453_ ) );
AOI22_X1 _17378_ ( .A1(_01308_ ), .A2(_01453_ ), .B1(_01312_ ), .B2(_04704_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ) );
AND4_X1 _17379_ ( .A1(\io_master_arid [1] ), .A2(_00571_ ), .A3(_00573_ ), .A4(_01320_ ), .ZN(_01454_ ) );
OAI21_X1 _17380_ ( .A(_01329_ ), .B1(_01330_ ), .B2(_01454_ ), .ZN(_01455_ ) );
AOI22_X1 _17381_ ( .A1(_01308_ ), .A2(_01455_ ), .B1(_01312_ ), .B2(_04682_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ) );
AND4_X1 _17382_ ( .A1(\io_master_arid [1] ), .A2(_00574_ ), .A3(_00576_ ), .A4(_01320_ ), .ZN(_01456_ ) );
OAI21_X1 _17383_ ( .A(_01329_ ), .B1(_01330_ ), .B2(_01456_ ), .ZN(_01457_ ) );
AOI22_X1 _17384_ ( .A1(_01308_ ), .A2(_01457_ ), .B1(_01312_ ), .B2(_04754_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ) );
AND4_X1 _17385_ ( .A1(\io_master_arid [1] ), .A2(_00577_ ), .A3(_00579_ ), .A4(_01320_ ), .ZN(_01458_ ) );
OAI21_X1 _17386_ ( .A(_01329_ ), .B1(_01330_ ), .B2(_01458_ ), .ZN(_01459_ ) );
AOI22_X1 _17387_ ( .A1(_01308_ ), .A2(_01459_ ), .B1(_01312_ ), .B2(_04731_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ) );
NOR3_X1 _17388_ ( .A1(_00582_ ), .A2(_06027_ ), .A3(_01278_ ), .ZN(_01460_ ) );
OAI21_X1 _17389_ ( .A(_01329_ ), .B1(_01330_ ), .B2(_01460_ ), .ZN(_01461_ ) );
NAND2_X1 _17390_ ( .A1(_01313_ ), .A2(_01461_ ), .ZN(_01462_ ) );
MUX2_X1 _17391_ ( .A(\EX_LS_result_reg [23] ), .B(_01462_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ) );
NOR3_X1 _17392_ ( .A1(_00585_ ), .A2(_06027_ ), .A3(_01278_ ), .ZN(_01463_ ) );
OAI21_X1 _17393_ ( .A(_01329_ ), .B1(_01330_ ), .B2(_01463_ ), .ZN(_01464_ ) );
AOI22_X1 _17394_ ( .A1(_01308_ ), .A2(_01464_ ), .B1(_01312_ ), .B2(_04539_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ) );
NOR3_X1 _17395_ ( .A1(_00484_ ), .A2(_06027_ ), .A3(_01278_ ), .ZN(_01465_ ) );
OAI21_X1 _17396_ ( .A(_01329_ ), .B1(_01330_ ), .B2(_01465_ ), .ZN(_01466_ ) );
NAND2_X1 _17397_ ( .A1(_01313_ ), .A2(_01466_ ), .ZN(_01467_ ) );
MUX2_X1 _17398_ ( .A(\EX_LS_result_reg [31] ), .B(_01467_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17399_ ( .A1(\LS_WB_waddr_reg [1] ), .A2(\LS_WB_waddr_reg [0] ), .ZN(_01468_ ) );
INV_X1 _17400_ ( .A(\LS_WB_waddr_reg [3] ), .ZN(_01469_ ) );
INV_X1 _17401_ ( .A(\LS_WB_waddr_reg [2] ), .ZN(_01470_ ) );
NAND3_X1 _17402_ ( .A1(_01468_ ), .A2(_01469_ ), .A3(_01470_ ), .ZN(_01471_ ) );
AND2_X1 _17403_ ( .A1(_01547_ ), .A2(LS_WB_wen_reg ), .ZN(_01472_ ) );
NAND2_X1 _17404_ ( .A1(_01471_ ), .A2(_01472_ ), .ZN(_01473_ ) );
BUF_X4 _17405_ ( .A(_01473_ ), .Z(_01474_ ) );
INV_X1 _17406_ ( .A(\LS_WB_waddr_reg [1] ), .ZN(_01475_ ) );
INV_X1 _17407_ ( .A(\LS_WB_waddr_reg [0] ), .ZN(_01476_ ) );
AOI21_X1 _17408_ ( .A(_01474_ ), .B1(_01475_ ), .B2(_01476_ ), .ZN(_01477_ ) );
NOR2_X1 _17409_ ( .A1(_01473_ ), .A2(_01469_ ), .ZN(_01478_ ) );
NOR4_X1 _17410_ ( .A1(_01477_ ), .A2(_01478_ ), .A3(_01470_ ), .A4(_01474_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ) );
NOR2_X1 _17411_ ( .A1(_01474_ ), .A2(_01470_ ), .ZN(_01479_ ) );
NOR2_X1 _17412_ ( .A1(_01474_ ), .A2(_01476_ ), .ZN(_01480_ ) );
AND4_X1 _17413_ ( .A1(_01469_ ), .A2(_01479_ ), .A3(_01480_ ), .A4(_01475_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ) );
AND4_X1 _17414_ ( .A1(_01470_ ), .A2(_01478_ ), .A3(_01480_ ), .A4(_01475_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ) );
NOR2_X1 _17415_ ( .A1(_01473_ ), .A2(_01475_ ), .ZN(_01481_ ) );
AND4_X1 _17416_ ( .A1(_01470_ ), .A2(_01478_ ), .A3(_01481_ ), .A4(_01476_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ) );
CLKBUF_X1 _17417_ ( .A(reset ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ) );
AOI21_X1 _17418_ ( .A(_01474_ ), .B1(_01469_ ), .B2(_01470_ ), .ZN(_01482_ ) );
NOR4_X1 _17419_ ( .A1(_01482_ ), .A2(_01481_ ), .A3(_01476_ ), .A4(_01474_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ) );
NOR4_X1 _17420_ ( .A1(_01482_ ), .A2(_01480_ ), .A3(_01475_ ), .A4(_01474_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ) );
AND4_X1 _17421_ ( .A1(_01469_ ), .A2(_01479_ ), .A3(_01481_ ), .A4(_01476_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _17422_ ( .A1(_01469_ ), .A2(_01479_ ), .A3(_01481_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ) );
NOR4_X1 _17423_ ( .A1(_01477_ ), .A2(_01479_ ), .A3(_01469_ ), .A4(_01474_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ) );
NOR4_X1 _17424_ ( .A1(_01477_ ), .A2(_01469_ ), .A3(_01470_ ), .A4(_01474_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ) );
AND4_X1 _17425_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01478_ ), .A3(_01480_ ), .A4(_01475_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17426_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01478_ ), .A3(_01481_ ), .A4(_01476_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ) );
AND4_X1 _17427_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01478_ ), .A3(_01480_ ), .A4(\LS_WB_waddr_reg [1] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ) );
AND4_X1 _17428_ ( .A1(_01470_ ), .A2(_01478_ ), .A3(_01481_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ) );
NOR4_X1 _17429_ ( .A1(_01482_ ), .A2(_01475_ ), .A3(_01476_ ), .A4(_01474_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ) );
NAND3_X1 _17430_ ( .A1(_01949_ ), .A2(_01618_ ), .A3(_01956_ ), .ZN(_01483_ ) );
NAND2_X1 _17431_ ( .A1(_01483_ ), .A2(_01618_ ), .ZN(\myminixbar.state_$_DFF_P__Q_1_D ) );
AOI211_X1 _17432_ ( .A(reset ), .B(_01949_ ), .C1(_01950_ ), .C2(_06039_ ), .ZN(\myminixbar.state_$_DFF_P__Q_D ) );
CLKBUF_X2 _17433_ ( .A(_01471_ ), .Z(_01484_ ) );
CLKBUF_X2 _17434_ ( .A(_01472_ ), .Z(_01485_ ) );
AND3_X1 _17435_ ( .A1(_01484_ ), .A2(\LS_WB_wdata_reg [21] ), .A3(_01485_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ) );
AND3_X1 _17436_ ( .A1(_01484_ ), .A2(\LS_WB_wdata_reg [20] ), .A3(_01485_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ) );
AND3_X1 _17437_ ( .A1(_01484_ ), .A2(\LS_WB_wdata_reg [19] ), .A3(_01485_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ) );
AND3_X1 _17438_ ( .A1(_01484_ ), .A2(\LS_WB_wdata_reg [18] ), .A3(_01485_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ) );
AND3_X1 _17439_ ( .A1(_01484_ ), .A2(\LS_WB_wdata_reg [17] ), .A3(_01485_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ) );
AND3_X1 _17440_ ( .A1(_01484_ ), .A2(\LS_WB_wdata_reg [16] ), .A3(_01485_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ) );
AND3_X1 _17441_ ( .A1(_01484_ ), .A2(\LS_WB_wdata_reg [15] ), .A3(_01485_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ) );
AND3_X1 _17442_ ( .A1(_01484_ ), .A2(\LS_WB_wdata_reg [14] ), .A3(_01485_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ) );
AND3_X1 _17443_ ( .A1(_01484_ ), .A2(\LS_WB_wdata_reg [13] ), .A3(_01485_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ) );
AND3_X1 _17444_ ( .A1(_01484_ ), .A2(\LS_WB_wdata_reg [12] ), .A3(_01485_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ) );
CLKBUF_X2 _17445_ ( .A(_01471_ ), .Z(_01486_ ) );
CLKBUF_X2 _17446_ ( .A(_01472_ ), .Z(_01487_ ) );
AND3_X1 _17447_ ( .A1(_01486_ ), .A2(\LS_WB_wdata_reg [30] ), .A3(_01487_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ) );
AND3_X1 _17448_ ( .A1(_01486_ ), .A2(\LS_WB_wdata_reg [11] ), .A3(_01487_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ) );
AND3_X1 _17449_ ( .A1(_01486_ ), .A2(\LS_WB_wdata_reg [10] ), .A3(_01487_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ) );
AND3_X1 _17450_ ( .A1(_01486_ ), .A2(\LS_WB_wdata_reg [9] ), .A3(_01487_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ) );
AND3_X1 _17451_ ( .A1(_01486_ ), .A2(\LS_WB_wdata_reg [8] ), .A3(_01487_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ) );
AND3_X1 _17452_ ( .A1(_01486_ ), .A2(\LS_WB_wdata_reg [7] ), .A3(_01487_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ) );
AND3_X1 _17453_ ( .A1(_01486_ ), .A2(\LS_WB_wdata_reg [6] ), .A3(_01487_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ) );
AND3_X1 _17454_ ( .A1(_01486_ ), .A2(\LS_WB_wdata_reg [5] ), .A3(_01487_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ) );
AND3_X1 _17455_ ( .A1(_01486_ ), .A2(\LS_WB_wdata_reg [4] ), .A3(_01487_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ) );
AND3_X1 _17456_ ( .A1(_01486_ ), .A2(\LS_WB_wdata_reg [3] ), .A3(_01487_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ) );
CLKBUF_X2 _17457_ ( .A(_01471_ ), .Z(_01488_ ) );
CLKBUF_X2 _17458_ ( .A(_01472_ ), .Z(_01489_ ) );
AND3_X1 _17459_ ( .A1(_01488_ ), .A2(\LS_WB_wdata_reg [2] ), .A3(_01489_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ) );
AND3_X1 _17460_ ( .A1(_01488_ ), .A2(\LS_WB_wdata_reg [29] ), .A3(_01489_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ) );
AND3_X1 _17461_ ( .A1(_01488_ ), .A2(\LS_WB_wdata_reg [1] ), .A3(_01489_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ) );
AND3_X1 _17462_ ( .A1(_01488_ ), .A2(\LS_WB_wdata_reg [0] ), .A3(_01489_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ) );
AND3_X1 _17463_ ( .A1(_01488_ ), .A2(\LS_WB_wdata_reg [28] ), .A3(_01489_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ) );
AND3_X1 _17464_ ( .A1(_01488_ ), .A2(\LS_WB_wdata_reg [27] ), .A3(_01489_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ) );
AND3_X1 _17465_ ( .A1(_01488_ ), .A2(\LS_WB_wdata_reg [26] ), .A3(_01489_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ) );
AND3_X1 _17466_ ( .A1(_01488_ ), .A2(\LS_WB_wdata_reg [25] ), .A3(_01489_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ) );
AND3_X1 _17467_ ( .A1(_01488_ ), .A2(\LS_WB_wdata_reg [24] ), .A3(_01489_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ) );
AND3_X1 _17468_ ( .A1(_01488_ ), .A2(\LS_WB_wdata_reg [23] ), .A3(_01489_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ) );
AND3_X1 _17469_ ( .A1(_01471_ ), .A2(\LS_WB_wdata_reg [22] ), .A3(_01472_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17470_ ( .A1(_01471_ ), .A2(\LS_WB_wdata_reg [31] ), .A3(_01472_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_D ) );
AND3_X1 _17471_ ( .A1(_01618_ ), .A2(\mysc.state [2] ), .A3(\mylsu.previous_load_done ), .ZN(\mysc.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _17472_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01490_ ) );
AND2_X1 _17473_ ( .A1(_01490_ ), .A2(\myidu.stall_quest_loaduse ), .ZN(_01491_ ) );
INV_X1 _17474_ ( .A(_01491_ ), .ZN(_01492_ ) );
NOR2_X1 _17475_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01493_ ) );
OAI211_X1 _17476_ ( .A(_01547_ ), .B(\mysc.state [0] ), .C1(_01492_ ), .C2(_01493_ ), .ZN(_01494_ ) );
INV_X1 _17477_ ( .A(_01494_ ), .ZN(_01495_ ) );
OR3_X1 _17478_ ( .A1(_01495_ ), .A2(reset ), .A3(\mysc.state [1] ), .ZN(\mysc.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _17479_ ( .A1(_01492_ ), .A2(reset ), .A3(_01493_ ), .ZN(_01496_ ) );
NAND2_X1 _17480_ ( .A1(_01496_ ), .A2(\mysc.state [0] ), .ZN(_01497_ ) );
OR3_X1 _17481_ ( .A1(_03871_ ), .A2(reset ), .A3(\mylsu.previous_load_done ), .ZN(_01498_ ) );
NAND2_X1 _17482_ ( .A1(_01497_ ), .A2(_01498_ ), .ZN(\mysc.state_$_DFF_P__Q_D ) );
CLKGATE_X1 _17483_ ( .CK(clock ), .E(\mylsu.previous_load_done ), .GCK(_07973_ ) );
CLKGATE_X1 _17484_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ), .GCK(_07974_ ) );
CLKGATE_X1 _17485_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ), .GCK(_07975_ ) );
CLKGATE_X1 _17486_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ), .GCK(_07976_ ) );
CLKGATE_X1 _17487_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ), .GCK(_07977_ ) );
CLKGATE_X1 _17488_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ), .GCK(_07978_ ) );
CLKGATE_X1 _17489_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ), .GCK(_07979_ ) );
CLKGATE_X1 _17490_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ), .GCK(_07980_ ) );
CLKGATE_X1 _17491_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ), .GCK(_07981_ ) );
CLKGATE_X1 _17492_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ), .GCK(_07982_ ) );
CLKGATE_X1 _17493_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ), .GCK(_07983_ ) );
CLKGATE_X1 _17494_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ), .GCK(_07984_ ) );
CLKGATE_X1 _17495_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ), .GCK(_07985_ ) );
CLKGATE_X1 _17496_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ), .GCK(_07986_ ) );
CLKGATE_X1 _17497_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ), .GCK(_07987_ ) );
CLKGATE_X1 _17498_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ), .GCK(_07988_ ) );
CLKGATE_X1 _17499_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ), .GCK(_07989_ ) );
CLKGATE_X1 _17500_ ( .CK(clock ), .E(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_07990_ ) );
CLKGATE_X1 _17501_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ), .GCK(_07991_ ) );
CLKGATE_X1 _17502_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ), .GCK(_07992_ ) );
CLKGATE_X1 _17503_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .GCK(_07993_ ) );
CLKGATE_X1 _17504_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_07994_ ) );
CLKGATE_X1 _17505_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .GCK(_07995_ ) );
CLKGATE_X1 _17506_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E ), .GCK(_07996_ ) );
CLKGATE_X1 _17507_ ( .CK(clock ), .E(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .GCK(_07997_ ) );
CLKGATE_X1 _17508_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP1P__Q_E ), .GCK(_07998_ ) );
CLKGATE_X1 _17509_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_07999_ ) );
CLKGATE_X1 _17510_ ( .CK(clock ), .E(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_08000_ ) );
CLKGATE_X1 _17511_ ( .CK(clock ), .E(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_08001_ ) );
CLKGATE_X1 _17512_ ( .CK(clock ), .E(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_08002_ ) );
CLKGATE_X1 _17513_ ( .CK(clock ), .E(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_08003_ ) );
CLKGATE_X1 _17514_ ( .CK(clock ), .E(\myifu.myicache.tag[3]_$_DFFE_PP__Q_E ), .GCK(_08004_ ) );
CLKGATE_X1 _17515_ ( .CK(clock ), .E(\myifu.myicache.tag[2]_$_DFFE_PP__Q_E ), .GCK(_08005_ ) );
CLKGATE_X1 _17516_ ( .CK(clock ), .E(\myifu.myicache.tag[1]_$_DFFE_PP__Q_E ), .GCK(_08006_ ) );
CLKGATE_X1 _17517_ ( .CK(clock ), .E(\myifu.myicache.tag[0]_$_DFFE_PP__Q_E ), .GCK(_08007_ ) );
CLKGATE_X1 _17518_ ( .CK(clock ), .E(\myifu.myicache.data[7]_$_DFFE_PP__Q_E ), .GCK(_08008_ ) );
CLKGATE_X1 _17519_ ( .CK(clock ), .E(\myifu.myicache.data[6]_$_DFFE_PP__Q_E ), .GCK(_08009_ ) );
CLKGATE_X1 _17520_ ( .CK(clock ), .E(\myifu.myicache.data[5]_$_DFFE_PP__Q_E ), .GCK(_08010_ ) );
CLKGATE_X1 _17521_ ( .CK(clock ), .E(\myifu.myicache.data[4]_$_DFFE_PP__Q_E ), .GCK(_08011_ ) );
CLKGATE_X1 _17522_ ( .CK(clock ), .E(\myifu.myicache.data[3]_$_DFFE_PP__Q_E ), .GCK(_08012_ ) );
CLKGATE_X1 _17523_ ( .CK(clock ), .E(\myifu.myicache.data[2]_$_DFFE_PP__Q_E ), .GCK(_08013_ ) );
CLKGATE_X1 _17524_ ( .CK(clock ), .E(\myifu.myicache.data[1]_$_DFFE_PP__Q_E ), .GCK(_08014_ ) );
CLKGATE_X1 _17525_ ( .CK(clock ), .E(\myifu.myicache.data[0]_$_DFFE_PP__Q_E ), .GCK(_08015_ ) );
CLKGATE_X1 _17526_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08016_ ) );
CLKGATE_X1 _17527_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E ), .GCK(_08017_ ) );
CLKGATE_X1 _17528_ ( .CK(clock ), .E(\myidu.typ_$_SDFFE_PP0P__Q_E ), .GCK(_08018_ ) );
CLKGATE_X1 _17529_ ( .CK(clock ), .E(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ), .GCK(_08019_ ) );
CLKGATE_X1 _17530_ ( .CK(clock ), .E(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .GCK(_08020_ ) );
CLKGATE_X1 _17531_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08021_ ) );
CLKGATE_X1 _17532_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08022_ ) );
CLKGATE_X1 _17533_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08023_ ) );
CLKGATE_X1 _17534_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ), .GCK(_08024_ ) );
CLKGATE_X1 _17535_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08025_ ) );
CLKGATE_X1 _17536_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ), .GCK(_08026_ ) );
CLKGATE_X1 _17537_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ), .GCK(_08027_ ) );
CLKGATE_X1 _17538_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ), .GCK(_08028_ ) );
CLKGATE_X1 _17539_ ( .CK(clock ), .E(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08029_ ) );
CLKGATE_X1 _17540_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y ), .GCK(_08030_ ) );
CLKGATE_X1 _17541_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ), .GCK(_08031_ ) );
CLKGATE_X1 _17542_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E ), .GCK(_08032_ ) );
CLKGATE_X1 _17543_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08033_ ) );
CLKGATE_X1 _17544_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__B_Y_$_ORNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08034_ ) );
CLKGATE_X1 _17545_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ), .GCK(_08035_ ) );
CLKGATE_X1 _17546_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ), .GCK(_08036_ ) );
CLKGATE_X1 _17547_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08037_ ) );
LOGIC1_X1 _17548_ ( .Z(\io_master_awid [0] ) );
LOGIC0_X1 _17549_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q ( .D(_00000_ ), .CK(clock ), .Q(\myclint.mtime [63] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_1 ( .D(_00001_ ), .CK(clock ), .Q(\myclint.mtime [62] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_10 ( .D(_00002_ ), .CK(clock ), .Q(\myclint.mtime [53] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_11 ( .D(_00003_ ), .CK(clock ), .Q(\myclint.mtime [52] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_12 ( .D(_00004_ ), .CK(clock ), .Q(\myclint.mtime [51] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_13 ( .D(_00005_ ), .CK(clock ), .Q(\myclint.mtime [50] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_14 ( .D(_00006_ ), .CK(clock ), .Q(\myclint.mtime [49] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_15 ( .D(_00007_ ), .CK(clock ), .Q(\myclint.mtime [48] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_16 ( .D(_00008_ ), .CK(clock ), .Q(\myclint.mtime [47] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_17 ( .D(_00009_ ), .CK(clock ), .Q(\myclint.mtime [46] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_18 ( .D(_00010_ ), .CK(clock ), .Q(\myclint.mtime [45] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_19 ( .D(_00011_ ), .CK(clock ), .Q(\myclint.mtime [44] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_2 ( .D(_00012_ ), .CK(clock ), .Q(\myclint.mtime [61] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_20 ( .D(_00013_ ), .CK(clock ), .Q(\myclint.mtime [43] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_21 ( .D(_00014_ ), .CK(clock ), .Q(\myclint.mtime [42] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_22 ( .D(_00015_ ), .CK(clock ), .Q(\myclint.mtime [41] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_23 ( .D(_00016_ ), .CK(clock ), .Q(\myclint.mtime [40] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_24 ( .D(_00017_ ), .CK(clock ), .Q(\myclint.mtime [39] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_25 ( .D(_00018_ ), .CK(clock ), .Q(\myclint.mtime [38] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_26 ( .D(_00019_ ), .CK(clock ), .Q(\myclint.mtime [37] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_27 ( .D(_00020_ ), .CK(clock ), .Q(\myclint.mtime [36] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_28 ( .D(_00021_ ), .CK(clock ), .Q(\myclint.mtime [35] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_29 ( .D(_00022_ ), .CK(clock ), .Q(\myclint.mtime [34] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_3 ( .D(_00023_ ), .CK(clock ), .Q(\myclint.mtime [60] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_30 ( .D(_00024_ ), .CK(clock ), .Q(\myclint.mtime [33] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_31 ( .D(_00025_ ), .CK(clock ), .Q(\myclint.mtime [32] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_32 ( .D(_00026_ ), .CK(clock ), .Q(\myclint.mtime [31] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_33 ( .D(_00027_ ), .CK(clock ), .Q(\myclint.mtime [30] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_34 ( .D(_00028_ ), .CK(clock ), .Q(\myclint.mtime [29] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_35 ( .D(_00029_ ), .CK(clock ), .Q(\myclint.mtime [28] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_36 ( .D(_00030_ ), .CK(clock ), .Q(\myclint.mtime [27] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_37 ( .D(_00031_ ), .CK(clock ), .Q(\myclint.mtime [26] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_38 ( .D(_00032_ ), .CK(clock ), .Q(\myclint.mtime [25] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_39 ( .D(_00033_ ), .CK(clock ), .Q(\myclint.mtime [24] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_4 ( .D(_00034_ ), .CK(clock ), .Q(\myclint.mtime [59] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_40 ( .D(_00035_ ), .CK(clock ), .Q(\myclint.mtime [23] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_41 ( .D(_00036_ ), .CK(clock ), .Q(\myclint.mtime [22] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_42 ( .D(_00037_ ), .CK(clock ), .Q(\myclint.mtime [21] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_43 ( .D(_00038_ ), .CK(clock ), .Q(\myclint.mtime [20] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_44 ( .D(_00039_ ), .CK(clock ), .Q(\myclint.mtime [19] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_45 ( .D(_00040_ ), .CK(clock ), .Q(\myclint.mtime [18] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_46 ( .D(_00041_ ), .CK(clock ), .Q(\myclint.mtime [17] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_47 ( .D(_00042_ ), .CK(clock ), .Q(\myclint.mtime [16] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_48 ( .D(_00043_ ), .CK(clock ), .Q(\myclint.mtime [15] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_49 ( .D(_00044_ ), .CK(clock ), .Q(\myclint.mtime [14] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_5 ( .D(_00045_ ), .CK(clock ), .Q(\myclint.mtime [58] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_50 ( .D(_00046_ ), .CK(clock ), .Q(\myclint.mtime [13] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_51 ( .D(_00047_ ), .CK(clock ), .Q(\myclint.mtime [12] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_52 ( .D(_00048_ ), .CK(clock ), .Q(\myclint.mtime [11] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_53 ( .D(_00049_ ), .CK(clock ), .Q(\myclint.mtime [10] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_54 ( .D(_00050_ ), .CK(clock ), .Q(\myclint.mtime [9] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_55 ( .D(_00051_ ), .CK(clock ), .Q(\myclint.mtime [8] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_56 ( .D(_00052_ ), .CK(clock ), .Q(\myclint.mtime [7] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_57 ( .D(_00053_ ), .CK(clock ), .Q(\myclint.mtime [6] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_58 ( .D(_00054_ ), .CK(clock ), .Q(\myclint.mtime [5] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_59 ( .D(_00055_ ), .CK(clock ), .Q(\myclint.mtime [4] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_6 ( .D(_00056_ ), .CK(clock ), .Q(\myclint.mtime [57] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_60 ( .D(_00057_ ), .CK(clock ), .Q(\myclint.mtime [3] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_61 ( .D(_00058_ ), .CK(clock ), .Q(\myclint.mtime [2] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_62 ( .D(_00059_ ), .CK(clock ), .Q(\myclint.mtime [1] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_63 ( .D(_00060_ ), .CK(clock ), .Q(\myclint.mtime [0] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_7 ( .D(_00061_ ), .CK(clock ), .Q(\myclint.mtime [56] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_8 ( .D(_00062_ ), .CK(clock ), .Q(\myclint.mtime [55] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_9 ( .D(_00063_ ), .CK(clock ), .Q(\myclint.mtime [54] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.state_r_$_SDFF_PP0__Q ( .D(_00064_ ), .CK(clock ), .Q(\myclint.rvalid ), .QN(\myclint.state_r_$_NOT__A_Y ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][31] ), .QN(_08268_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][30] ), .QN(_08269_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][21] ), .QN(_08270_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][20] ), .QN(_08271_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][19] ), .QN(_08272_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][18] ), .QN(_08273_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][17] ), .QN(_08274_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][16] ), .QN(_08275_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][15] ), .QN(_08276_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][14] ), .QN(_08277_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][13] ), .QN(_08278_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][12] ), .QN(_08279_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][29] ), .QN(_08280_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][11] ), .QN(_08281_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][10] ), .QN(_08282_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][9] ), .QN(_08283_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][8] ), .QN(_08284_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][7] ), .QN(_08285_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][6] ), .QN(_08286_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][5] ), .QN(_08287_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][4] ), .QN(_08288_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][3] ), .QN(_08289_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][2] ), .QN(_08290_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][28] ), .QN(_08291_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][1] ), .QN(_08292_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][0] ), .QN(_08293_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][27] ), .QN(_08294_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][26] ), .QN(_08295_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][25] ), .QN(_08296_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][24] ), .QN(_08297_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][23] ), .QN(_08298_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08037_ ), .Q(\mycsreg.CSReg[0][22] ), .QN(_08299_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08036_ ), .Q(\mtvec [31] ), .QN(_08300_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08036_ ), .Q(\mtvec [30] ), .QN(_08301_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08036_ ), .Q(\mtvec [21] ), .QN(_08302_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08036_ ), .Q(\mtvec [20] ), .QN(_08303_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08036_ ), .Q(\mtvec [19] ), .QN(_08304_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08036_ ), .Q(\mtvec [18] ), .QN(_08305_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08036_ ), .Q(\mtvec [17] ), .QN(_08306_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08036_ ), .Q(\mtvec [16] ), .QN(_08307_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08036_ ), .Q(\mtvec [15] ), .QN(_08308_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08036_ ), .Q(\mtvec [14] ), .QN(_08309_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08036_ ), .Q(\mtvec [13] ), .QN(_08310_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08036_ ), .Q(\mtvec [12] ), .QN(_08311_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08036_ ), .Q(\mtvec [29] ), .QN(_08312_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08036_ ), .Q(\mtvec [11] ), .QN(_08313_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08036_ ), .Q(\mtvec [10] ), .QN(_08314_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08036_ ), .Q(\mtvec [9] ), .QN(_08315_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08036_ ), .Q(\mtvec [8] ), .QN(_08316_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08036_ ), .Q(\mtvec [7] ), .QN(_08317_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08036_ ), .Q(\mtvec [6] ), .QN(_08318_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08036_ ), .Q(\mtvec [5] ), .QN(_08319_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08036_ ), .Q(\mtvec [4] ), .QN(_08320_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08036_ ), .Q(\mtvec [3] ), .QN(_08321_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08036_ ), .Q(\mtvec [2] ), .QN(_08322_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08036_ ), .Q(\mtvec [28] ), .QN(_08323_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08036_ ), .Q(\mtvec [1] ), .QN(_08324_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08036_ ), .Q(\mtvec [0] ), .QN(_08325_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08036_ ), .Q(\mtvec [27] ), .QN(_08326_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08036_ ), .Q(\mtvec [26] ), .QN(_08327_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08036_ ), .Q(\mtvec [25] ), .QN(_08328_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08036_ ), .Q(\mtvec [24] ), .QN(_08329_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08036_ ), .Q(\mtvec [23] ), .QN(_08330_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08036_ ), .Q(\mtvec [22] ), .QN(_08331_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08035_ ), .Q(\mepc [31] ), .QN(_08332_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08035_ ), .Q(\mepc [30] ), .QN(_08333_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08035_ ), .Q(\mepc [21] ), .QN(_08334_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08035_ ), .Q(\mepc [20] ), .QN(_08335_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08035_ ), .Q(\mepc [19] ), .QN(_08336_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08035_ ), .Q(\mepc [18] ), .QN(_08337_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08035_ ), .Q(\mepc [17] ), .QN(_08338_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08035_ ), .Q(\mepc [16] ), .QN(_08339_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08035_ ), .Q(\mepc [15] ), .QN(_08340_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08035_ ), .Q(\mepc [14] ), .QN(_08341_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08035_ ), .Q(\mepc [13] ), .QN(_08342_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08035_ ), .Q(\mepc [12] ), .QN(_08343_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08035_ ), .Q(\mepc [29] ), .QN(_08344_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08035_ ), .Q(\mepc [11] ), .QN(_08345_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08035_ ), .Q(\mepc [10] ), .QN(_08346_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08035_ ), .Q(\mepc [9] ), .QN(_08347_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08035_ ), .Q(\mepc [8] ), .QN(_08348_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08035_ ), .Q(\mepc [7] ), .QN(_08349_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08035_ ), .Q(\mepc [6] ), .QN(_08350_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08035_ ), .Q(\mepc [5] ), .QN(_08351_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08035_ ), .Q(\mepc [4] ), .QN(_08352_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08035_ ), .Q(\mepc [3] ), .QN(_08353_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08035_ ), .Q(\mepc [2] ), .QN(_08354_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08035_ ), .Q(\mepc [28] ), .QN(_08355_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08035_ ), .Q(\mepc [1] ), .QN(_08356_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08035_ ), .Q(\mepc [0] ), .QN(_08357_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08035_ ), .Q(\mepc [27] ), .QN(_08358_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08035_ ), .Q(\mepc [26] ), .QN(_08359_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08035_ ), .Q(\mepc [25] ), .QN(_08360_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08035_ ), .Q(\mepc [24] ), .QN(_08361_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08035_ ), .Q(\mepc [23] ), .QN(_08362_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08035_ ), .Q(\mepc [22] ), .QN(_08363_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][3] ), .QN(_08364_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_1 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][2] ), .QN(_08365_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_2 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][1] ), .QN(_08366_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_3 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][0] ), .QN(_08267_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q ( .D(_00065_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][31] ), .QN(_08266_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][30] ), .QN(_08265_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][21] ), .QN(_08264_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][20] ), .QN(_08263_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][19] ), .QN(_08262_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][18] ), .QN(_08261_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][17] ), .QN(_08260_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][16] ), .QN(_08259_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][15] ), .QN(_08258_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][14] ), .QN(_08257_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][13] ), .QN(_08256_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][12] ), .QN(_08255_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][29] ), .QN(_08254_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][11] ), .QN(_08253_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][10] ), .QN(_08252_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][9] ), .QN(_08251_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][8] ), .QN(_08250_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][7] ), .QN(_08249_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][6] ), .QN(_08248_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][5] ), .QN(_08247_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][4] ), .QN(_08246_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_3 ( .D(_00086_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][28] ), .QN(_08245_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_4 ( .D(_00087_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][27] ), .QN(_08244_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_5 ( .D(_00088_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][26] ), .QN(_08243_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_6 ( .D(_00089_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][25] ), .QN(_08242_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_7 ( .D(_00090_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][24] ), .QN(_08241_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_8 ( .D(_00091_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][23] ), .QN(_08240_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_9 ( .D(_00092_ ), .CK(_08034_ ), .Q(\mycsreg.CSReg[3][22] ), .QN(_08367_ ) );
DFF_X1 \mycsreg.excp_written_$_SDFF_PN0__Q ( .D(_00093_ ), .CK(clock ), .Q(excp_written ), .QN(_08368_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [31] ), .QN(_08239_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_1 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [30] ), .QN(_08369_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_10 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [21] ), .QN(_08370_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_11 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [20] ), .QN(_08371_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_12 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [19] ), .QN(_08372_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_13 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [18] ), .QN(_08373_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_14 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [17] ), .QN(_08374_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_15 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [16] ), .QN(_08375_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_16 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [15] ), .QN(_08376_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_17 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [14] ), .QN(_08377_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_18 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [13] ), .QN(_08378_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_19 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [12] ), .QN(_08379_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_2 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [29] ), .QN(_08380_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_20 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [11] ), .QN(_08381_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_21 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [10] ), .QN(_08382_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_22 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [9] ), .QN(_08383_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_23 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [8] ), .QN(_08384_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_24 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [7] ), .QN(_08385_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_25 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [6] ), .QN(_08386_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_26 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [5] ), .QN(_08387_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_27 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [4] ), .QN(_08388_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_28 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [3] ), .QN(_08389_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_29 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [2] ), .QN(_08390_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_3 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [28] ), .QN(_08391_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_30 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [1] ), .QN(_08392_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_31 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [0] ), .QN(_08393_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_4 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [27] ), .QN(_08394_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_5 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [26] ), .QN(_08395_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_6 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [25] ), .QN(_08396_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_7 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [24] ), .QN(_08397_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_8 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [23] ), .QN(_08398_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_9 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ), .CK(_08033_ ), .Q(\myec.mepc_tmp [22] ), .QN(_08238_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q ( .D(_00094_ ), .CK(_08032_ ), .Q(\myec.state [1] ), .QN(_08237_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q_1 ( .D(_00095_ ), .CK(_08032_ ), .Q(\myec.state [0] ), .QN(_08399_ ) );
DFF_X1 \myexu.check_quest_$_SDFF_PN0__Q ( .D(_00096_ ), .CK(clock ), .Q(check_quest ), .QN(_08400_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(_08236_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(_08401_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(_08402_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(_08403_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(_08404_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(_08405_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(_08406_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(_08407_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(_08408_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(_08409_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(_08410_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(_08235_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q ( .D(_00097_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(_08234_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_1 ( .D(_00098_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(_08233_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_10 ( .D(_00099_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(_08232_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_11 ( .D(_00100_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(_08231_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_12 ( .D(_00101_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(_08230_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_13 ( .D(_00102_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(_08229_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_14 ( .D(_00103_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(_08228_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_15 ( .D(_00104_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(_08227_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_16 ( .D(_00105_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(_08226_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_17 ( .D(_00106_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(_08225_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_18 ( .D(_00107_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(_08224_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_19 ( .D(_00108_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(_08223_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_2 ( .D(_00109_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(_08222_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_3 ( .D(_00110_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(_08221_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_4 ( .D(_00111_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(_08220_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_5 ( .D(_00112_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(_08219_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_6 ( .D(_00113_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(_08218_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_7 ( .D(_00114_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(_08217_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_8 ( .D(_00115_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(_08216_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_9 ( .D(_00116_ ), .CK(_08031_ ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(_08215_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q ( .D(_00117_ ), .CK(_08030_ ), .Q(\EX_LS_dest_reg [4] ), .QN(_08214_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_1 ( .D(_00118_ ), .CK(_08030_ ), .Q(\EX_LS_dest_reg [3] ), .QN(_08213_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_2 ( .D(_00119_ ), .CK(_08030_ ), .Q(\EX_LS_dest_reg [2] ), .QN(_08212_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_3 ( .D(_00120_ ), .CK(_08030_ ), .Q(\EX_LS_dest_reg [1] ), .QN(_08211_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_4 ( .D(_00121_ ), .CK(_08030_ ), .Q(\EX_LS_dest_reg [0] ), .QN(_08210_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q ( .D(_00122_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [30] ), .QN(_08209_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_1 ( .D(_00123_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [29] ), .QN(_08208_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_10 ( .D(_00124_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [20] ), .QN(_08207_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_11 ( .D(_00125_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [19] ), .QN(_08206_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_12 ( .D(_00126_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [18] ), .QN(_08205_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_13 ( .D(_00127_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [17] ), .QN(_08204_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_14 ( .D(_00128_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [16] ), .QN(_08203_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_15 ( .D(_00129_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [15] ), .QN(_08202_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_16 ( .D(_00130_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [14] ), .QN(_08201_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_17 ( .D(_00131_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [13] ), .QN(_08200_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_18 ( .D(_00132_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [12] ), .QN(_08199_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_19 ( .D(_00133_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [11] ), .QN(_08198_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_2 ( .D(_00134_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [28] ), .QN(_08197_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_20 ( .D(_00135_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [10] ), .QN(_08196_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_21 ( .D(_00136_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [9] ), .QN(_08195_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_22 ( .D(_00137_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [8] ), .QN(_08194_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_23 ( .D(_00138_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [7] ), .QN(_08193_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_24 ( .D(_00139_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [6] ), .QN(_08192_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_25 ( .D(_00140_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [5] ), .QN(_08191_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_26 ( .D(_00141_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [4] ), .QN(_08190_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_27 ( .D(_00142_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [3] ), .QN(_08189_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_28 ( .D(_00143_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [2] ), .QN(_08188_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_29 ( .D(_00144_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [1] ), .QN(_08187_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_3 ( .D(_00145_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [27] ), .QN(_08186_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_30 ( .D(_00146_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [0] ), .QN(_08185_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_4 ( .D(_00147_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [26] ), .QN(_08184_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_5 ( .D(_00148_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [25] ), .QN(_08183_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_6 ( .D(_00149_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [24] ), .QN(_08182_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_7 ( .D(_00150_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [23] ), .QN(_08181_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_8 ( .D(_00151_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [22] ), .QN(_08180_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_9 ( .D(_00152_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [21] ), .QN(_08179_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN1P__Q ( .D(_00153_ ), .CK(_08029_ ), .Q(\myexu.pc_jump [31] ), .QN(_08178_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q ( .D(_00154_ ), .CK(_08030_ ), .Q(\EX_LS_pc [31] ), .QN(_08177_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_1 ( .D(_00155_ ), .CK(_08030_ ), .Q(\EX_LS_pc [30] ), .QN(_08176_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_10 ( .D(_00156_ ), .CK(_08030_ ), .Q(\EX_LS_pc [21] ), .QN(_08175_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_11 ( .D(_00157_ ), .CK(_08030_ ), .Q(\EX_LS_pc [20] ), .QN(_08174_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_12 ( .D(_00158_ ), .CK(_08030_ ), .Q(\EX_LS_pc [19] ), .QN(_08173_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_13 ( .D(_00159_ ), .CK(_08030_ ), .Q(\EX_LS_pc [18] ), .QN(_08172_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_14 ( .D(_00160_ ), .CK(_08030_ ), .Q(\EX_LS_pc [17] ), .QN(_08171_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_15 ( .D(_00161_ ), .CK(_08030_ ), .Q(\EX_LS_pc [16] ), .QN(_08170_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_16 ( .D(_00162_ ), .CK(_08030_ ), .Q(\EX_LS_pc [15] ), .QN(_08169_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_17 ( .D(_00163_ ), .CK(_08030_ ), .Q(\EX_LS_pc [14] ), .QN(_08168_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_18 ( .D(_00164_ ), .CK(_08030_ ), .Q(\EX_LS_pc [13] ), .QN(_08167_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_19 ( .D(_00165_ ), .CK(_08030_ ), .Q(\EX_LS_pc [12] ), .QN(_08166_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_2 ( .D(_00166_ ), .CK(_08030_ ), .Q(\EX_LS_pc [29] ), .QN(_08165_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_20 ( .D(_00167_ ), .CK(_08030_ ), .Q(\EX_LS_pc [11] ), .QN(_08164_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_21 ( .D(_00168_ ), .CK(_08030_ ), .Q(\EX_LS_pc [10] ), .QN(_08163_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_22 ( .D(_00169_ ), .CK(_08030_ ), .Q(\EX_LS_pc [9] ), .QN(_08162_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_23 ( .D(_00170_ ), .CK(_08030_ ), .Q(\EX_LS_pc [8] ), .QN(_08161_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_24 ( .D(_00171_ ), .CK(_08030_ ), .Q(\EX_LS_pc [7] ), .QN(_08160_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_25 ( .D(_00172_ ), .CK(_08030_ ), .Q(\EX_LS_pc [6] ), .QN(_08159_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_26 ( .D(_00173_ ), .CK(_08030_ ), .Q(\EX_LS_pc [5] ), .QN(_08158_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_27 ( .D(_00174_ ), .CK(_08030_ ), .Q(\EX_LS_pc [4] ), .QN(_08157_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_28 ( .D(_00175_ ), .CK(_08030_ ), .Q(\EX_LS_pc [3] ), .QN(_08156_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_29 ( .D(_00176_ ), .CK(_08030_ ), .Q(\EX_LS_pc [2] ), .QN(_08155_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_3 ( .D(_00177_ ), .CK(_08030_ ), .Q(\EX_LS_pc [28] ), .QN(_08154_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_30 ( .D(_00178_ ), .CK(_08030_ ), .Q(\EX_LS_pc [1] ), .QN(_08153_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_31 ( .D(_00179_ ), .CK(_08030_ ), .Q(\EX_LS_pc [0] ), .QN(_08152_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_4 ( .D(_00180_ ), .CK(_08030_ ), .Q(\EX_LS_pc [27] ), .QN(_08151_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_5 ( .D(_00181_ ), .CK(_08030_ ), .Q(\EX_LS_pc [26] ), .QN(_08150_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_6 ( .D(_00182_ ), .CK(_08030_ ), .Q(\EX_LS_pc [25] ), .QN(_08149_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_7 ( .D(_00183_ ), .CK(_08030_ ), .Q(\EX_LS_pc [24] ), .QN(_08148_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_8 ( .D(_00184_ ), .CK(_08030_ ), .Q(\EX_LS_pc [23] ), .QN(_08147_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_9 ( .D(_00185_ ), .CK(_08030_ ), .Q(\EX_LS_pc [22] ), .QN(_08411_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(_08412_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(_08413_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(_08414_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(_08415_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_12 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(_08416_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_13 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(_08417_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_14 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(_08418_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_15 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(_08419_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_16 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(_08420_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_17 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(_08421_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_18 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(_08422_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_19 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(_08423_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(_08424_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_20 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(_08425_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_21 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(_08426_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_22 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(_08427_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_23 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(_08428_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_24 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(_08429_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_25 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(_08430_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_26 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(_08431_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_27 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(_08432_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_28 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(_08433_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_29 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(_08434_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(_08435_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_30 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(_08436_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_31 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(_08437_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(_08438_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(_08439_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(_08440_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(_08441_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(_08442_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08031_ ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(_08443_ ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q ( .D(\myexu.result_reg_$_DFFE_PP__Q_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_1 ( .D(\myexu.result_reg_$_DFFE_PP__Q_1_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_10 ( .D(\myexu.result_reg_$_DFFE_PP__Q_10_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_11 ( .D(\myexu.result_reg_$_DFFE_PP__Q_11_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_12 ( .D(\myexu.result_reg_$_DFFE_PP__Q_12_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_13 ( .D(\myexu.result_reg_$_DFFE_PP__Q_13_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_14 ( .D(\myexu.result_reg_$_DFFE_PP__Q_14_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_15 ( .D(\myexu.result_reg_$_DFFE_PP__Q_15_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_16 ( .D(\myexu.result_reg_$_DFFE_PP__Q_16_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_17 ( .D(\myexu.result_reg_$_DFFE_PP__Q_17_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_18 ( .D(\myexu.result_reg_$_DFFE_PP__Q_18_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_19 ( .D(\myexu.result_reg_$_DFFE_PP__Q_19_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_2 ( .D(\myexu.result_reg_$_DFFE_PP__Q_2_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_20 ( .D(\myexu.result_reg_$_DFFE_PP__Q_20_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_21 ( .D(\myexu.result_reg_$_DFFE_PP__Q_21_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_22 ( .D(\myexu.result_reg_$_DFFE_PP__Q_22_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_23 ( .D(\myexu.result_reg_$_DFFE_PP__Q_23_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_24 ( .D(\myexu.result_reg_$_DFFE_PP__Q_24_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_25 ( .D(\myexu.result_reg_$_DFFE_PP__Q_25_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_26 ( .D(\myexu.result_reg_$_DFFE_PP__Q_26_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_27 ( .D(\myexu.result_reg_$_DFFE_PP__Q_27_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_28 ( .D(\myexu.result_reg_$_DFFE_PP__Q_28_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_29 ( .D(\myexu.result_reg_$_DFFE_PP__Q_29_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_3 ( .D(\myexu.result_reg_$_DFFE_PP__Q_3_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_30 ( .D(\myexu.result_reg_$_DFFE_PP__Q_30_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_31 ( .D(\myexu.result_reg_$_DFFE_PP__Q_31_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_4 ( .D(\myexu.result_reg_$_DFFE_PP__Q_4_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_5 ( .D(\myexu.result_reg_$_DFFE_PP__Q_5_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_6 ( .D(\myexu.result_reg_$_DFFE_PP__Q_6_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_7 ( .D(\myexu.result_reg_$_DFFE_PP__Q_7_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_8 ( .D(\myexu.result_reg_$_DFFE_PP__Q_8_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_9 ( .D(\myexu.result_reg_$_DFFE_PP__Q_9_D ), .CK(_08031_ ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.state_$_SDFF_PN0__Q ( .D(_00187_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q ( .D(_00186_ ), .CK(_08030_ ), .Q(\EX_LS_flag [2] ), .QN(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_1 ( .D(_00188_ ), .CK(_08030_ ), .Q(\EX_LS_flag [1] ), .QN(_08146_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_2 ( .D(_00189_ ), .CK(_08030_ ), .Q(\EX_LS_flag [0] ), .QN(_08145_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_3 ( .D(_00190_ ), .CK(_08030_ ), .Q(\EX_LS_typ [4] ), .QN(_08144_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_4 ( .D(_00191_ ), .CK(_08030_ ), .Q(\EX_LS_typ [3] ), .QN(_08143_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_5 ( .D(_00192_ ), .CK(_08030_ ), .Q(\EX_LS_typ [2] ), .QN(_08142_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_6 ( .D(_00193_ ), .CK(_08030_ ), .Q(\EX_LS_typ [1] ), .QN(_08141_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_7 ( .D(_00194_ ), .CK(_08030_ ), .Q(\EX_LS_typ [0] ), .QN(_08140_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q ( .D(_00195_ ), .CK(_08028_ ), .Q(\ID_EX_csr [11] ), .QN(_08139_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_1 ( .D(_00196_ ), .CK(_08028_ ), .Q(\ID_EX_csr [10] ), .QN(_08138_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_10 ( .D(_00197_ ), .CK(_08028_ ), .Q(\ID_EX_csr [1] ), .QN(_08137_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_11 ( .D(_00198_ ), .CK(_08028_ ), .Q(\ID_EX_csr [0] ), .QN(_08136_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_2 ( .D(_00199_ ), .CK(_08028_ ), .Q(\ID_EX_csr [9] ), .QN(_08135_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_3 ( .D(_00200_ ), .CK(_08028_ ), .Q(\ID_EX_csr [8] ), .QN(_08134_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_4 ( .D(_00201_ ), .CK(_08028_ ), .Q(\ID_EX_csr [7] ), .QN(_08133_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_5 ( .D(_00202_ ), .CK(_08028_ ), .Q(\ID_EX_csr [6] ), .QN(_08132_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_6 ( .D(_00203_ ), .CK(_08028_ ), .Q(\ID_EX_csr [5] ), .QN(_08131_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_7 ( .D(_00204_ ), .CK(_08028_ ), .Q(\ID_EX_csr [4] ), .QN(_08130_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_8 ( .D(_00205_ ), .CK(_08028_ ), .Q(\ID_EX_csr [3] ), .QN(_08129_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_9 ( .D(_00206_ ), .CK(_08028_ ), .Q(\ID_EX_csr [2] ), .QN(_08128_ ) );
DFF_X1 \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q ( .D(_00207_ ), .CK(_08027_ ), .Q(exception_quest_IDU ), .QN(_08127_ ) );
DFF_X1 \myidu.fc_disenable_$_SDFFE_PP0P__Q ( .D(_00208_ ), .CK(_08026_ ), .Q(fc_disenable ), .QN(\myidu.fc_disenable_$_NOT__A_Y ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ), .CK(_08025_ ), .Q(\ID_EX_imm [31] ), .QN(_08444_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ), .CK(_08025_ ), .Q(\ID_EX_imm [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ), .CK(_08025_ ), .Q(\ID_EX_imm [21] ), .QN(_08445_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ), .CK(_08025_ ), .Q(\ID_EX_imm [20] ), .QN(_08446_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ), .CK(_08025_ ), .Q(\ID_EX_imm [19] ), .QN(_08447_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ), .CK(_08025_ ), .Q(\ID_EX_imm [18] ), .QN(_08448_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ), .CK(_08025_ ), .Q(\ID_EX_imm [17] ), .QN(_08449_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ), .CK(_08025_ ), .Q(\ID_EX_imm [16] ), .QN(_08450_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ), .CK(_08025_ ), .Q(\ID_EX_imm [15] ), .QN(_08451_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ), .CK(_08025_ ), .Q(\ID_EX_imm [14] ), .QN(_08452_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ), .CK(_08025_ ), .Q(\ID_EX_imm [13] ), .QN(_08453_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ), .CK(_08025_ ), .Q(\ID_EX_imm [12] ), .QN(_08454_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ), .CK(_08025_ ), .Q(\ID_EX_imm [29] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ), .CK(_08025_ ), .Q(\ID_EX_imm [11] ), .QN(_08455_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ), .CK(_08025_ ), .Q(\ID_EX_imm [10] ), .QN(_08456_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ), .CK(_08025_ ), .Q(\ID_EX_imm [9] ), .QN(_08457_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ), .CK(_08025_ ), .Q(\ID_EX_imm [8] ), .QN(_08458_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ), .CK(_08025_ ), .Q(\ID_EX_imm [7] ), .QN(_08459_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ), .CK(_08025_ ), .Q(\ID_EX_imm [6] ), .QN(_08460_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ), .CK(_08025_ ), .Q(\ID_EX_imm [5] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ), .CK(_08025_ ), .Q(\ID_EX_imm [4] ), .QN(_08461_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ), .CK(_08025_ ), .Q(\ID_EX_imm [3] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ), .CK(_08025_ ), .Q(\ID_EX_imm [2] ), .QN(_08462_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ), .CK(_08025_ ), .Q(\ID_EX_imm [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ), .CK(_08025_ ), .Q(\ID_EX_imm [1] ), .QN(_08463_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ), .CK(_08025_ ), .Q(\ID_EX_imm [0] ), .QN(_08464_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ), .CK(_08025_ ), .Q(\ID_EX_imm [27] ), .QN(_08465_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ), .CK(_08025_ ), .Q(\ID_EX_imm [26] ), .QN(_08466_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ), .CK(_08025_ ), .Q(\ID_EX_imm [25] ), .QN(_08467_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ), .CK(_08025_ ), .Q(\ID_EX_imm [24] ), .QN(_08468_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ), .CK(_08025_ ), .Q(\ID_EX_imm [23] ), .QN(_08469_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ), .CK(_08025_ ), .Q(\ID_EX_imm [22] ), .QN(_08470_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08024_ ), .Q(\ID_EX_pc [31] ), .QN(_08471_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08024_ ), .Q(\ID_EX_pc [30] ), .QN(_08472_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08024_ ), .Q(\ID_EX_pc [21] ), .QN(_08473_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08024_ ), .Q(\ID_EX_pc [20] ), .QN(_08474_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08024_ ), .Q(\ID_EX_pc [19] ), .QN(_08475_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08024_ ), .Q(\ID_EX_pc [18] ), .QN(_08476_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08024_ ), .Q(\ID_EX_pc [17] ), .QN(_08477_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08024_ ), .Q(\ID_EX_pc [16] ), .QN(_08478_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08024_ ), .Q(\ID_EX_pc [15] ), .QN(_08479_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08024_ ), .Q(\ID_EX_pc [14] ), .QN(_08480_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08024_ ), .Q(\ID_EX_pc [13] ), .QN(_08481_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08024_ ), .Q(\ID_EX_pc [12] ), .QN(_08482_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08024_ ), .Q(\ID_EX_pc [29] ), .QN(_08483_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08024_ ), .Q(\ID_EX_pc [11] ), .QN(_08484_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08024_ ), .Q(\ID_EX_pc [10] ), .QN(_08485_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08024_ ), .Q(\ID_EX_pc [9] ), .QN(_08486_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08024_ ), .Q(\ID_EX_pc [8] ), .QN(_08487_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08024_ ), .Q(\ID_EX_pc [7] ), .QN(_08488_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08024_ ), .Q(\ID_EX_pc [6] ), .QN(_08489_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08024_ ), .Q(\ID_EX_pc [5] ), .QN(_08490_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_08024_ ), .Q(\ID_EX_pc [4] ), .QN(_08491_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_28 ( .D(\IF_ID_pc [3] ), .CK(_08024_ ), .Q(\ID_EX_pc [3] ), .QN(_08492_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_29 ( .D(\IF_ID_pc [2] ), .CK(_08024_ ), .Q(\ID_EX_pc [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08024_ ), .Q(\ID_EX_pc [28] ), .QN(_08493_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_30 ( .D(\IF_ID_pc [1] ), .CK(_08024_ ), .Q(\ID_EX_pc [1] ), .QN(_08494_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_31 ( .D(\IF_ID_pc [0] ), .CK(_08024_ ), .Q(\ID_EX_pc [0] ), .QN(_08495_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08024_ ), .Q(\ID_EX_pc [27] ), .QN(_08496_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08024_ ), .Q(\ID_EX_pc [26] ), .QN(_08497_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08024_ ), .Q(\ID_EX_pc [25] ), .QN(_08498_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08024_ ), .Q(\ID_EX_pc [24] ), .QN(_08499_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08024_ ), .Q(\ID_EX_pc [23] ), .QN(_08500_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08024_ ), .Q(\ID_EX_pc [22] ), .QN(_08126_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q ( .D(_00209_ ), .CK(_08023_ ), .Q(\ID_EX_rd [4] ), .QN(_08125_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_1 ( .D(_00210_ ), .CK(_08023_ ), .Q(\ID_EX_rd [3] ), .QN(_08124_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_2 ( .D(_00211_ ), .CK(_08023_ ), .Q(\ID_EX_rd [2] ), .QN(_08123_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_3 ( .D(_00212_ ), .CK(_08023_ ), .Q(\ID_EX_rd [1] ), .QN(_08122_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_4 ( .D(_00213_ ), .CK(_08023_ ), .Q(\ID_EX_rd [0] ), .QN(_08121_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q ( .D(_00214_ ), .CK(_08022_ ), .Q(\ID_EX_rs1 [4] ), .QN(_08120_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1 ( .D(_00215_ ), .CK(_08022_ ), .Q(\ID_EX_rs1 [3] ), .QN(_08119_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00217_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08117_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2 ( .D(_00216_ ), .CK(_08022_ ), .Q(\ID_EX_rs1 [2] ), .QN(_08118_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00219_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08115_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3 ( .D(_00218_ ), .CK(_08022_ ), .Q(\ID_EX_rs1 [1] ), .QN(_08116_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00221_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08113_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4 ( .D(_00220_ ), .CK(_08022_ ), .Q(\ID_EX_rs1 [0] ), .QN(_08114_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00223_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08111_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q ( .D(_00222_ ), .CK(_08021_ ), .Q(\ID_EX_rs2 [4] ), .QN(_08112_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1 ( .D(_00224_ ), .CK(_08021_ ), .Q(\ID_EX_rs2 [3] ), .QN(_08110_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00226_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08108_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2 ( .D(_00225_ ), .CK(_08021_ ), .Q(\ID_EX_rs2 [2] ), .QN(_08109_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00228_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08106_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3 ( .D(_00227_ ), .CK(_08021_ ), .Q(\ID_EX_rs2 [1] ), .QN(_08107_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00230_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08104_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4 ( .D(_00229_ ), .CK(_08021_ ), .Q(\ID_EX_rs2 [0] ), .QN(_08105_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00232_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08102_ ) );
DFF_X1 \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q ( .D(_00231_ ), .CK(_08020_ ), .Q(\myidu.stall_quest_fencei ), .QN(_08103_ ) );
DFF_X1 \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q ( .D(_00233_ ), .CK(_08019_ ), .Q(\myidu.stall_quest_loaduse ), .QN(_08101_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q ( .D(\myidu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myidu.state [2] ), .QN(_08502_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q_1 ( .D(\myidu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \myidu.state_$_DFF_P__Q_2 ( .D(\myidu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q ( .D(_00234_ ), .CK(_08018_ ), .Q(\ID_EX_typ [7] ), .QN(_08501_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_1 ( .D(_00235_ ), .CK(_08018_ ), .Q(\ID_EX_typ [6] ), .QN(_08100_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_2 ( .D(_00236_ ), .CK(_08018_ ), .Q(\ID_EX_typ [5] ), .QN(_08099_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_3 ( .D(_00237_ ), .CK(_08018_ ), .Q(\ID_EX_typ [4] ), .QN(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_4 ( .D(_00238_ ), .CK(_08018_ ), .Q(\ID_EX_typ [3] ), .QN(_08098_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_5 ( .D(_00239_ ), .CK(_08018_ ), .Q(\ID_EX_typ [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_6 ( .D(_00240_ ), .CK(_08018_ ), .Q(\ID_EX_typ [1] ), .QN(_08097_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_7 ( .D(_00241_ ), .CK(_08018_ ), .Q(\ID_EX_typ [0] ), .QN(_08503_ ) );
DFF_X1 \myifu.check_assert_$_DFFE_PP__Q ( .D(\myifu.state [1] ), .CK(_08017_ ), .Q(check_assert ), .QN(_08504_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ), .CK(_08016_ ), .Q(\IF_ID_inst [31] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ), .CK(_08016_ ), .Q(\IF_ID_inst [30] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ), .CK(_08016_ ), .Q(\IF_ID_inst [21] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ), .CK(_08016_ ), .Q(\IF_ID_inst [20] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ), .CK(_08016_ ), .Q(\IF_ID_inst [19] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ), .CK(_08016_ ), .Q(\IF_ID_inst [18] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ), .CK(_08016_ ), .Q(\IF_ID_inst [17] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ), .CK(_08016_ ), .Q(\IF_ID_inst [16] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ), .CK(_08016_ ), .Q(\IF_ID_inst [15] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ), .CK(_08016_ ), .Q(\IF_ID_inst [14] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ), .CK(_08016_ ), .Q(\IF_ID_inst [13] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ), .CK(_08016_ ), .Q(\IF_ID_inst [12] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ), .CK(_08016_ ), .Q(\IF_ID_inst [29] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ), .CK(_08016_ ), .Q(\IF_ID_inst [11] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ), .CK(_08016_ ), .Q(\IF_ID_inst [10] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ), .CK(_08016_ ), .Q(\IF_ID_inst [9] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ), .CK(_08016_ ), .Q(\IF_ID_inst [8] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ), .CK(_08016_ ), .Q(\IF_ID_inst [7] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ), .CK(_08016_ ), .Q(\IF_ID_inst [6] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ), .CK(_08016_ ), .Q(\IF_ID_inst [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ), .CK(_08016_ ), .Q(\IF_ID_inst [4] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ), .CK(_08016_ ), .Q(\IF_ID_inst [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ), .CK(_08016_ ), .Q(\IF_ID_inst [2] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ), .CK(_08016_ ), .Q(\IF_ID_inst [28] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ), .CK(_08016_ ), .Q(\IF_ID_inst [1] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ), .CK(_08016_ ), .Q(\IF_ID_inst [0] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ), .CK(_08016_ ), .Q(\IF_ID_inst [27] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ), .CK(_08016_ ), .Q(\IF_ID_inst [26] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ), .CK(_08016_ ), .Q(\IF_ID_inst [25] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ), .CK(_08016_ ), .Q(\IF_ID_inst [24] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ), .CK(_08016_ ), .Q(\IF_ID_inst [23] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ), .CK(_08016_ ), .Q(\IF_ID_inst [22] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][31] ), .QN(_08505_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][30] ), .QN(_08506_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][21] ), .QN(_08507_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][20] ), .QN(_08508_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][19] ), .QN(_08509_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][18] ), .QN(_08510_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][17] ), .QN(_08511_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][16] ), .QN(_08512_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][15] ), .QN(_08513_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][14] ), .QN(_08514_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][13] ), .QN(_08515_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][12] ), .QN(_08516_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][29] ), .QN(_08517_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][11] ), .QN(_08518_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][10] ), .QN(_08519_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][9] ), .QN(_08520_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][8] ), .QN(_08521_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][7] ), .QN(_08522_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][6] ), .QN(_08523_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][5] ), .QN(_08524_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][4] ), .QN(_08525_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][3] ), .QN(_08526_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][2] ), .QN(_08527_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][28] ), .QN(_08528_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][1] ), .QN(_08529_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][0] ), .QN(_08530_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][27] ), .QN(_08531_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][26] ), .QN(_08532_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][25] ), .QN(_08533_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][24] ), .QN(_08534_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][23] ), .QN(_08535_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08015_ ), .Q(\myifu.myicache.data[0][22] ), .QN(_08536_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][31] ), .QN(_08537_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][30] ), .QN(_08538_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][21] ), .QN(_08539_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][20] ), .QN(_08540_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][19] ), .QN(_08541_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][18] ), .QN(_08542_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][17] ), .QN(_08543_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][16] ), .QN(_08544_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][15] ), .QN(_08545_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][14] ), .QN(_08546_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][13] ), .QN(_08547_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][12] ), .QN(_08548_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][29] ), .QN(_08549_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][11] ), .QN(_08550_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][10] ), .QN(_08551_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][9] ), .QN(_08552_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][8] ), .QN(_08553_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][7] ), .QN(_08554_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][6] ), .QN(_08555_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][5] ), .QN(_08556_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][4] ), .QN(_08557_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][3] ), .QN(_08558_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][2] ), .QN(_08559_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][28] ), .QN(_08560_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][1] ), .QN(_08561_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][0] ), .QN(_08562_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][27] ), .QN(_08563_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][26] ), .QN(_08564_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][25] ), .QN(_08565_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][24] ), .QN(_08566_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][23] ), .QN(_08567_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08014_ ), .Q(\myifu.myicache.data[1][22] ), .QN(_08568_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][31] ), .QN(_08569_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][30] ), .QN(_08570_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][21] ), .QN(_08571_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][20] ), .QN(_08572_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][19] ), .QN(_08573_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][18] ), .QN(_08574_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][17] ), .QN(_08575_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][16] ), .QN(_08576_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][15] ), .QN(_08577_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][14] ), .QN(_08578_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][13] ), .QN(_08579_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][12] ), .QN(_08580_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][29] ), .QN(_08581_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][11] ), .QN(_08582_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][10] ), .QN(_08583_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][9] ), .QN(_08584_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][8] ), .QN(_08585_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][7] ), .QN(_08586_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][6] ), .QN(_08587_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][5] ), .QN(_08588_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][4] ), .QN(_08589_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][3] ), .QN(_08590_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][2] ), .QN(_08591_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][28] ), .QN(_08592_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][1] ), .QN(_08593_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][0] ), .QN(_08594_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][27] ), .QN(_08595_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][26] ), .QN(_08596_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][25] ), .QN(_08597_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][24] ), .QN(_08598_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][23] ), .QN(_08599_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08013_ ), .Q(\myifu.myicache.data[2][22] ), .QN(_08600_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][31] ), .QN(_08601_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][30] ), .QN(_08602_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][21] ), .QN(_08603_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][20] ), .QN(_08604_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][19] ), .QN(_08605_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][18] ), .QN(_08606_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][17] ), .QN(_08607_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][16] ), .QN(_08608_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][15] ), .QN(_08609_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][14] ), .QN(_08610_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][13] ), .QN(_08611_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][12] ), .QN(_08612_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][29] ), .QN(_08613_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][11] ), .QN(_08614_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][10] ), .QN(_08615_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][9] ), .QN(_08616_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][8] ), .QN(_08617_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][7] ), .QN(_08618_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][6] ), .QN(_08619_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][5] ), .QN(_08620_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][4] ), .QN(_08621_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][3] ), .QN(_08622_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][2] ), .QN(_08623_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][28] ), .QN(_08624_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][1] ), .QN(_08625_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][0] ), .QN(_08626_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][27] ), .QN(_08627_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][26] ), .QN(_08628_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][25] ), .QN(_08629_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][24] ), .QN(_08630_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][23] ), .QN(_08631_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08012_ ), .Q(\myifu.myicache.data[3][22] ), .QN(_08632_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][31] ), .QN(_08633_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][30] ), .QN(_08634_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][21] ), .QN(_08635_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][20] ), .QN(_08636_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][19] ), .QN(_08637_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][18] ), .QN(_08638_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][17] ), .QN(_08639_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][16] ), .QN(_08640_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][15] ), .QN(_08641_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][14] ), .QN(_08642_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][13] ), .QN(_08643_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][12] ), .QN(_08644_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][29] ), .QN(_08645_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][11] ), .QN(_08646_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][10] ), .QN(_08647_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][9] ), .QN(_08648_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][8] ), .QN(_08649_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][7] ), .QN(_08650_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][6] ), .QN(_08651_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][5] ), .QN(_08652_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][4] ), .QN(_08653_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][3] ), .QN(_08654_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][2] ), .QN(_08655_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][28] ), .QN(_08656_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][1] ), .QN(_08657_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][0] ), .QN(_08658_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][27] ), .QN(_08659_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][26] ), .QN(_08660_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][25] ), .QN(_08661_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][24] ), .QN(_08662_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][23] ), .QN(_08663_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08011_ ), .Q(\myifu.myicache.data[4][22] ), .QN(_08664_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][31] ), .QN(_08665_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][30] ), .QN(_08666_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][21] ), .QN(_08667_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][20] ), .QN(_08668_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][19] ), .QN(_08669_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][18] ), .QN(_08670_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][17] ), .QN(_08671_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][16] ), .QN(_08672_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][15] ), .QN(_08673_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][14] ), .QN(_08674_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][13] ), .QN(_08675_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][12] ), .QN(_08676_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][29] ), .QN(_08677_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][11] ), .QN(_08678_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][10] ), .QN(_08679_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][9] ), .QN(_08680_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][8] ), .QN(_08681_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][7] ), .QN(_08682_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][6] ), .QN(_08683_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][5] ), .QN(_08684_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][4] ), .QN(_08685_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][3] ), .QN(_08686_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][2] ), .QN(_08687_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][28] ), .QN(_08688_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][1] ), .QN(_08689_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][0] ), .QN(_08690_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][27] ), .QN(_08691_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][26] ), .QN(_08692_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][25] ), .QN(_08693_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][24] ), .QN(_08694_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][23] ), .QN(_08695_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08010_ ), .Q(\myifu.myicache.data[5][22] ), .QN(_08696_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][31] ), .QN(_08697_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][30] ), .QN(_08698_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][21] ), .QN(_08699_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][20] ), .QN(_08700_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][19] ), .QN(_08701_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][18] ), .QN(_08702_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][17] ), .QN(_08703_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][16] ), .QN(_08704_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][15] ), .QN(_08705_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][14] ), .QN(_08706_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][13] ), .QN(_08707_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][12] ), .QN(_08708_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][29] ), .QN(_08709_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][11] ), .QN(_08710_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][10] ), .QN(_08711_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][9] ), .QN(_08712_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][8] ), .QN(_08713_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][7] ), .QN(_08714_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][6] ), .QN(_08715_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][5] ), .QN(_08716_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][4] ), .QN(_08717_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][3] ), .QN(_08718_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][2] ), .QN(_08719_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][28] ), .QN(_08720_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][1] ), .QN(_08721_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][0] ), .QN(_08722_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][27] ), .QN(_08723_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][26] ), .QN(_08724_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][25] ), .QN(_08725_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][24] ), .QN(_08726_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][23] ), .QN(_08727_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08009_ ), .Q(\myifu.myicache.data[6][22] ), .QN(_08728_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][31] ), .QN(_08729_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][30] ), .QN(_08730_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][21] ), .QN(_08731_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][20] ), .QN(_08732_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][19] ), .QN(_08733_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][18] ), .QN(_08734_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][17] ), .QN(_08735_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][16] ), .QN(_08736_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][15] ), .QN(_08737_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][14] ), .QN(_08738_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][13] ), .QN(_08739_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][12] ), .QN(_08740_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][29] ), .QN(_08741_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][11] ), .QN(_08742_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][10] ), .QN(_08743_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][9] ), .QN(_08744_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][8] ), .QN(_08745_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][7] ), .QN(_08746_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][6] ), .QN(_08747_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][5] ), .QN(_08748_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][4] ), .QN(_08749_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][3] ), .QN(_08750_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][2] ), .QN(_08751_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][28] ), .QN(_08752_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][1] ), .QN(_08753_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][0] ), .QN(_08754_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][27] ), .QN(_08755_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][26] ), .QN(_08756_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][25] ), .QN(_08757_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][24] ), .QN(_08758_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][23] ), .QN(_08759_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08008_ ), .Q(\myifu.myicache.data[7][22] ), .QN(_08760_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][26] ), .QN(_08761_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][25] ), .QN(_08762_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][16] ), .QN(_08763_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][15] ), .QN(_08764_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][14] ), .QN(_08765_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][13] ), .QN(_08766_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][12] ), .QN(_08767_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][11] ), .QN(_08768_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][10] ), .QN(_08769_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][9] ), .QN(_08770_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][8] ), .QN(_08771_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][7] ), .QN(_08772_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][24] ), .QN(_08773_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][6] ), .QN(_08774_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][5] ), .QN(_08775_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][4] ), .QN(_08776_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][3] ), .QN(_08777_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][2] ), .QN(_08778_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][1] ), .QN(_08779_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][0] ), .QN(_08780_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][23] ), .QN(_08781_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][22] ), .QN(_08782_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][21] ), .QN(_08783_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][20] ), .QN(_08784_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][19] ), .QN(_08785_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][18] ), .QN(_08786_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08007_ ), .Q(\myifu.myicache.tag[0][17] ), .QN(_08787_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][26] ), .QN(_08788_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][25] ), .QN(_08789_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][16] ), .QN(_08790_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][15] ), .QN(_08791_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][14] ), .QN(_08792_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][13] ), .QN(_08793_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][12] ), .QN(_08794_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][11] ), .QN(_08795_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][10] ), .QN(_08796_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][9] ), .QN(_08797_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][8] ), .QN(_08798_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][7] ), .QN(_08799_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][24] ), .QN(_08800_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][6] ), .QN(_08801_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][5] ), .QN(_08802_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][4] ), .QN(_08803_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][3] ), .QN(_08804_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][2] ), .QN(_08805_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][1] ), .QN(_08806_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][0] ), .QN(_08807_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][23] ), .QN(_08808_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][22] ), .QN(_08809_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][21] ), .QN(_08810_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][20] ), .QN(_08811_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][19] ), .QN(_08812_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][18] ), .QN(_08813_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08006_ ), .Q(\myifu.myicache.tag[1][17] ), .QN(_08814_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][26] ), .QN(_08815_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][25] ), .QN(_08816_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][16] ), .QN(_08817_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][15] ), .QN(_08818_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][14] ), .QN(_08819_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][13] ), .QN(_08820_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][12] ), .QN(_08821_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][11] ), .QN(_08822_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][10] ), .QN(_08823_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][9] ), .QN(_08824_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][8] ), .QN(_08825_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][7] ), .QN(_08826_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][24] ), .QN(_08827_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][6] ), .QN(_08828_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][5] ), .QN(_08829_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][4] ), .QN(_08830_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][3] ), .QN(_08831_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][2] ), .QN(_08832_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][1] ), .QN(_08833_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][0] ), .QN(_08834_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][23] ), .QN(_08835_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][22] ), .QN(_08836_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][21] ), .QN(_08837_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][20] ), .QN(_08838_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][19] ), .QN(_08839_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][18] ), .QN(_08840_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08005_ ), .Q(\myifu.myicache.tag[2][17] ), .QN(_08841_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][26] ), .QN(_08842_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][25] ), .QN(_08843_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][16] ), .QN(_08844_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][15] ), .QN(_08845_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][14] ), .QN(_08846_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][13] ), .QN(_08847_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][12] ), .QN(_08848_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][11] ), .QN(_08849_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][10] ), .QN(_08850_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][9] ), .QN(_08851_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][8] ), .QN(_08852_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][7] ), .QN(_08853_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][24] ), .QN(_08854_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][6] ), .QN(_08855_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][5] ), .QN(_08856_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][4] ), .QN(_08857_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][3] ), .QN(_08858_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][2] ), .QN(_08859_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][1] ), .QN(_08860_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][0] ), .QN(_08861_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][23] ), .QN(_08862_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][22] ), .QN(_08863_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][21] ), .QN(_08864_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][20] ), .QN(_08865_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][19] ), .QN(_08866_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][18] ), .QN(_08867_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08004_ ), .Q(\myifu.myicache.tag[3][17] ), .QN(_08096_ ) );
DFF_X1 \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_00242_ ), .CK(_08003_ ), .Q(\myifu.myicache.valid [0] ), .QN(_08095_ ) );
DFF_X1 \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_00243_ ), .CK(_08002_ ), .Q(\myifu.myicache.valid [1] ), .QN(_08094_ ) );
DFF_X1 \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_00244_ ), .CK(_08001_ ), .Q(\myifu.myicache.valid [2] ), .QN(_08868_ ) );
DFF_X1 \myifu.myicache.valid[3]_$_DFFE_PP__Q ( .D(\myifu.wen_$_ANDNOT__A_Y ), .CK(_08000_ ), .Q(\myifu.myicache.valid [3] ), .QN(_08093_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q ( .D(_00245_ ), .CK(_07999_ ), .Q(\IF_ID_pc [0] ), .QN(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00246_ ), .CK(_07998_ ), .Q(\IF_ID_pc [30] ), .QN(_08092_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00247_ ), .CK(_07998_ ), .Q(\IF_ID_pc [21] ), .QN(_08091_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00248_ ), .CK(_07998_ ), .Q(\IF_ID_pc [20] ), .QN(_08090_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00249_ ), .CK(_07998_ ), .Q(\IF_ID_pc [19] ), .QN(_08089_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00250_ ), .CK(_07998_ ), .Q(\IF_ID_pc [18] ), .QN(_08088_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00251_ ), .CK(_07998_ ), .Q(\IF_ID_pc [17] ), .QN(_08087_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00252_ ), .CK(_07998_ ), .Q(\IF_ID_pc [16] ), .QN(_08086_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00253_ ), .CK(_07998_ ), .Q(\IF_ID_pc [15] ), .QN(_08085_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00254_ ), .CK(_07998_ ), .Q(\IF_ID_pc [14] ), .QN(_08084_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00255_ ), .CK(_07998_ ), .Q(\IF_ID_pc [13] ), .QN(_08083_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00256_ ), .CK(_07998_ ), .Q(\IF_ID_pc [12] ), .QN(_08082_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00257_ ), .CK(_07998_ ), .Q(\IF_ID_pc [29] ), .QN(_08081_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00258_ ), .CK(_07998_ ), .Q(\IF_ID_pc [11] ), .QN(_08080_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00259_ ), .CK(_07998_ ), .Q(\IF_ID_pc [10] ), .QN(_08079_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00260_ ), .CK(_07998_ ), .Q(\IF_ID_pc [9] ), .QN(_08078_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00261_ ), .CK(_07998_ ), .Q(\IF_ID_pc [8] ), .QN(_08077_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00262_ ), .CK(_07998_ ), .Q(\IF_ID_pc [7] ), .QN(_08076_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00263_ ), .CK(_07998_ ), .Q(\IF_ID_pc [6] ), .QN(_08075_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00264_ ), .CK(_07998_ ), .Q(\IF_ID_pc [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00265_ ), .CK(_07998_ ), .Q(\IF_ID_pc [4] ), .QN(_08074_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00267_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08073_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00266_ ), .CK(_07998_ ), .Q(\IF_ID_pc [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00269_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08071_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00268_ ), .CK(_07998_ ), .Q(\IF_ID_pc [2] ), .QN(_08072_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00270_ ), .CK(_07998_ ), .Q(\IF_ID_pc [28] ), .QN(_08070_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00271_ ), .CK(_07998_ ), .Q(\IF_ID_pc [1] ), .QN(_08069_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00272_ ), .CK(_07998_ ), .Q(\IF_ID_pc [27] ), .QN(_08068_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00273_ ), .CK(_07998_ ), .Q(\IF_ID_pc [26] ), .QN(_08067_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00274_ ), .CK(_07998_ ), .Q(\IF_ID_pc [25] ), .QN(_08066_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00275_ ), .CK(_07998_ ), .Q(\IF_ID_pc [24] ), .QN(_08065_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00276_ ), .CK(_07998_ ), .Q(\IF_ID_pc [23] ), .QN(_08064_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00277_ ), .CK(_07998_ ), .Q(\IF_ID_pc [22] ), .QN(_08063_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP1P__Q ( .D(_00278_ ), .CK(_07998_ ), .Q(\IF_ID_pc [31] ), .QN(_08062_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q ( .D(\myifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myifu.state [2] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.state_$_DFF_P__Q_1 ( .D(\myifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myifu.state [1] ), .QN(_08870_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q_2 ( .D(\myifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\myifu.state [0] ), .QN(_08061_ ) );
DFF_X1 \myifu.tmp_offset_$_SDFFE_PP0P__Q ( .D(_00279_ ), .CK(_07997_ ), .Q(\myifu.tmp_offset [2] ), .QN(_08869_ ) );
DFF_X1 \myifu.to_reset_$_SDFF_PP0__Q ( .D(_00281_ ), .CK(clock ), .Q(\myifu.to_reset ), .QN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ) );
DFF_X1 \myifu.wen_$_SDFFE_PP0P__Q ( .D(_00280_ ), .CK(_07996_ ), .Q(\myifu.myicache.valid_data_in ), .QN(_08060_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [31] ), .QN(_08871_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [30] ), .QN(_08872_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [21] ), .QN(_08873_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [20] ), .QN(_08874_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [19] ), .QN(_08875_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [18] ), .QN(_08876_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [17] ), .QN(_08877_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [16] ), .QN(_08878_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [15] ), .QN(_08879_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [14] ), .QN(_08880_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [13] ), .QN(_08881_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [12] ), .QN(_08882_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [29] ), .QN(_08883_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [11] ), .QN(_08884_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [10] ), .QN(_08885_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [9] ), .QN(_08886_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [8] ), .QN(_08887_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [7] ), .QN(_08888_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [6] ), .QN(_08889_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [5] ), .QN(_08890_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [4] ), .QN(_08891_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [3] ), .QN(_08892_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [2] ), .QN(_08893_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [28] ), .QN(_08894_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_30 ( .D(fanout_net_4 ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [1] ), .QN(_08895_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [0] ), .QN(_08896_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [27] ), .QN(_08897_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [26] ), .QN(_08898_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [25] ), .QN(_08899_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [24] ), .QN(_08900_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [23] ), .QN(_08901_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_07995_ ), .Q(\mylsu.araddr_tmp [22] ), .QN(_08902_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [31] ), .QN(_08903_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [30] ), .QN(_08904_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [21] ), .QN(_08905_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [20] ), .QN(_08906_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [19] ), .QN(_08907_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [18] ), .QN(_08908_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [17] ), .QN(_08909_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [16] ), .QN(_08910_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [15] ), .QN(_08911_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [14] ), .QN(_08912_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [13] ), .QN(_08913_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [12] ), .QN(_08914_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [29] ), .QN(_08915_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [11] ), .QN(_08916_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [10] ), .QN(_08917_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [9] ), .QN(_08918_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [8] ), .QN(_08919_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [7] ), .QN(_08920_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [6] ), .QN(_08921_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [5] ), .QN(_08922_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [4] ), .QN(_08923_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [3] ), .QN(_08924_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [2] ), .QN(_08925_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [28] ), .QN(_08926_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [1] ), .QN(_08927_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [0] ), .QN(_08928_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [27] ), .QN(_08929_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [26] ), .QN(_08930_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [25] ), .QN(_08931_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [24] ), .QN(_08932_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [23] ), .QN(_08933_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_07994_ ), .Q(\mylsu.awaddr_tmp [22] ), .QN(_08059_ ) );
DFF_X1 \mylsu.pc_out_$_SDFFE_PN0P__Q ( .D(_00282_ ), .CK(_07993_ ), .Q(LS_WB_pc ), .QN(_08058_ ) );
DFF_X1 \mylsu.previous_load_done_$_SDFFE_PN0P__Q ( .D(_00283_ ), .CK(_07992_ ), .Q(\mylsu.previous_load_done ), .QN(_08934_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q ( .D(\mylsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mylsu.state [4] ), .QN(_08935_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_1 ( .D(\mylsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mylsu.state [3] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_2 ( .D(\mylsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mylsu.state [2] ), .QN(_08936_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_3 ( .D(\mylsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\mylsu.state [1] ), .QN(_08937_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_4 ( .D(\mylsu.state_$_DFF_P__Q_4_D ), .CK(clock ), .Q(\mylsu.state [0] ), .QN(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q ( .D(\EX_LS_typ [2] ), .CK(_07995_ ), .Q(\mylsu.typ_tmp [2] ), .QN(\mylsu.typ_tmp_$_NOT__A_Y ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_typ [1] ), .CK(_07995_ ), .Q(\mylsu.typ_tmp [1] ), .QN(_08938_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_typ [0] ), .CK(_07995_ ), .Q(\mylsu.typ_tmp [0] ), .QN(_08057_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q ( .D(_00284_ ), .CK(_07995_ ), .Q(\LS_WB_waddr_csreg [11] ), .QN(_08056_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_1 ( .D(_00285_ ), .CK(_07995_ ), .Q(\LS_WB_waddr_csreg [10] ), .QN(_08055_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_2 ( .D(_00286_ ), .CK(_07995_ ), .Q(\LS_WB_waddr_csreg [7] ), .QN(_08054_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_3 ( .D(_00287_ ), .CK(_07995_ ), .Q(\LS_WB_waddr_csreg [5] ), .QN(_08053_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_4 ( .D(_00288_ ), .CK(_07995_ ), .Q(\LS_WB_waddr_csreg [4] ), .QN(_08052_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_5 ( .D(_00289_ ), .CK(_07995_ ), .Q(\LS_WB_waddr_csreg [3] ), .QN(_08051_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_6 ( .D(_00290_ ), .CK(_07995_ ), .Q(\LS_WB_waddr_csreg [2] ), .QN(_08050_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_7 ( .D(_00291_ ), .CK(_07995_ ), .Q(\LS_WB_waddr_csreg [1] ), .QN(_08049_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q ( .D(_00292_ ), .CK(_07995_ ), .Q(\LS_WB_waddr_csreg [9] ), .QN(_08048_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_1 ( .D(_00293_ ), .CK(_07995_ ), .Q(\LS_WB_waddr_csreg [8] ), .QN(_08047_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_2 ( .D(_00294_ ), .CK(_07995_ ), .Q(\LS_WB_waddr_csreg [6] ), .QN(_08046_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_3 ( .D(_00295_ ), .CK(_07995_ ), .Q(\LS_WB_waddr_csreg [0] ), .QN(_08939_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q ( .D(\EX_LS_dest_reg [3] ), .CK(_07995_ ), .Q(\LS_WB_waddr_reg [3] ), .QN(_08940_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_reg [2] ), .CK(_07995_ ), .Q(\LS_WB_waddr_reg [2] ), .QN(_08941_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_reg [1] ), .CK(_07995_ ), .Q(\LS_WB_waddr_reg [1] ), .QN(_08942_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_reg [0] ), .CK(_07995_ ), .Q(\LS_WB_waddr_reg [0] ), .QN(_08943_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [31] ), .QN(_08944_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [30] ), .QN(_08945_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [21] ), .QN(_08946_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [20] ), .QN(_08947_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [19] ), .QN(_08948_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [18] ), .QN(_08949_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [17] ), .QN(_08950_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [16] ), .QN(_08951_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [15] ), .QN(_08952_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [14] ), .QN(_08953_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [13] ), .QN(_08954_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [12] ), .QN(_08955_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [29] ), .QN(_08956_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [11] ), .QN(_08957_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [10] ), .QN(_08958_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [9] ), .QN(_08959_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [8] ), .QN(_08960_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [7] ), .QN(_08961_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [6] ), .QN(_08962_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [5] ), .QN(_08963_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [4] ), .QN(_08964_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [3] ), .QN(_08965_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [2] ), .QN(_08966_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [28] ), .QN(_08967_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [1] ), .QN(_08968_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [0] ), .QN(_08969_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [27] ), .QN(_08970_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [26] ), .QN(_08971_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [25] ), .QN(_08972_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [24] ), .QN(_08973_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [23] ), .QN(_08974_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ), .CK(_07995_ ), .Q(\LS_WB_wdata_csreg [22] ), .QN(_08975_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [31] ), .QN(_08976_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [30] ), .QN(_08977_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [21] ), .QN(_08978_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [20] ), .QN(_08979_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [19] ), .QN(_08980_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [18] ), .QN(_08981_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [17] ), .QN(_08982_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [16] ), .QN(_08983_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [15] ), .QN(_08984_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [14] ), .QN(_08985_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [13] ), .QN(_08986_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [12] ), .QN(_08987_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [29] ), .QN(_08988_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [11] ), .QN(_08989_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [10] ), .QN(_08990_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [9] ), .QN(_08991_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [8] ), .QN(_08992_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [7] ), .QN(_08993_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [6] ), .QN(_08994_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [5] ), .QN(_08995_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [4] ), .QN(_08996_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [3] ), .QN(_08997_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [2] ), .QN(_08998_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [28] ), .QN(_08999_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [1] ), .QN(_09000_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [0] ), .QN(_09001_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [27] ), .QN(_09002_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [26] ), .QN(_09003_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [25] ), .QN(_09004_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [24] ), .QN(_09005_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [23] ), .QN(_09006_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ), .CK(_07991_ ), .Q(\LS_WB_wdata_reg [22] ), .QN(_08045_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q ( .D(_00296_ ), .CK(_07990_ ), .Q(\LS_WB_wen_csreg [7] ), .QN(_08044_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_1 ( .D(_00297_ ), .CK(_07990_ ), .Q(\LS_WB_wen_csreg [6] ), .QN(_08043_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_2 ( .D(_00298_ ), .CK(_07990_ ), .Q(\LS_WB_wen_csreg [3] ), .QN(_08042_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_3 ( .D(_00299_ ), .CK(_07990_ ), .Q(\LS_WB_wen_csreg [2] ), .QN(_08041_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_4 ( .D(_00300_ ), .CK(_07990_ ), .Q(\LS_WB_wen_csreg [1] ), .QN(_08040_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_5 ( .D(_00301_ ), .CK(_07990_ ), .Q(\LS_WB_wen_csreg [0] ), .QN(_08039_ ) );
DFF_X1 \mylsu.wen_reg_$_SDFFE_PN0P__Q ( .D(_00302_ ), .CK(_07990_ ), .Q(LS_WB_wen_reg ), .QN(_09007_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q ( .D(\myminixbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myminixbar.state [2] ), .QN(_09008_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q_1 ( .D(\myminixbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myminixbar.state [0] ), .QN(_09009_ ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07989_ ), .Q(\myreg.Reg[0][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07988_ ), .Q(\myreg.Reg[10][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07987_ ), .Q(\myreg.Reg[11][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07986_ ), .Q(\myreg.Reg[12][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07985_ ), .Q(\myreg.Reg[13][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07984_ ), .Q(\myreg.Reg[14][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07983_ ), .Q(\myreg.Reg[15][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07982_ ), .Q(\myreg.Reg[1][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07981_ ), .Q(\myreg.Reg[2][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07980_ ), .Q(\myreg.Reg[3][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07979_ ), .Q(\myreg.Reg[4][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07978_ ), .Q(\myreg.Reg[5][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07977_ ), .Q(\myreg.Reg[6][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07976_ ), .Q(\myreg.Reg[7][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07975_ ), .Q(\myreg.Reg[8][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07974_ ), .Q(\myreg.Reg[9][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mysc.loaduse_clear_$_SDFFE_PP0P__Q ( .D(_00303_ ), .CK(_07973_ ), .Q(loaduse_clear ), .QN(_09010_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q ( .D(\mysc.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mysc.state [2] ), .QN(_09011_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_1 ( .D(\mysc.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mysc.state [1] ), .QN(_09012_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_2 ( .D(\mysc.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mysc.state [0] ), .QN(_08038_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(\EX_LS_dest_csreg_mem [1] ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\ID_EX_typ [4] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_40 ) );
BUF_X8 fanout_buf_41 ( .A(\myifu.to_reset ), .Z(fanout_net_41 ) );
BUF_X8 fanout_buf_42 ( .A(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .Z(fanout_net_42 ) );

endmodule
